module core (clock,
    io_load_store_unsigned,
    io_meip,
    io_memory_read,
    io_memory_write,
    reset,
    io_fetch_address,
    io_fetch_data,
    io_memory_address,
    io_memory_read_data,
    io_memory_size,
    io_memory_write_data);
 input clock;
 output io_load_store_unsigned;
 input io_meip;
 output io_memory_read;
 output io_memory_write;
 input reset;
 output [31:0] io_fetch_address;
 input [31:0] io_fetch_data;
 output [31:0] io_memory_address;
 input [31:0] io_memory_read_data;
 output [1:0] io_memory_size;
 output [31:0] io_memory_write_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire \csr._csr_read_data_T_8[10] ;
 wire \csr._csr_read_data_T_8[11] ;
 wire \csr._csr_read_data_T_8[12] ;
 wire \csr._csr_read_data_T_8[13] ;
 wire \csr._csr_read_data_T_8[14] ;
 wire \csr._csr_read_data_T_8[15] ;
 wire \csr._csr_read_data_T_8[16] ;
 wire \csr._csr_read_data_T_8[17] ;
 wire \csr._csr_read_data_T_8[18] ;
 wire \csr._csr_read_data_T_8[19] ;
 wire \csr._csr_read_data_T_8[20] ;
 wire \csr._csr_read_data_T_8[21] ;
 wire \csr._csr_read_data_T_8[22] ;
 wire \csr._csr_read_data_T_8[23] ;
 wire \csr._csr_read_data_T_8[24] ;
 wire \csr._csr_read_data_T_8[25] ;
 wire \csr._csr_read_data_T_8[26] ;
 wire \csr._csr_read_data_T_8[27] ;
 wire \csr._csr_read_data_T_8[28] ;
 wire \csr._csr_read_data_T_8[29] ;
 wire \csr._csr_read_data_T_8[2] ;
 wire \csr._csr_read_data_T_8[30] ;
 wire \csr._csr_read_data_T_8[31] ;
 wire \csr._csr_read_data_T_8[3] ;
 wire \csr._csr_read_data_T_8[4] ;
 wire \csr._csr_read_data_T_8[5] ;
 wire \csr._csr_read_data_T_8[6] ;
 wire \csr._csr_read_data_T_8[7] ;
 wire \csr._csr_read_data_T_8[8] ;
 wire \csr._csr_read_data_T_8[9] ;
 wire \csr._csr_read_data_T_9[0] ;
 wire \csr._csr_read_data_T_9[1] ;
 wire \csr._csr_read_data_T_9[2] ;
 wire \csr._csr_read_data_T_9[31] ;
 wire \csr._csr_read_data_T_9[3] ;
 wire \csr._mcycle_T_2[0] ;
 wire \csr._mcycle_T_2[10] ;
 wire \csr._mcycle_T_2[11] ;
 wire \csr._mcycle_T_2[12] ;
 wire \csr._mcycle_T_2[13] ;
 wire \csr._mcycle_T_2[14] ;
 wire \csr._mcycle_T_2[15] ;
 wire \csr._mcycle_T_2[16] ;
 wire \csr._mcycle_T_2[17] ;
 wire \csr._mcycle_T_2[18] ;
 wire \csr._mcycle_T_2[19] ;
 wire \csr._mcycle_T_2[1] ;
 wire \csr._mcycle_T_2[20] ;
 wire \csr._mcycle_T_2[21] ;
 wire \csr._mcycle_T_2[22] ;
 wire \csr._mcycle_T_2[23] ;
 wire \csr._mcycle_T_2[24] ;
 wire \csr._mcycle_T_2[25] ;
 wire \csr._mcycle_T_2[26] ;
 wire \csr._mcycle_T_2[27] ;
 wire \csr._mcycle_T_2[28] ;
 wire \csr._mcycle_T_2[29] ;
 wire \csr._mcycle_T_2[2] ;
 wire \csr._mcycle_T_2[30] ;
 wire \csr._mcycle_T_2[31] ;
 wire \csr._mcycle_T_2[3] ;
 wire \csr._mcycle_T_2[4] ;
 wire \csr._mcycle_T_2[5] ;
 wire \csr._mcycle_T_2[6] ;
 wire \csr._mcycle_T_2[7] ;
 wire \csr._mcycle_T_2[8] ;
 wire \csr._mcycle_T_2[9] ;
 wire \csr._mcycle_T_3[32] ;
 wire \csr._mcycle_T_3[33] ;
 wire \csr._mcycle_T_3[34] ;
 wire \csr._mcycle_T_3[35] ;
 wire \csr._mcycle_T_3[36] ;
 wire \csr._mcycle_T_3[37] ;
 wire \csr._mcycle_T_3[38] ;
 wire \csr._mcycle_T_3[39] ;
 wire \csr._mcycle_T_3[40] ;
 wire \csr._mcycle_T_3[41] ;
 wire \csr._mcycle_T_3[42] ;
 wire \csr._mcycle_T_3[43] ;
 wire \csr._mcycle_T_3[44] ;
 wire \csr._mcycle_T_3[45] ;
 wire \csr._mcycle_T_3[46] ;
 wire \csr._mcycle_T_3[47] ;
 wire \csr._mcycle_T_3[48] ;
 wire \csr._mcycle_T_3[49] ;
 wire \csr._mcycle_T_3[50] ;
 wire \csr._mcycle_T_3[51] ;
 wire \csr._mcycle_T_3[52] ;
 wire \csr._mcycle_T_3[53] ;
 wire \csr._mcycle_T_3[54] ;
 wire \csr._mcycle_T_3[55] ;
 wire \csr._mcycle_T_3[56] ;
 wire \csr._mcycle_T_3[57] ;
 wire \csr._mcycle_T_3[58] ;
 wire \csr._mcycle_T_3[59] ;
 wire \csr._mcycle_T_3[60] ;
 wire \csr._mcycle_T_3[61] ;
 wire \csr._mcycle_T_3[62] ;
 wire \csr._mcycle_T_3[63] ;
 wire \csr._minstret_T_3[32] ;
 wire \csr._minstret_T_3[33] ;
 wire \csr._minstret_T_3[34] ;
 wire \csr._minstret_T_3[35] ;
 wire \csr._minstret_T_3[36] ;
 wire \csr._minstret_T_3[37] ;
 wire \csr._minstret_T_3[38] ;
 wire \csr._minstret_T_3[39] ;
 wire \csr._minstret_T_3[40] ;
 wire \csr._minstret_T_3[41] ;
 wire \csr._minstret_T_3[42] ;
 wire \csr._minstret_T_3[43] ;
 wire \csr._minstret_T_3[44] ;
 wire \csr._minstret_T_3[45] ;
 wire \csr._minstret_T_3[46] ;
 wire \csr._minstret_T_3[47] ;
 wire \csr._minstret_T_3[48] ;
 wire \csr._minstret_T_3[49] ;
 wire \csr._minstret_T_3[50] ;
 wire \csr._minstret_T_3[51] ;
 wire \csr._minstret_T_3[52] ;
 wire \csr._minstret_T_3[53] ;
 wire \csr._minstret_T_3[54] ;
 wire \csr._minstret_T_3[55] ;
 wire \csr._minstret_T_3[56] ;
 wire \csr._minstret_T_3[57] ;
 wire \csr._minstret_T_3[58] ;
 wire \csr._minstret_T_3[59] ;
 wire \csr._minstret_T_3[60] ;
 wire \csr._minstret_T_3[61] ;
 wire \csr._minstret_T_3[62] ;
 wire \csr._minstret_T_3[63] ;
 wire \csr.ie ;
 wire \csr.io_csr_address[0] ;
 wire \csr.io_csr_address[10] ;
 wire \csr.io_csr_address[11] ;
 wire \csr.io_csr_address[1] ;
 wire \csr.io_csr_address[2] ;
 wire \csr.io_csr_address[3] ;
 wire \csr.io_csr_address[4] ;
 wire \csr.io_csr_address[5] ;
 wire \csr.io_csr_address[6] ;
 wire \csr.io_csr_address[7] ;
 wire \csr.io_csr_address[8] ;
 wire \csr.io_csr_address[9] ;
 wire \csr.io_csr_write_address[0] ;
 wire \csr.io_csr_write_address[10] ;
 wire \csr.io_csr_write_address[11] ;
 wire \csr.io_csr_write_address[1] ;
 wire \csr.io_csr_write_address[2] ;
 wire \csr.io_csr_write_address[3] ;
 wire \csr.io_csr_write_address[4] ;
 wire \csr.io_csr_write_address[5] ;
 wire \csr.io_csr_write_address[6] ;
 wire \csr.io_csr_write_address[7] ;
 wire \csr.io_csr_write_address[8] ;
 wire \csr.io_csr_write_address[9] ;
 wire \csr.io_csr_write_enable ;
 wire \csr.io_ecause[0] ;
 wire \csr.io_ecause[1] ;
 wire \csr.io_ecause[2] ;
 wire \csr.io_inst_retired ;
 wire \csr.io_interrupt ;
 wire \csr.io_mem_pc[0] ;
 wire \csr.io_mem_pc[10] ;
 wire \csr.io_mem_pc[11] ;
 wire \csr.io_mem_pc[12] ;
 wire \csr.io_mem_pc[13] ;
 wire \csr.io_mem_pc[14] ;
 wire \csr.io_mem_pc[15] ;
 wire \csr.io_mem_pc[16] ;
 wire \csr.io_mem_pc[17] ;
 wire \csr.io_mem_pc[18] ;
 wire \csr.io_mem_pc[19] ;
 wire \csr.io_mem_pc[1] ;
 wire \csr.io_mem_pc[20] ;
 wire \csr.io_mem_pc[21] ;
 wire \csr.io_mem_pc[22] ;
 wire \csr.io_mem_pc[23] ;
 wire \csr.io_mem_pc[24] ;
 wire \csr.io_mem_pc[25] ;
 wire \csr.io_mem_pc[26] ;
 wire \csr.io_mem_pc[27] ;
 wire \csr.io_mem_pc[28] ;
 wire \csr.io_mem_pc[29] ;
 wire \csr.io_mem_pc[2] ;
 wire \csr.io_mem_pc[30] ;
 wire \csr.io_mem_pc[31] ;
 wire \csr.io_mem_pc[3] ;
 wire \csr.io_mem_pc[4] ;
 wire \csr.io_mem_pc[5] ;
 wire \csr.io_mem_pc[6] ;
 wire \csr.io_mem_pc[7] ;
 wire \csr.io_mem_pc[8] ;
 wire \csr.io_mem_pc[9] ;
 wire \csr.io_mret ;
 wire \csr.io_mret_vector[0] ;
 wire \csr.io_mret_vector[10] ;
 wire \csr.io_mret_vector[11] ;
 wire \csr.io_mret_vector[12] ;
 wire \csr.io_mret_vector[13] ;
 wire \csr.io_mret_vector[14] ;
 wire \csr.io_mret_vector[15] ;
 wire \csr.io_mret_vector[16] ;
 wire \csr.io_mret_vector[17] ;
 wire \csr.io_mret_vector[18] ;
 wire \csr.io_mret_vector[19] ;
 wire \csr.io_mret_vector[1] ;
 wire \csr.io_mret_vector[20] ;
 wire \csr.io_mret_vector[21] ;
 wire \csr.io_mret_vector[22] ;
 wire \csr.io_mret_vector[23] ;
 wire \csr.io_mret_vector[24] ;
 wire \csr.io_mret_vector[25] ;
 wire \csr.io_mret_vector[26] ;
 wire \csr.io_mret_vector[27] ;
 wire \csr.io_mret_vector[28] ;
 wire \csr.io_mret_vector[29] ;
 wire \csr.io_mret_vector[2] ;
 wire \csr.io_mret_vector[30] ;
 wire \csr.io_mret_vector[31] ;
 wire \csr.io_mret_vector[3] ;
 wire \csr.io_mret_vector[4] ;
 wire \csr.io_mret_vector[5] ;
 wire \csr.io_mret_vector[6] ;
 wire \csr.io_mret_vector[7] ;
 wire \csr.io_mret_vector[8] ;
 wire \csr.io_mret_vector[9] ;
 wire \csr.io_trapped ;
 wire \csr.mcycle[0] ;
 wire \csr.mcycle[10] ;
 wire \csr.mcycle[11] ;
 wire \csr.mcycle[12] ;
 wire \csr.mcycle[13] ;
 wire \csr.mcycle[14] ;
 wire \csr.mcycle[15] ;
 wire \csr.mcycle[16] ;
 wire \csr.mcycle[17] ;
 wire \csr.mcycle[18] ;
 wire \csr.mcycle[19] ;
 wire \csr.mcycle[1] ;
 wire \csr.mcycle[20] ;
 wire \csr.mcycle[21] ;
 wire \csr.mcycle[22] ;
 wire \csr.mcycle[23] ;
 wire \csr.mcycle[24] ;
 wire \csr.mcycle[25] ;
 wire \csr.mcycle[26] ;
 wire \csr.mcycle[27] ;
 wire \csr.mcycle[28] ;
 wire \csr.mcycle[29] ;
 wire \csr.mcycle[2] ;
 wire \csr.mcycle[30] ;
 wire \csr.mcycle[31] ;
 wire \csr.mcycle[3] ;
 wire \csr.mcycle[4] ;
 wire \csr.mcycle[5] ;
 wire \csr.mcycle[6] ;
 wire \csr.mcycle[7] ;
 wire \csr.mcycle[8] ;
 wire \csr.mcycle[9] ;
 wire \csr.meie ;
 wire \csr.minstret[0] ;
 wire \csr.minstret[10] ;
 wire \csr.minstret[11] ;
 wire \csr.minstret[12] ;
 wire \csr.minstret[13] ;
 wire \csr.minstret[14] ;
 wire \csr.minstret[15] ;
 wire \csr.minstret[16] ;
 wire \csr.minstret[17] ;
 wire \csr.minstret[18] ;
 wire \csr.minstret[19] ;
 wire \csr.minstret[1] ;
 wire \csr.minstret[20] ;
 wire \csr.minstret[21] ;
 wire \csr.minstret[22] ;
 wire \csr.minstret[23] ;
 wire \csr.minstret[24] ;
 wire \csr.minstret[25] ;
 wire \csr.minstret[26] ;
 wire \csr.minstret[27] ;
 wire \csr.minstret[28] ;
 wire \csr.minstret[29] ;
 wire \csr.minstret[2] ;
 wire \csr.minstret[30] ;
 wire \csr.minstret[31] ;
 wire \csr.minstret[3] ;
 wire \csr.minstret[4] ;
 wire \csr.minstret[5] ;
 wire \csr.minstret[6] ;
 wire \csr.minstret[7] ;
 wire \csr.minstret[8] ;
 wire \csr.minstret[9] ;
 wire \csr.mscratch[0] ;
 wire \csr.mscratch[10] ;
 wire \csr.mscratch[11] ;
 wire \csr.mscratch[12] ;
 wire \csr.mscratch[13] ;
 wire \csr.mscratch[14] ;
 wire \csr.mscratch[15] ;
 wire \csr.mscratch[16] ;
 wire \csr.mscratch[17] ;
 wire \csr.mscratch[18] ;
 wire \csr.mscratch[19] ;
 wire \csr.mscratch[1] ;
 wire \csr.mscratch[20] ;
 wire \csr.mscratch[21] ;
 wire \csr.mscratch[22] ;
 wire \csr.mscratch[23] ;
 wire \csr.mscratch[24] ;
 wire \csr.mscratch[25] ;
 wire \csr.mscratch[26] ;
 wire \csr.mscratch[27] ;
 wire \csr.mscratch[28] ;
 wire \csr.mscratch[29] ;
 wire \csr.mscratch[2] ;
 wire \csr.mscratch[30] ;
 wire \csr.mscratch[31] ;
 wire \csr.mscratch[3] ;
 wire \csr.mscratch[4] ;
 wire \csr.mscratch[5] ;
 wire \csr.mscratch[6] ;
 wire \csr.mscratch[7] ;
 wire \csr.mscratch[8] ;
 wire \csr.mscratch[9] ;
 wire \csr.msie ;
 wire \csr.msip ;
 wire \csr.mtie ;
 wire \csr.mtip ;
 wire \csr.pie ;
 wire \decode.control.io_funct3[0] ;
 wire \decode.control.io_funct3[1] ;
 wire \decode.control.io_funct3[2] ;
 wire \decode.control.io_funct7[0] ;
 wire \decode.control.io_funct7[1] ;
 wire \decode.control.io_funct7[2] ;
 wire \decode.control.io_funct7[3] ;
 wire \decode.control.io_funct7[4] ;
 wire \decode.control.io_funct7[5] ;
 wire \decode.control.io_funct7[6] ;
 wire \decode.control.io_opcode[0] ;
 wire \decode.control.io_opcode[1] ;
 wire \decode.control.io_opcode[2] ;
 wire \decode.control.io_opcode[3] ;
 wire \decode.control.io_opcode[4] ;
 wire \decode.control.io_opcode[5] ;
 wire \decode.control.io_opcode[6] ;
 wire \decode.csr_read_reg ;
 wire \decode.csr_write_reg ;
 wire \decode.exception_out_reg ;
 wire \decode.id_ex_aluop_reg[0] ;
 wire \decode.id_ex_aluop_reg[1] ;
 wire \decode.id_ex_aluop_reg[2] ;
 wire \decode.id_ex_aluop_reg[3] ;
 wire \decode.id_ex_ex_rd_reg[0] ;
 wire \decode.id_ex_ex_rd_reg[1] ;
 wire \decode.id_ex_ex_rd_reg[2] ;
 wire \decode.id_ex_ex_rd_reg[3] ;
 wire \decode.id_ex_ex_rd_reg[4] ;
 wire \decode.id_ex_ex_rs1_reg[0] ;
 wire \decode.id_ex_ex_rs1_reg[1] ;
 wire \decode.id_ex_ex_rs1_reg[2] ;
 wire \decode.id_ex_ex_rs1_reg[3] ;
 wire \decode.id_ex_ex_rs1_reg[4] ;
 wire \decode.id_ex_ex_use_rs1_reg ;
 wire \decode.id_ex_ex_use_rs2_reg ;
 wire \decode.id_ex_funct3_reg[0] ;
 wire \decode.id_ex_funct3_reg[1] ;
 wire \decode.id_ex_funct3_reg[2] ;
 wire \decode.id_ex_imm_reg[0] ;
 wire \decode.id_ex_imm_reg[10] ;
 wire \decode.id_ex_imm_reg[11] ;
 wire \decode.id_ex_imm_reg[12] ;
 wire \decode.id_ex_imm_reg[13] ;
 wire \decode.id_ex_imm_reg[14] ;
 wire \decode.id_ex_imm_reg[15] ;
 wire \decode.id_ex_imm_reg[16] ;
 wire \decode.id_ex_imm_reg[17] ;
 wire \decode.id_ex_imm_reg[18] ;
 wire \decode.id_ex_imm_reg[19] ;
 wire \decode.id_ex_imm_reg[1] ;
 wire \decode.id_ex_imm_reg[20] ;
 wire \decode.id_ex_imm_reg[21] ;
 wire \decode.id_ex_imm_reg[22] ;
 wire \decode.id_ex_imm_reg[23] ;
 wire \decode.id_ex_imm_reg[24] ;
 wire \decode.id_ex_imm_reg[25] ;
 wire \decode.id_ex_imm_reg[26] ;
 wire \decode.id_ex_imm_reg[27] ;
 wire \decode.id_ex_imm_reg[28] ;
 wire \decode.id_ex_imm_reg[29] ;
 wire \decode.id_ex_imm_reg[2] ;
 wire \decode.id_ex_imm_reg[30] ;
 wire \decode.id_ex_imm_reg[31] ;
 wire \decode.id_ex_imm_reg[3] ;
 wire \decode.id_ex_imm_reg[4] ;
 wire \decode.id_ex_imm_reg[5] ;
 wire \decode.id_ex_imm_reg[6] ;
 wire \decode.id_ex_imm_reg[7] ;
 wire \decode.id_ex_imm_reg[8] ;
 wire \decode.id_ex_imm_reg[9] ;
 wire \decode.id_ex_immsrc_reg ;
 wire \decode.id_ex_isbranch_reg ;
 wire \decode.id_ex_isjump_reg ;
 wire \decode.id_ex_islui_reg ;
 wire \decode.id_ex_memread_reg ;
 wire \decode.id_ex_memtoreg_reg[0] ;
 wire \decode.id_ex_memtoreg_reg[1] ;
 wire \decode.id_ex_memwrite_reg ;
 wire \decode.id_ex_pc_reg[0] ;
 wire \decode.id_ex_pc_reg[10] ;
 wire \decode.id_ex_pc_reg[11] ;
 wire \decode.id_ex_pc_reg[12] ;
 wire \decode.id_ex_pc_reg[13] ;
 wire \decode.id_ex_pc_reg[14] ;
 wire \decode.id_ex_pc_reg[15] ;
 wire \decode.id_ex_pc_reg[16] ;
 wire \decode.id_ex_pc_reg[17] ;
 wire \decode.id_ex_pc_reg[18] ;
 wire \decode.id_ex_pc_reg[19] ;
 wire \decode.id_ex_pc_reg[1] ;
 wire \decode.id_ex_pc_reg[20] ;
 wire \decode.id_ex_pc_reg[21] ;
 wire \decode.id_ex_pc_reg[22] ;
 wire \decode.id_ex_pc_reg[23] ;
 wire \decode.id_ex_pc_reg[24] ;
 wire \decode.id_ex_pc_reg[25] ;
 wire \decode.id_ex_pc_reg[26] ;
 wire \decode.id_ex_pc_reg[27] ;
 wire \decode.id_ex_pc_reg[28] ;
 wire \decode.id_ex_pc_reg[29] ;
 wire \decode.id_ex_pc_reg[2] ;
 wire \decode.id_ex_pc_reg[30] ;
 wire \decode.id_ex_pc_reg[31] ;
 wire \decode.id_ex_pc_reg[3] ;
 wire \decode.id_ex_pc_reg[4] ;
 wire \decode.id_ex_pc_reg[5] ;
 wire \decode.id_ex_pc_reg[6] ;
 wire \decode.id_ex_pc_reg[7] ;
 wire \decode.id_ex_pc_reg[8] ;
 wire \decode.id_ex_pc_reg[9] ;
 wire \decode.id_ex_pcsel_reg ;
 wire \decode.id_ex_rdsel_reg ;
 wire \decode.id_ex_regwrite_reg ;
 wire \decode.id_ex_rs1_data_reg[0] ;
 wire \decode.id_ex_rs1_data_reg[10] ;
 wire \decode.id_ex_rs1_data_reg[11] ;
 wire \decode.id_ex_rs1_data_reg[12] ;
 wire \decode.id_ex_rs1_data_reg[13] ;
 wire \decode.id_ex_rs1_data_reg[14] ;
 wire \decode.id_ex_rs1_data_reg[15] ;
 wire \decode.id_ex_rs1_data_reg[16] ;
 wire \decode.id_ex_rs1_data_reg[17] ;
 wire \decode.id_ex_rs1_data_reg[18] ;
 wire \decode.id_ex_rs1_data_reg[19] ;
 wire \decode.id_ex_rs1_data_reg[1] ;
 wire \decode.id_ex_rs1_data_reg[20] ;
 wire \decode.id_ex_rs1_data_reg[21] ;
 wire \decode.id_ex_rs1_data_reg[22] ;
 wire \decode.id_ex_rs1_data_reg[23] ;
 wire \decode.id_ex_rs1_data_reg[24] ;
 wire \decode.id_ex_rs1_data_reg[25] ;
 wire \decode.id_ex_rs1_data_reg[26] ;
 wire \decode.id_ex_rs1_data_reg[27] ;
 wire \decode.id_ex_rs1_data_reg[28] ;
 wire \decode.id_ex_rs1_data_reg[29] ;
 wire \decode.id_ex_rs1_data_reg[2] ;
 wire \decode.id_ex_rs1_data_reg[30] ;
 wire \decode.id_ex_rs1_data_reg[31] ;
 wire \decode.id_ex_rs1_data_reg[3] ;
 wire \decode.id_ex_rs1_data_reg[4] ;
 wire \decode.id_ex_rs1_data_reg[5] ;
 wire \decode.id_ex_rs1_data_reg[6] ;
 wire \decode.id_ex_rs1_data_reg[7] ;
 wire \decode.id_ex_rs1_data_reg[8] ;
 wire \decode.id_ex_rs1_data_reg[9] ;
 wire \decode.id_ex_rs2_data_reg[0] ;
 wire \decode.id_ex_rs2_data_reg[10] ;
 wire \decode.id_ex_rs2_data_reg[11] ;
 wire \decode.id_ex_rs2_data_reg[12] ;
 wire \decode.id_ex_rs2_data_reg[13] ;
 wire \decode.id_ex_rs2_data_reg[14] ;
 wire \decode.id_ex_rs2_data_reg[15] ;
 wire \decode.id_ex_rs2_data_reg[16] ;
 wire \decode.id_ex_rs2_data_reg[17] ;
 wire \decode.id_ex_rs2_data_reg[18] ;
 wire \decode.id_ex_rs2_data_reg[19] ;
 wire \decode.id_ex_rs2_data_reg[1] ;
 wire \decode.id_ex_rs2_data_reg[20] ;
 wire \decode.id_ex_rs2_data_reg[21] ;
 wire \decode.id_ex_rs2_data_reg[22] ;
 wire \decode.id_ex_rs2_data_reg[23] ;
 wire \decode.id_ex_rs2_data_reg[24] ;
 wire \decode.id_ex_rs2_data_reg[25] ;
 wire \decode.id_ex_rs2_data_reg[26] ;
 wire \decode.id_ex_rs2_data_reg[27] ;
 wire \decode.id_ex_rs2_data_reg[28] ;
 wire \decode.id_ex_rs2_data_reg[29] ;
 wire \decode.id_ex_rs2_data_reg[2] ;
 wire \decode.id_ex_rs2_data_reg[30] ;
 wire \decode.id_ex_rs2_data_reg[31] ;
 wire \decode.id_ex_rs2_data_reg[3] ;
 wire \decode.id_ex_rs2_data_reg[4] ;
 wire \decode.id_ex_rs2_data_reg[5] ;
 wire \decode.id_ex_rs2_data_reg[6] ;
 wire \decode.id_ex_rs2_data_reg[7] ;
 wire \decode.id_ex_rs2_data_reg[8] ;
 wire \decode.id_ex_rs2_data_reg[9] ;
 wire \decode.immGen._imm_T_10[0] ;
 wire \decode.immGen._imm_T_10[1] ;
 wire \decode.immGen._imm_T_10[2] ;
 wire \decode.immGen._imm_T_10[3] ;
 wire \decode.immGen._imm_T_10[4] ;
 wire \decode.immGen._imm_T_24[11] ;
 wire \decode.immGen._imm_T_24[15] ;
 wire \decode.immGen._imm_T_24[16] ;
 wire \decode.immGen._imm_T_24[17] ;
 wire \decode.immGen._imm_T_24[18] ;
 wire \decode.immGen._imm_T_24[19] ;
 wire \decode.immGen._imm_T_24[1] ;
 wire \decode.immGen._imm_T_24[2] ;
 wire \decode.immGen._imm_T_24[3] ;
 wire \decode.immGen._imm_T_24[4] ;
 wire \decode.io_id_pc[0] ;
 wire \decode.io_id_pc[10] ;
 wire \decode.io_id_pc[11] ;
 wire \decode.io_id_pc[12] ;
 wire \decode.io_id_pc[13] ;
 wire \decode.io_id_pc[14] ;
 wire \decode.io_id_pc[15] ;
 wire \decode.io_id_pc[16] ;
 wire \decode.io_id_pc[17] ;
 wire \decode.io_id_pc[18] ;
 wire \decode.io_id_pc[19] ;
 wire \decode.io_id_pc[1] ;
 wire \decode.io_id_pc[20] ;
 wire \decode.io_id_pc[21] ;
 wire \decode.io_id_pc[22] ;
 wire \decode.io_id_pc[23] ;
 wire \decode.io_id_pc[24] ;
 wire \decode.io_id_pc[25] ;
 wire \decode.io_id_pc[26] ;
 wire \decode.io_id_pc[27] ;
 wire \decode.io_id_pc[28] ;
 wire \decode.io_id_pc[29] ;
 wire \decode.io_id_pc[2] ;
 wire \decode.io_id_pc[30] ;
 wire \decode.io_id_pc[31] ;
 wire \decode.io_id_pc[3] ;
 wire \decode.io_id_pc[4] ;
 wire \decode.io_id_pc[5] ;
 wire \decode.io_id_pc[6] ;
 wire \decode.io_id_pc[7] ;
 wire \decode.io_id_pc[8] ;
 wire \decode.io_id_pc[9] ;
 wire \decode.io_mret_out ;
 wire \decode.io_wb_rd[0] ;
 wire \decode.io_wb_rd[1] ;
 wire \decode.io_wb_rd[2] ;
 wire \decode.io_wb_rd[3] ;
 wire \decode.io_wb_rd[4] ;
 wire \decode.io_wb_regwrite ;
 wire \decode.io_wfi_out ;
 wire \decode.regfile.registers_0[0] ;
 wire \decode.regfile.registers_0[10] ;
 wire \decode.regfile.registers_0[11] ;
 wire \decode.regfile.registers_0[12] ;
 wire \decode.regfile.registers_0[13] ;
 wire \decode.regfile.registers_0[14] ;
 wire \decode.regfile.registers_0[15] ;
 wire \decode.regfile.registers_0[16] ;
 wire \decode.regfile.registers_0[17] ;
 wire \decode.regfile.registers_0[18] ;
 wire \decode.regfile.registers_0[19] ;
 wire \decode.regfile.registers_0[1] ;
 wire \decode.regfile.registers_0[20] ;
 wire \decode.regfile.registers_0[21] ;
 wire \decode.regfile.registers_0[22] ;
 wire \decode.regfile.registers_0[23] ;
 wire \decode.regfile.registers_0[24] ;
 wire \decode.regfile.registers_0[25] ;
 wire \decode.regfile.registers_0[26] ;
 wire \decode.regfile.registers_0[27] ;
 wire \decode.regfile.registers_0[28] ;
 wire \decode.regfile.registers_0[29] ;
 wire \decode.regfile.registers_0[2] ;
 wire \decode.regfile.registers_0[30] ;
 wire \decode.regfile.registers_0[31] ;
 wire \decode.regfile.registers_0[3] ;
 wire \decode.regfile.registers_0[4] ;
 wire \decode.regfile.registers_0[5] ;
 wire \decode.regfile.registers_0[6] ;
 wire \decode.regfile.registers_0[7] ;
 wire \decode.regfile.registers_0[8] ;
 wire \decode.regfile.registers_0[9] ;
 wire \decode.regfile.registers_10[0] ;
 wire \decode.regfile.registers_10[10] ;
 wire \decode.regfile.registers_10[11] ;
 wire \decode.regfile.registers_10[12] ;
 wire \decode.regfile.registers_10[13] ;
 wire \decode.regfile.registers_10[14] ;
 wire \decode.regfile.registers_10[15] ;
 wire \decode.regfile.registers_10[16] ;
 wire \decode.regfile.registers_10[17] ;
 wire \decode.regfile.registers_10[18] ;
 wire \decode.regfile.registers_10[19] ;
 wire \decode.regfile.registers_10[1] ;
 wire \decode.regfile.registers_10[20] ;
 wire \decode.regfile.registers_10[21] ;
 wire \decode.regfile.registers_10[22] ;
 wire \decode.regfile.registers_10[23] ;
 wire \decode.regfile.registers_10[24] ;
 wire \decode.regfile.registers_10[25] ;
 wire \decode.regfile.registers_10[26] ;
 wire \decode.regfile.registers_10[27] ;
 wire \decode.regfile.registers_10[28] ;
 wire \decode.regfile.registers_10[29] ;
 wire \decode.regfile.registers_10[2] ;
 wire \decode.regfile.registers_10[30] ;
 wire \decode.regfile.registers_10[31] ;
 wire \decode.regfile.registers_10[3] ;
 wire \decode.regfile.registers_10[4] ;
 wire \decode.regfile.registers_10[5] ;
 wire \decode.regfile.registers_10[6] ;
 wire \decode.regfile.registers_10[7] ;
 wire \decode.regfile.registers_10[8] ;
 wire \decode.regfile.registers_10[9] ;
 wire \decode.regfile.registers_11[0] ;
 wire \decode.regfile.registers_11[10] ;
 wire \decode.regfile.registers_11[11] ;
 wire \decode.regfile.registers_11[12] ;
 wire \decode.regfile.registers_11[13] ;
 wire \decode.regfile.registers_11[14] ;
 wire \decode.regfile.registers_11[15] ;
 wire \decode.regfile.registers_11[16] ;
 wire \decode.regfile.registers_11[17] ;
 wire \decode.regfile.registers_11[18] ;
 wire \decode.regfile.registers_11[19] ;
 wire \decode.regfile.registers_11[1] ;
 wire \decode.regfile.registers_11[20] ;
 wire \decode.regfile.registers_11[21] ;
 wire \decode.regfile.registers_11[22] ;
 wire \decode.regfile.registers_11[23] ;
 wire \decode.regfile.registers_11[24] ;
 wire \decode.regfile.registers_11[25] ;
 wire \decode.regfile.registers_11[26] ;
 wire \decode.regfile.registers_11[27] ;
 wire \decode.regfile.registers_11[28] ;
 wire \decode.regfile.registers_11[29] ;
 wire \decode.regfile.registers_11[2] ;
 wire \decode.regfile.registers_11[30] ;
 wire \decode.regfile.registers_11[31] ;
 wire \decode.regfile.registers_11[3] ;
 wire \decode.regfile.registers_11[4] ;
 wire \decode.regfile.registers_11[5] ;
 wire \decode.regfile.registers_11[6] ;
 wire \decode.regfile.registers_11[7] ;
 wire \decode.regfile.registers_11[8] ;
 wire \decode.regfile.registers_11[9] ;
 wire \decode.regfile.registers_12[0] ;
 wire \decode.regfile.registers_12[10] ;
 wire \decode.regfile.registers_12[11] ;
 wire \decode.regfile.registers_12[12] ;
 wire \decode.regfile.registers_12[13] ;
 wire \decode.regfile.registers_12[14] ;
 wire \decode.regfile.registers_12[15] ;
 wire \decode.regfile.registers_12[16] ;
 wire \decode.regfile.registers_12[17] ;
 wire \decode.regfile.registers_12[18] ;
 wire \decode.regfile.registers_12[19] ;
 wire \decode.regfile.registers_12[1] ;
 wire \decode.regfile.registers_12[20] ;
 wire \decode.regfile.registers_12[21] ;
 wire \decode.regfile.registers_12[22] ;
 wire \decode.regfile.registers_12[23] ;
 wire \decode.regfile.registers_12[24] ;
 wire \decode.regfile.registers_12[25] ;
 wire \decode.regfile.registers_12[26] ;
 wire \decode.regfile.registers_12[27] ;
 wire \decode.regfile.registers_12[28] ;
 wire \decode.regfile.registers_12[29] ;
 wire \decode.regfile.registers_12[2] ;
 wire \decode.regfile.registers_12[30] ;
 wire \decode.regfile.registers_12[31] ;
 wire \decode.regfile.registers_12[3] ;
 wire \decode.regfile.registers_12[4] ;
 wire \decode.regfile.registers_12[5] ;
 wire \decode.regfile.registers_12[6] ;
 wire \decode.regfile.registers_12[7] ;
 wire \decode.regfile.registers_12[8] ;
 wire \decode.regfile.registers_12[9] ;
 wire \decode.regfile.registers_13[0] ;
 wire \decode.regfile.registers_13[10] ;
 wire \decode.regfile.registers_13[11] ;
 wire \decode.regfile.registers_13[12] ;
 wire \decode.regfile.registers_13[13] ;
 wire \decode.regfile.registers_13[14] ;
 wire \decode.regfile.registers_13[15] ;
 wire \decode.regfile.registers_13[16] ;
 wire \decode.regfile.registers_13[17] ;
 wire \decode.regfile.registers_13[18] ;
 wire \decode.regfile.registers_13[19] ;
 wire \decode.regfile.registers_13[1] ;
 wire \decode.regfile.registers_13[20] ;
 wire \decode.regfile.registers_13[21] ;
 wire \decode.regfile.registers_13[22] ;
 wire \decode.regfile.registers_13[23] ;
 wire \decode.regfile.registers_13[24] ;
 wire \decode.regfile.registers_13[25] ;
 wire \decode.regfile.registers_13[26] ;
 wire \decode.regfile.registers_13[27] ;
 wire \decode.regfile.registers_13[28] ;
 wire \decode.regfile.registers_13[29] ;
 wire \decode.regfile.registers_13[2] ;
 wire \decode.regfile.registers_13[30] ;
 wire \decode.regfile.registers_13[31] ;
 wire \decode.regfile.registers_13[3] ;
 wire \decode.regfile.registers_13[4] ;
 wire \decode.regfile.registers_13[5] ;
 wire \decode.regfile.registers_13[6] ;
 wire \decode.regfile.registers_13[7] ;
 wire \decode.regfile.registers_13[8] ;
 wire \decode.regfile.registers_13[9] ;
 wire \decode.regfile.registers_14[0] ;
 wire \decode.regfile.registers_14[10] ;
 wire \decode.regfile.registers_14[11] ;
 wire \decode.regfile.registers_14[12] ;
 wire \decode.regfile.registers_14[13] ;
 wire \decode.regfile.registers_14[14] ;
 wire \decode.regfile.registers_14[15] ;
 wire \decode.regfile.registers_14[16] ;
 wire \decode.regfile.registers_14[17] ;
 wire \decode.regfile.registers_14[18] ;
 wire \decode.regfile.registers_14[19] ;
 wire \decode.regfile.registers_14[1] ;
 wire \decode.regfile.registers_14[20] ;
 wire \decode.regfile.registers_14[21] ;
 wire \decode.regfile.registers_14[22] ;
 wire \decode.regfile.registers_14[23] ;
 wire \decode.regfile.registers_14[24] ;
 wire \decode.regfile.registers_14[25] ;
 wire \decode.regfile.registers_14[26] ;
 wire \decode.regfile.registers_14[27] ;
 wire \decode.regfile.registers_14[28] ;
 wire \decode.regfile.registers_14[29] ;
 wire \decode.regfile.registers_14[2] ;
 wire \decode.regfile.registers_14[30] ;
 wire \decode.regfile.registers_14[31] ;
 wire \decode.regfile.registers_14[3] ;
 wire \decode.regfile.registers_14[4] ;
 wire \decode.regfile.registers_14[5] ;
 wire \decode.regfile.registers_14[6] ;
 wire \decode.regfile.registers_14[7] ;
 wire \decode.regfile.registers_14[8] ;
 wire \decode.regfile.registers_14[9] ;
 wire \decode.regfile.registers_15[0] ;
 wire \decode.regfile.registers_15[10] ;
 wire \decode.regfile.registers_15[11] ;
 wire \decode.regfile.registers_15[12] ;
 wire \decode.regfile.registers_15[13] ;
 wire \decode.regfile.registers_15[14] ;
 wire \decode.regfile.registers_15[15] ;
 wire \decode.regfile.registers_15[16] ;
 wire \decode.regfile.registers_15[17] ;
 wire \decode.regfile.registers_15[18] ;
 wire \decode.regfile.registers_15[19] ;
 wire \decode.regfile.registers_15[1] ;
 wire \decode.regfile.registers_15[20] ;
 wire \decode.regfile.registers_15[21] ;
 wire \decode.regfile.registers_15[22] ;
 wire \decode.regfile.registers_15[23] ;
 wire \decode.regfile.registers_15[24] ;
 wire \decode.regfile.registers_15[25] ;
 wire \decode.regfile.registers_15[26] ;
 wire \decode.regfile.registers_15[27] ;
 wire \decode.regfile.registers_15[28] ;
 wire \decode.regfile.registers_15[29] ;
 wire \decode.regfile.registers_15[2] ;
 wire \decode.regfile.registers_15[30] ;
 wire \decode.regfile.registers_15[31] ;
 wire \decode.regfile.registers_15[3] ;
 wire \decode.regfile.registers_15[4] ;
 wire \decode.regfile.registers_15[5] ;
 wire \decode.regfile.registers_15[6] ;
 wire \decode.regfile.registers_15[7] ;
 wire \decode.regfile.registers_15[8] ;
 wire \decode.regfile.registers_15[9] ;
 wire \decode.regfile.registers_16[0] ;
 wire \decode.regfile.registers_16[10] ;
 wire \decode.regfile.registers_16[11] ;
 wire \decode.regfile.registers_16[12] ;
 wire \decode.regfile.registers_16[13] ;
 wire \decode.regfile.registers_16[14] ;
 wire \decode.regfile.registers_16[15] ;
 wire \decode.regfile.registers_16[16] ;
 wire \decode.regfile.registers_16[17] ;
 wire \decode.regfile.registers_16[18] ;
 wire \decode.regfile.registers_16[19] ;
 wire \decode.regfile.registers_16[1] ;
 wire \decode.regfile.registers_16[20] ;
 wire \decode.regfile.registers_16[21] ;
 wire \decode.regfile.registers_16[22] ;
 wire \decode.regfile.registers_16[23] ;
 wire \decode.regfile.registers_16[24] ;
 wire \decode.regfile.registers_16[25] ;
 wire \decode.regfile.registers_16[26] ;
 wire \decode.regfile.registers_16[27] ;
 wire \decode.regfile.registers_16[28] ;
 wire \decode.regfile.registers_16[29] ;
 wire \decode.regfile.registers_16[2] ;
 wire \decode.regfile.registers_16[30] ;
 wire \decode.regfile.registers_16[31] ;
 wire \decode.regfile.registers_16[3] ;
 wire \decode.regfile.registers_16[4] ;
 wire \decode.regfile.registers_16[5] ;
 wire \decode.regfile.registers_16[6] ;
 wire \decode.regfile.registers_16[7] ;
 wire \decode.regfile.registers_16[8] ;
 wire \decode.regfile.registers_16[9] ;
 wire \decode.regfile.registers_17[0] ;
 wire \decode.regfile.registers_17[10] ;
 wire \decode.regfile.registers_17[11] ;
 wire \decode.regfile.registers_17[12] ;
 wire \decode.regfile.registers_17[13] ;
 wire \decode.regfile.registers_17[14] ;
 wire \decode.regfile.registers_17[15] ;
 wire \decode.regfile.registers_17[16] ;
 wire \decode.regfile.registers_17[17] ;
 wire \decode.regfile.registers_17[18] ;
 wire \decode.regfile.registers_17[19] ;
 wire \decode.regfile.registers_17[1] ;
 wire \decode.regfile.registers_17[20] ;
 wire \decode.regfile.registers_17[21] ;
 wire \decode.regfile.registers_17[22] ;
 wire \decode.regfile.registers_17[23] ;
 wire \decode.regfile.registers_17[24] ;
 wire \decode.regfile.registers_17[25] ;
 wire \decode.regfile.registers_17[26] ;
 wire \decode.regfile.registers_17[27] ;
 wire \decode.regfile.registers_17[28] ;
 wire \decode.regfile.registers_17[29] ;
 wire \decode.regfile.registers_17[2] ;
 wire \decode.regfile.registers_17[30] ;
 wire \decode.regfile.registers_17[31] ;
 wire \decode.regfile.registers_17[3] ;
 wire \decode.regfile.registers_17[4] ;
 wire \decode.regfile.registers_17[5] ;
 wire \decode.regfile.registers_17[6] ;
 wire \decode.regfile.registers_17[7] ;
 wire \decode.regfile.registers_17[8] ;
 wire \decode.regfile.registers_17[9] ;
 wire \decode.regfile.registers_18[0] ;
 wire \decode.regfile.registers_18[10] ;
 wire \decode.regfile.registers_18[11] ;
 wire \decode.regfile.registers_18[12] ;
 wire \decode.regfile.registers_18[13] ;
 wire \decode.regfile.registers_18[14] ;
 wire \decode.regfile.registers_18[15] ;
 wire \decode.regfile.registers_18[16] ;
 wire \decode.regfile.registers_18[17] ;
 wire \decode.regfile.registers_18[18] ;
 wire \decode.regfile.registers_18[19] ;
 wire \decode.regfile.registers_18[1] ;
 wire \decode.regfile.registers_18[20] ;
 wire \decode.regfile.registers_18[21] ;
 wire \decode.regfile.registers_18[22] ;
 wire \decode.regfile.registers_18[23] ;
 wire \decode.regfile.registers_18[24] ;
 wire \decode.regfile.registers_18[25] ;
 wire \decode.regfile.registers_18[26] ;
 wire \decode.regfile.registers_18[27] ;
 wire \decode.regfile.registers_18[28] ;
 wire \decode.regfile.registers_18[29] ;
 wire \decode.regfile.registers_18[2] ;
 wire \decode.regfile.registers_18[30] ;
 wire \decode.regfile.registers_18[31] ;
 wire \decode.regfile.registers_18[3] ;
 wire \decode.regfile.registers_18[4] ;
 wire \decode.regfile.registers_18[5] ;
 wire \decode.regfile.registers_18[6] ;
 wire \decode.regfile.registers_18[7] ;
 wire \decode.regfile.registers_18[8] ;
 wire \decode.regfile.registers_18[9] ;
 wire \decode.regfile.registers_19[0] ;
 wire \decode.regfile.registers_19[10] ;
 wire \decode.regfile.registers_19[11] ;
 wire \decode.regfile.registers_19[12] ;
 wire \decode.regfile.registers_19[13] ;
 wire \decode.regfile.registers_19[14] ;
 wire \decode.regfile.registers_19[15] ;
 wire \decode.regfile.registers_19[16] ;
 wire \decode.regfile.registers_19[17] ;
 wire \decode.regfile.registers_19[18] ;
 wire \decode.regfile.registers_19[19] ;
 wire \decode.regfile.registers_19[1] ;
 wire \decode.regfile.registers_19[20] ;
 wire \decode.regfile.registers_19[21] ;
 wire \decode.regfile.registers_19[22] ;
 wire \decode.regfile.registers_19[23] ;
 wire \decode.regfile.registers_19[24] ;
 wire \decode.regfile.registers_19[25] ;
 wire \decode.regfile.registers_19[26] ;
 wire \decode.regfile.registers_19[27] ;
 wire \decode.regfile.registers_19[28] ;
 wire \decode.regfile.registers_19[29] ;
 wire \decode.regfile.registers_19[2] ;
 wire \decode.regfile.registers_19[30] ;
 wire \decode.regfile.registers_19[31] ;
 wire \decode.regfile.registers_19[3] ;
 wire \decode.regfile.registers_19[4] ;
 wire \decode.regfile.registers_19[5] ;
 wire \decode.regfile.registers_19[6] ;
 wire \decode.regfile.registers_19[7] ;
 wire \decode.regfile.registers_19[8] ;
 wire \decode.regfile.registers_19[9] ;
 wire \decode.regfile.registers_1[0] ;
 wire \decode.regfile.registers_1[10] ;
 wire \decode.regfile.registers_1[11] ;
 wire \decode.regfile.registers_1[12] ;
 wire \decode.regfile.registers_1[13] ;
 wire \decode.regfile.registers_1[14] ;
 wire \decode.regfile.registers_1[15] ;
 wire \decode.regfile.registers_1[16] ;
 wire \decode.regfile.registers_1[17] ;
 wire \decode.regfile.registers_1[18] ;
 wire \decode.regfile.registers_1[19] ;
 wire \decode.regfile.registers_1[1] ;
 wire \decode.regfile.registers_1[20] ;
 wire \decode.regfile.registers_1[21] ;
 wire \decode.regfile.registers_1[22] ;
 wire \decode.regfile.registers_1[23] ;
 wire \decode.regfile.registers_1[24] ;
 wire \decode.regfile.registers_1[25] ;
 wire \decode.regfile.registers_1[26] ;
 wire \decode.regfile.registers_1[27] ;
 wire \decode.regfile.registers_1[28] ;
 wire \decode.regfile.registers_1[29] ;
 wire \decode.regfile.registers_1[2] ;
 wire \decode.regfile.registers_1[30] ;
 wire \decode.regfile.registers_1[31] ;
 wire \decode.regfile.registers_1[3] ;
 wire \decode.regfile.registers_1[4] ;
 wire \decode.regfile.registers_1[5] ;
 wire \decode.regfile.registers_1[6] ;
 wire \decode.regfile.registers_1[7] ;
 wire \decode.regfile.registers_1[8] ;
 wire \decode.regfile.registers_1[9] ;
 wire \decode.regfile.registers_20[0] ;
 wire \decode.regfile.registers_20[10] ;
 wire \decode.regfile.registers_20[11] ;
 wire \decode.regfile.registers_20[12] ;
 wire \decode.regfile.registers_20[13] ;
 wire \decode.regfile.registers_20[14] ;
 wire \decode.regfile.registers_20[15] ;
 wire \decode.regfile.registers_20[16] ;
 wire \decode.regfile.registers_20[17] ;
 wire \decode.regfile.registers_20[18] ;
 wire \decode.regfile.registers_20[19] ;
 wire \decode.regfile.registers_20[1] ;
 wire \decode.regfile.registers_20[20] ;
 wire \decode.regfile.registers_20[21] ;
 wire \decode.regfile.registers_20[22] ;
 wire \decode.regfile.registers_20[23] ;
 wire \decode.regfile.registers_20[24] ;
 wire \decode.regfile.registers_20[25] ;
 wire \decode.regfile.registers_20[26] ;
 wire \decode.regfile.registers_20[27] ;
 wire \decode.regfile.registers_20[28] ;
 wire \decode.regfile.registers_20[29] ;
 wire \decode.regfile.registers_20[2] ;
 wire \decode.regfile.registers_20[30] ;
 wire \decode.regfile.registers_20[31] ;
 wire \decode.regfile.registers_20[3] ;
 wire \decode.regfile.registers_20[4] ;
 wire \decode.regfile.registers_20[5] ;
 wire \decode.regfile.registers_20[6] ;
 wire \decode.regfile.registers_20[7] ;
 wire \decode.regfile.registers_20[8] ;
 wire \decode.regfile.registers_20[9] ;
 wire \decode.regfile.registers_21[0] ;
 wire \decode.regfile.registers_21[10] ;
 wire \decode.regfile.registers_21[11] ;
 wire \decode.regfile.registers_21[12] ;
 wire \decode.regfile.registers_21[13] ;
 wire \decode.regfile.registers_21[14] ;
 wire \decode.regfile.registers_21[15] ;
 wire \decode.regfile.registers_21[16] ;
 wire \decode.regfile.registers_21[17] ;
 wire \decode.regfile.registers_21[18] ;
 wire \decode.regfile.registers_21[19] ;
 wire \decode.regfile.registers_21[1] ;
 wire \decode.regfile.registers_21[20] ;
 wire \decode.regfile.registers_21[21] ;
 wire \decode.regfile.registers_21[22] ;
 wire \decode.regfile.registers_21[23] ;
 wire \decode.regfile.registers_21[24] ;
 wire \decode.regfile.registers_21[25] ;
 wire \decode.regfile.registers_21[26] ;
 wire \decode.regfile.registers_21[27] ;
 wire \decode.regfile.registers_21[28] ;
 wire \decode.regfile.registers_21[29] ;
 wire \decode.regfile.registers_21[2] ;
 wire \decode.regfile.registers_21[30] ;
 wire \decode.regfile.registers_21[31] ;
 wire \decode.regfile.registers_21[3] ;
 wire \decode.regfile.registers_21[4] ;
 wire \decode.regfile.registers_21[5] ;
 wire \decode.regfile.registers_21[6] ;
 wire \decode.regfile.registers_21[7] ;
 wire \decode.regfile.registers_21[8] ;
 wire \decode.regfile.registers_21[9] ;
 wire \decode.regfile.registers_22[0] ;
 wire \decode.regfile.registers_22[10] ;
 wire \decode.regfile.registers_22[11] ;
 wire \decode.regfile.registers_22[12] ;
 wire \decode.regfile.registers_22[13] ;
 wire \decode.regfile.registers_22[14] ;
 wire \decode.regfile.registers_22[15] ;
 wire \decode.regfile.registers_22[16] ;
 wire \decode.regfile.registers_22[17] ;
 wire \decode.regfile.registers_22[18] ;
 wire \decode.regfile.registers_22[19] ;
 wire \decode.regfile.registers_22[1] ;
 wire \decode.regfile.registers_22[20] ;
 wire \decode.regfile.registers_22[21] ;
 wire \decode.regfile.registers_22[22] ;
 wire \decode.regfile.registers_22[23] ;
 wire \decode.regfile.registers_22[24] ;
 wire \decode.regfile.registers_22[25] ;
 wire \decode.regfile.registers_22[26] ;
 wire \decode.regfile.registers_22[27] ;
 wire \decode.regfile.registers_22[28] ;
 wire \decode.regfile.registers_22[29] ;
 wire \decode.regfile.registers_22[2] ;
 wire \decode.regfile.registers_22[30] ;
 wire \decode.regfile.registers_22[31] ;
 wire \decode.regfile.registers_22[3] ;
 wire \decode.regfile.registers_22[4] ;
 wire \decode.regfile.registers_22[5] ;
 wire \decode.regfile.registers_22[6] ;
 wire \decode.regfile.registers_22[7] ;
 wire \decode.regfile.registers_22[8] ;
 wire \decode.regfile.registers_22[9] ;
 wire \decode.regfile.registers_23[0] ;
 wire \decode.regfile.registers_23[10] ;
 wire \decode.regfile.registers_23[11] ;
 wire \decode.regfile.registers_23[12] ;
 wire \decode.regfile.registers_23[13] ;
 wire \decode.regfile.registers_23[14] ;
 wire \decode.regfile.registers_23[15] ;
 wire \decode.regfile.registers_23[16] ;
 wire \decode.regfile.registers_23[17] ;
 wire \decode.regfile.registers_23[18] ;
 wire \decode.regfile.registers_23[19] ;
 wire \decode.regfile.registers_23[1] ;
 wire \decode.regfile.registers_23[20] ;
 wire \decode.regfile.registers_23[21] ;
 wire \decode.regfile.registers_23[22] ;
 wire \decode.regfile.registers_23[23] ;
 wire \decode.regfile.registers_23[24] ;
 wire \decode.regfile.registers_23[25] ;
 wire \decode.regfile.registers_23[26] ;
 wire \decode.regfile.registers_23[27] ;
 wire \decode.regfile.registers_23[28] ;
 wire \decode.regfile.registers_23[29] ;
 wire \decode.regfile.registers_23[2] ;
 wire \decode.regfile.registers_23[30] ;
 wire \decode.regfile.registers_23[31] ;
 wire \decode.regfile.registers_23[3] ;
 wire \decode.regfile.registers_23[4] ;
 wire \decode.regfile.registers_23[5] ;
 wire \decode.regfile.registers_23[6] ;
 wire \decode.regfile.registers_23[7] ;
 wire \decode.regfile.registers_23[8] ;
 wire \decode.regfile.registers_23[9] ;
 wire \decode.regfile.registers_24[0] ;
 wire \decode.regfile.registers_24[10] ;
 wire \decode.regfile.registers_24[11] ;
 wire \decode.regfile.registers_24[12] ;
 wire \decode.regfile.registers_24[13] ;
 wire \decode.regfile.registers_24[14] ;
 wire \decode.regfile.registers_24[15] ;
 wire \decode.regfile.registers_24[16] ;
 wire \decode.regfile.registers_24[17] ;
 wire \decode.regfile.registers_24[18] ;
 wire \decode.regfile.registers_24[19] ;
 wire \decode.regfile.registers_24[1] ;
 wire \decode.regfile.registers_24[20] ;
 wire \decode.regfile.registers_24[21] ;
 wire \decode.regfile.registers_24[22] ;
 wire \decode.regfile.registers_24[23] ;
 wire \decode.regfile.registers_24[24] ;
 wire \decode.regfile.registers_24[25] ;
 wire \decode.regfile.registers_24[26] ;
 wire \decode.regfile.registers_24[27] ;
 wire \decode.regfile.registers_24[28] ;
 wire \decode.regfile.registers_24[29] ;
 wire \decode.regfile.registers_24[2] ;
 wire \decode.regfile.registers_24[30] ;
 wire \decode.regfile.registers_24[31] ;
 wire \decode.regfile.registers_24[3] ;
 wire \decode.regfile.registers_24[4] ;
 wire \decode.regfile.registers_24[5] ;
 wire \decode.regfile.registers_24[6] ;
 wire \decode.regfile.registers_24[7] ;
 wire \decode.regfile.registers_24[8] ;
 wire \decode.regfile.registers_24[9] ;
 wire \decode.regfile.registers_25[0] ;
 wire \decode.regfile.registers_25[10] ;
 wire \decode.regfile.registers_25[11] ;
 wire \decode.regfile.registers_25[12] ;
 wire \decode.regfile.registers_25[13] ;
 wire \decode.regfile.registers_25[14] ;
 wire \decode.regfile.registers_25[15] ;
 wire \decode.regfile.registers_25[16] ;
 wire \decode.regfile.registers_25[17] ;
 wire \decode.regfile.registers_25[18] ;
 wire \decode.regfile.registers_25[19] ;
 wire \decode.regfile.registers_25[1] ;
 wire \decode.regfile.registers_25[20] ;
 wire \decode.regfile.registers_25[21] ;
 wire \decode.regfile.registers_25[22] ;
 wire \decode.regfile.registers_25[23] ;
 wire \decode.regfile.registers_25[24] ;
 wire \decode.regfile.registers_25[25] ;
 wire \decode.regfile.registers_25[26] ;
 wire \decode.regfile.registers_25[27] ;
 wire \decode.regfile.registers_25[28] ;
 wire \decode.regfile.registers_25[29] ;
 wire \decode.regfile.registers_25[2] ;
 wire \decode.regfile.registers_25[30] ;
 wire \decode.regfile.registers_25[31] ;
 wire \decode.regfile.registers_25[3] ;
 wire \decode.regfile.registers_25[4] ;
 wire \decode.regfile.registers_25[5] ;
 wire \decode.regfile.registers_25[6] ;
 wire \decode.regfile.registers_25[7] ;
 wire \decode.regfile.registers_25[8] ;
 wire \decode.regfile.registers_25[9] ;
 wire \decode.regfile.registers_26[0] ;
 wire \decode.regfile.registers_26[10] ;
 wire \decode.regfile.registers_26[11] ;
 wire \decode.regfile.registers_26[12] ;
 wire \decode.regfile.registers_26[13] ;
 wire \decode.regfile.registers_26[14] ;
 wire \decode.regfile.registers_26[15] ;
 wire \decode.regfile.registers_26[16] ;
 wire \decode.regfile.registers_26[17] ;
 wire \decode.regfile.registers_26[18] ;
 wire \decode.regfile.registers_26[19] ;
 wire \decode.regfile.registers_26[1] ;
 wire \decode.regfile.registers_26[20] ;
 wire \decode.regfile.registers_26[21] ;
 wire \decode.regfile.registers_26[22] ;
 wire \decode.regfile.registers_26[23] ;
 wire \decode.regfile.registers_26[24] ;
 wire \decode.regfile.registers_26[25] ;
 wire \decode.regfile.registers_26[26] ;
 wire \decode.regfile.registers_26[27] ;
 wire \decode.regfile.registers_26[28] ;
 wire \decode.regfile.registers_26[29] ;
 wire \decode.regfile.registers_26[2] ;
 wire \decode.regfile.registers_26[30] ;
 wire \decode.regfile.registers_26[31] ;
 wire \decode.regfile.registers_26[3] ;
 wire \decode.regfile.registers_26[4] ;
 wire \decode.regfile.registers_26[5] ;
 wire \decode.regfile.registers_26[6] ;
 wire \decode.regfile.registers_26[7] ;
 wire \decode.regfile.registers_26[8] ;
 wire \decode.regfile.registers_26[9] ;
 wire \decode.regfile.registers_27[0] ;
 wire \decode.regfile.registers_27[10] ;
 wire \decode.regfile.registers_27[11] ;
 wire \decode.regfile.registers_27[12] ;
 wire \decode.regfile.registers_27[13] ;
 wire \decode.regfile.registers_27[14] ;
 wire \decode.regfile.registers_27[15] ;
 wire \decode.regfile.registers_27[16] ;
 wire \decode.regfile.registers_27[17] ;
 wire \decode.regfile.registers_27[18] ;
 wire \decode.regfile.registers_27[19] ;
 wire \decode.regfile.registers_27[1] ;
 wire \decode.regfile.registers_27[20] ;
 wire \decode.regfile.registers_27[21] ;
 wire \decode.regfile.registers_27[22] ;
 wire \decode.regfile.registers_27[23] ;
 wire \decode.regfile.registers_27[24] ;
 wire \decode.regfile.registers_27[25] ;
 wire \decode.regfile.registers_27[26] ;
 wire \decode.regfile.registers_27[27] ;
 wire \decode.regfile.registers_27[28] ;
 wire \decode.regfile.registers_27[29] ;
 wire \decode.regfile.registers_27[2] ;
 wire \decode.regfile.registers_27[30] ;
 wire \decode.regfile.registers_27[31] ;
 wire \decode.regfile.registers_27[3] ;
 wire \decode.regfile.registers_27[4] ;
 wire \decode.regfile.registers_27[5] ;
 wire \decode.regfile.registers_27[6] ;
 wire \decode.regfile.registers_27[7] ;
 wire \decode.regfile.registers_27[8] ;
 wire \decode.regfile.registers_27[9] ;
 wire \decode.regfile.registers_28[0] ;
 wire \decode.regfile.registers_28[10] ;
 wire \decode.regfile.registers_28[11] ;
 wire \decode.regfile.registers_28[12] ;
 wire \decode.regfile.registers_28[13] ;
 wire \decode.regfile.registers_28[14] ;
 wire \decode.regfile.registers_28[15] ;
 wire \decode.regfile.registers_28[16] ;
 wire \decode.regfile.registers_28[17] ;
 wire \decode.regfile.registers_28[18] ;
 wire \decode.regfile.registers_28[19] ;
 wire \decode.regfile.registers_28[1] ;
 wire \decode.regfile.registers_28[20] ;
 wire \decode.regfile.registers_28[21] ;
 wire \decode.regfile.registers_28[22] ;
 wire \decode.regfile.registers_28[23] ;
 wire \decode.regfile.registers_28[24] ;
 wire \decode.regfile.registers_28[25] ;
 wire \decode.regfile.registers_28[26] ;
 wire \decode.regfile.registers_28[27] ;
 wire \decode.regfile.registers_28[28] ;
 wire \decode.regfile.registers_28[29] ;
 wire \decode.regfile.registers_28[2] ;
 wire \decode.regfile.registers_28[30] ;
 wire \decode.regfile.registers_28[31] ;
 wire \decode.regfile.registers_28[3] ;
 wire \decode.regfile.registers_28[4] ;
 wire \decode.regfile.registers_28[5] ;
 wire \decode.regfile.registers_28[6] ;
 wire \decode.regfile.registers_28[7] ;
 wire \decode.regfile.registers_28[8] ;
 wire \decode.regfile.registers_28[9] ;
 wire \decode.regfile.registers_29[0] ;
 wire \decode.regfile.registers_29[10] ;
 wire \decode.regfile.registers_29[11] ;
 wire \decode.regfile.registers_29[12] ;
 wire \decode.regfile.registers_29[13] ;
 wire \decode.regfile.registers_29[14] ;
 wire \decode.regfile.registers_29[15] ;
 wire \decode.regfile.registers_29[16] ;
 wire \decode.regfile.registers_29[17] ;
 wire \decode.regfile.registers_29[18] ;
 wire \decode.regfile.registers_29[19] ;
 wire \decode.regfile.registers_29[1] ;
 wire \decode.regfile.registers_29[20] ;
 wire \decode.regfile.registers_29[21] ;
 wire \decode.regfile.registers_29[22] ;
 wire \decode.regfile.registers_29[23] ;
 wire \decode.regfile.registers_29[24] ;
 wire \decode.regfile.registers_29[25] ;
 wire \decode.regfile.registers_29[26] ;
 wire \decode.regfile.registers_29[27] ;
 wire \decode.regfile.registers_29[28] ;
 wire \decode.regfile.registers_29[29] ;
 wire \decode.regfile.registers_29[2] ;
 wire \decode.regfile.registers_29[30] ;
 wire \decode.regfile.registers_29[31] ;
 wire \decode.regfile.registers_29[3] ;
 wire \decode.regfile.registers_29[4] ;
 wire \decode.regfile.registers_29[5] ;
 wire \decode.regfile.registers_29[6] ;
 wire \decode.regfile.registers_29[7] ;
 wire \decode.regfile.registers_29[8] ;
 wire \decode.regfile.registers_29[9] ;
 wire \decode.regfile.registers_2[0] ;
 wire \decode.regfile.registers_2[10] ;
 wire \decode.regfile.registers_2[11] ;
 wire \decode.regfile.registers_2[12] ;
 wire \decode.regfile.registers_2[13] ;
 wire \decode.regfile.registers_2[14] ;
 wire \decode.regfile.registers_2[15] ;
 wire \decode.regfile.registers_2[16] ;
 wire \decode.regfile.registers_2[17] ;
 wire \decode.regfile.registers_2[18] ;
 wire \decode.regfile.registers_2[19] ;
 wire \decode.regfile.registers_2[1] ;
 wire \decode.regfile.registers_2[20] ;
 wire \decode.regfile.registers_2[21] ;
 wire \decode.regfile.registers_2[22] ;
 wire \decode.regfile.registers_2[23] ;
 wire \decode.regfile.registers_2[24] ;
 wire \decode.regfile.registers_2[25] ;
 wire \decode.regfile.registers_2[26] ;
 wire \decode.regfile.registers_2[27] ;
 wire \decode.regfile.registers_2[28] ;
 wire \decode.regfile.registers_2[29] ;
 wire \decode.regfile.registers_2[2] ;
 wire \decode.regfile.registers_2[30] ;
 wire \decode.regfile.registers_2[31] ;
 wire \decode.regfile.registers_2[3] ;
 wire \decode.regfile.registers_2[4] ;
 wire \decode.regfile.registers_2[5] ;
 wire \decode.regfile.registers_2[6] ;
 wire \decode.regfile.registers_2[7] ;
 wire \decode.regfile.registers_2[8] ;
 wire \decode.regfile.registers_2[9] ;
 wire \decode.regfile.registers_30[0] ;
 wire \decode.regfile.registers_30[10] ;
 wire \decode.regfile.registers_30[11] ;
 wire \decode.regfile.registers_30[12] ;
 wire \decode.regfile.registers_30[13] ;
 wire \decode.regfile.registers_30[14] ;
 wire \decode.regfile.registers_30[15] ;
 wire \decode.regfile.registers_30[16] ;
 wire \decode.regfile.registers_30[17] ;
 wire \decode.regfile.registers_30[18] ;
 wire \decode.regfile.registers_30[19] ;
 wire \decode.regfile.registers_30[1] ;
 wire \decode.regfile.registers_30[20] ;
 wire \decode.regfile.registers_30[21] ;
 wire \decode.regfile.registers_30[22] ;
 wire \decode.regfile.registers_30[23] ;
 wire \decode.regfile.registers_30[24] ;
 wire \decode.regfile.registers_30[25] ;
 wire \decode.regfile.registers_30[26] ;
 wire \decode.regfile.registers_30[27] ;
 wire \decode.regfile.registers_30[28] ;
 wire \decode.regfile.registers_30[29] ;
 wire \decode.regfile.registers_30[2] ;
 wire \decode.regfile.registers_30[30] ;
 wire \decode.regfile.registers_30[31] ;
 wire \decode.regfile.registers_30[3] ;
 wire \decode.regfile.registers_30[4] ;
 wire \decode.regfile.registers_30[5] ;
 wire \decode.regfile.registers_30[6] ;
 wire \decode.regfile.registers_30[7] ;
 wire \decode.regfile.registers_30[8] ;
 wire \decode.regfile.registers_30[9] ;
 wire \decode.regfile.registers_31[0] ;
 wire \decode.regfile.registers_31[10] ;
 wire \decode.regfile.registers_31[11] ;
 wire \decode.regfile.registers_31[12] ;
 wire \decode.regfile.registers_31[13] ;
 wire \decode.regfile.registers_31[14] ;
 wire \decode.regfile.registers_31[15] ;
 wire \decode.regfile.registers_31[16] ;
 wire \decode.regfile.registers_31[17] ;
 wire \decode.regfile.registers_31[18] ;
 wire \decode.regfile.registers_31[19] ;
 wire \decode.regfile.registers_31[1] ;
 wire \decode.regfile.registers_31[20] ;
 wire \decode.regfile.registers_31[21] ;
 wire \decode.regfile.registers_31[22] ;
 wire \decode.regfile.registers_31[23] ;
 wire \decode.regfile.registers_31[24] ;
 wire \decode.regfile.registers_31[25] ;
 wire \decode.regfile.registers_31[26] ;
 wire \decode.regfile.registers_31[27] ;
 wire \decode.regfile.registers_31[28] ;
 wire \decode.regfile.registers_31[29] ;
 wire \decode.regfile.registers_31[2] ;
 wire \decode.regfile.registers_31[30] ;
 wire \decode.regfile.registers_31[31] ;
 wire \decode.regfile.registers_31[3] ;
 wire \decode.regfile.registers_31[4] ;
 wire \decode.regfile.registers_31[5] ;
 wire \decode.regfile.registers_31[6] ;
 wire \decode.regfile.registers_31[7] ;
 wire \decode.regfile.registers_31[8] ;
 wire \decode.regfile.registers_31[9] ;
 wire \decode.regfile.registers_3[0] ;
 wire \decode.regfile.registers_3[10] ;
 wire \decode.regfile.registers_3[11] ;
 wire \decode.regfile.registers_3[12] ;
 wire \decode.regfile.registers_3[13] ;
 wire \decode.regfile.registers_3[14] ;
 wire \decode.regfile.registers_3[15] ;
 wire \decode.regfile.registers_3[16] ;
 wire \decode.regfile.registers_3[17] ;
 wire \decode.regfile.registers_3[18] ;
 wire \decode.regfile.registers_3[19] ;
 wire \decode.regfile.registers_3[1] ;
 wire \decode.regfile.registers_3[20] ;
 wire \decode.regfile.registers_3[21] ;
 wire \decode.regfile.registers_3[22] ;
 wire \decode.regfile.registers_3[23] ;
 wire \decode.regfile.registers_3[24] ;
 wire \decode.regfile.registers_3[25] ;
 wire \decode.regfile.registers_3[26] ;
 wire \decode.regfile.registers_3[27] ;
 wire \decode.regfile.registers_3[28] ;
 wire \decode.regfile.registers_3[29] ;
 wire \decode.regfile.registers_3[2] ;
 wire \decode.regfile.registers_3[30] ;
 wire \decode.regfile.registers_3[31] ;
 wire \decode.regfile.registers_3[3] ;
 wire \decode.regfile.registers_3[4] ;
 wire \decode.regfile.registers_3[5] ;
 wire \decode.regfile.registers_3[6] ;
 wire \decode.regfile.registers_3[7] ;
 wire \decode.regfile.registers_3[8] ;
 wire \decode.regfile.registers_3[9] ;
 wire \decode.regfile.registers_4[0] ;
 wire \decode.regfile.registers_4[10] ;
 wire \decode.regfile.registers_4[11] ;
 wire \decode.regfile.registers_4[12] ;
 wire \decode.regfile.registers_4[13] ;
 wire \decode.regfile.registers_4[14] ;
 wire \decode.regfile.registers_4[15] ;
 wire \decode.regfile.registers_4[16] ;
 wire \decode.regfile.registers_4[17] ;
 wire \decode.regfile.registers_4[18] ;
 wire \decode.regfile.registers_4[19] ;
 wire \decode.regfile.registers_4[1] ;
 wire \decode.regfile.registers_4[20] ;
 wire \decode.regfile.registers_4[21] ;
 wire \decode.regfile.registers_4[22] ;
 wire \decode.regfile.registers_4[23] ;
 wire \decode.regfile.registers_4[24] ;
 wire \decode.regfile.registers_4[25] ;
 wire \decode.regfile.registers_4[26] ;
 wire \decode.regfile.registers_4[27] ;
 wire \decode.regfile.registers_4[28] ;
 wire \decode.regfile.registers_4[29] ;
 wire \decode.regfile.registers_4[2] ;
 wire \decode.regfile.registers_4[30] ;
 wire \decode.regfile.registers_4[31] ;
 wire \decode.regfile.registers_4[3] ;
 wire \decode.regfile.registers_4[4] ;
 wire \decode.regfile.registers_4[5] ;
 wire \decode.regfile.registers_4[6] ;
 wire \decode.regfile.registers_4[7] ;
 wire \decode.regfile.registers_4[8] ;
 wire \decode.regfile.registers_4[9] ;
 wire \decode.regfile.registers_5[0] ;
 wire \decode.regfile.registers_5[10] ;
 wire \decode.regfile.registers_5[11] ;
 wire \decode.regfile.registers_5[12] ;
 wire \decode.regfile.registers_5[13] ;
 wire \decode.regfile.registers_5[14] ;
 wire \decode.regfile.registers_5[15] ;
 wire \decode.regfile.registers_5[16] ;
 wire \decode.regfile.registers_5[17] ;
 wire \decode.regfile.registers_5[18] ;
 wire \decode.regfile.registers_5[19] ;
 wire \decode.regfile.registers_5[1] ;
 wire \decode.regfile.registers_5[20] ;
 wire \decode.regfile.registers_5[21] ;
 wire \decode.regfile.registers_5[22] ;
 wire \decode.regfile.registers_5[23] ;
 wire \decode.regfile.registers_5[24] ;
 wire \decode.regfile.registers_5[25] ;
 wire \decode.regfile.registers_5[26] ;
 wire \decode.regfile.registers_5[27] ;
 wire \decode.regfile.registers_5[28] ;
 wire \decode.regfile.registers_5[29] ;
 wire \decode.regfile.registers_5[2] ;
 wire \decode.regfile.registers_5[30] ;
 wire \decode.regfile.registers_5[31] ;
 wire \decode.regfile.registers_5[3] ;
 wire \decode.regfile.registers_5[4] ;
 wire \decode.regfile.registers_5[5] ;
 wire \decode.regfile.registers_5[6] ;
 wire \decode.regfile.registers_5[7] ;
 wire \decode.regfile.registers_5[8] ;
 wire \decode.regfile.registers_5[9] ;
 wire \decode.regfile.registers_6[0] ;
 wire \decode.regfile.registers_6[10] ;
 wire \decode.regfile.registers_6[11] ;
 wire \decode.regfile.registers_6[12] ;
 wire \decode.regfile.registers_6[13] ;
 wire \decode.regfile.registers_6[14] ;
 wire \decode.regfile.registers_6[15] ;
 wire \decode.regfile.registers_6[16] ;
 wire \decode.regfile.registers_6[17] ;
 wire \decode.regfile.registers_6[18] ;
 wire \decode.regfile.registers_6[19] ;
 wire \decode.regfile.registers_6[1] ;
 wire \decode.regfile.registers_6[20] ;
 wire \decode.regfile.registers_6[21] ;
 wire \decode.regfile.registers_6[22] ;
 wire \decode.regfile.registers_6[23] ;
 wire \decode.regfile.registers_6[24] ;
 wire \decode.regfile.registers_6[25] ;
 wire \decode.regfile.registers_6[26] ;
 wire \decode.regfile.registers_6[27] ;
 wire \decode.regfile.registers_6[28] ;
 wire \decode.regfile.registers_6[29] ;
 wire \decode.regfile.registers_6[2] ;
 wire \decode.regfile.registers_6[30] ;
 wire \decode.regfile.registers_6[31] ;
 wire \decode.regfile.registers_6[3] ;
 wire \decode.regfile.registers_6[4] ;
 wire \decode.regfile.registers_6[5] ;
 wire \decode.regfile.registers_6[6] ;
 wire \decode.regfile.registers_6[7] ;
 wire \decode.regfile.registers_6[8] ;
 wire \decode.regfile.registers_6[9] ;
 wire \decode.regfile.registers_7[0] ;
 wire \decode.regfile.registers_7[10] ;
 wire \decode.regfile.registers_7[11] ;
 wire \decode.regfile.registers_7[12] ;
 wire \decode.regfile.registers_7[13] ;
 wire \decode.regfile.registers_7[14] ;
 wire \decode.regfile.registers_7[15] ;
 wire \decode.regfile.registers_7[16] ;
 wire \decode.regfile.registers_7[17] ;
 wire \decode.regfile.registers_7[18] ;
 wire \decode.regfile.registers_7[19] ;
 wire \decode.regfile.registers_7[1] ;
 wire \decode.regfile.registers_7[20] ;
 wire \decode.regfile.registers_7[21] ;
 wire \decode.regfile.registers_7[22] ;
 wire \decode.regfile.registers_7[23] ;
 wire \decode.regfile.registers_7[24] ;
 wire \decode.regfile.registers_7[25] ;
 wire \decode.regfile.registers_7[26] ;
 wire \decode.regfile.registers_7[27] ;
 wire \decode.regfile.registers_7[28] ;
 wire \decode.regfile.registers_7[29] ;
 wire \decode.regfile.registers_7[2] ;
 wire \decode.regfile.registers_7[30] ;
 wire \decode.regfile.registers_7[31] ;
 wire \decode.regfile.registers_7[3] ;
 wire \decode.regfile.registers_7[4] ;
 wire \decode.regfile.registers_7[5] ;
 wire \decode.regfile.registers_7[6] ;
 wire \decode.regfile.registers_7[7] ;
 wire \decode.regfile.registers_7[8] ;
 wire \decode.regfile.registers_7[9] ;
 wire \decode.regfile.registers_8[0] ;
 wire \decode.regfile.registers_8[10] ;
 wire \decode.regfile.registers_8[11] ;
 wire \decode.regfile.registers_8[12] ;
 wire \decode.regfile.registers_8[13] ;
 wire \decode.regfile.registers_8[14] ;
 wire \decode.regfile.registers_8[15] ;
 wire \decode.regfile.registers_8[16] ;
 wire \decode.regfile.registers_8[17] ;
 wire \decode.regfile.registers_8[18] ;
 wire \decode.regfile.registers_8[19] ;
 wire \decode.regfile.registers_8[1] ;
 wire \decode.regfile.registers_8[20] ;
 wire \decode.regfile.registers_8[21] ;
 wire \decode.regfile.registers_8[22] ;
 wire \decode.regfile.registers_8[23] ;
 wire \decode.regfile.registers_8[24] ;
 wire \decode.regfile.registers_8[25] ;
 wire \decode.regfile.registers_8[26] ;
 wire \decode.regfile.registers_8[27] ;
 wire \decode.regfile.registers_8[28] ;
 wire \decode.regfile.registers_8[29] ;
 wire \decode.regfile.registers_8[2] ;
 wire \decode.regfile.registers_8[30] ;
 wire \decode.regfile.registers_8[31] ;
 wire \decode.regfile.registers_8[3] ;
 wire \decode.regfile.registers_8[4] ;
 wire \decode.regfile.registers_8[5] ;
 wire \decode.regfile.registers_8[6] ;
 wire \decode.regfile.registers_8[7] ;
 wire \decode.regfile.registers_8[8] ;
 wire \decode.regfile.registers_8[9] ;
 wire \decode.regfile.registers_9[0] ;
 wire \decode.regfile.registers_9[10] ;
 wire \decode.regfile.registers_9[11] ;
 wire \decode.regfile.registers_9[12] ;
 wire \decode.regfile.registers_9[13] ;
 wire \decode.regfile.registers_9[14] ;
 wire \decode.regfile.registers_9[15] ;
 wire \decode.regfile.registers_9[16] ;
 wire \decode.regfile.registers_9[17] ;
 wire \decode.regfile.registers_9[18] ;
 wire \decode.regfile.registers_9[19] ;
 wire \decode.regfile.registers_9[1] ;
 wire \decode.regfile.registers_9[20] ;
 wire \decode.regfile.registers_9[21] ;
 wire \decode.regfile.registers_9[22] ;
 wire \decode.regfile.registers_9[23] ;
 wire \decode.regfile.registers_9[24] ;
 wire \decode.regfile.registers_9[25] ;
 wire \decode.regfile.registers_9[26] ;
 wire \decode.regfile.registers_9[27] ;
 wire \decode.regfile.registers_9[28] ;
 wire \decode.regfile.registers_9[29] ;
 wire \decode.regfile.registers_9[2] ;
 wire \decode.regfile.registers_9[30] ;
 wire \decode.regfile.registers_9[31] ;
 wire \decode.regfile.registers_9[3] ;
 wire \decode.regfile.registers_9[4] ;
 wire \decode.regfile.registers_9[5] ;
 wire \decode.regfile.registers_9[6] ;
 wire \decode.regfile.registers_9[7] ;
 wire \decode.regfile.registers_9[8] ;
 wire \decode.regfile.registers_9[9] ;
 wire \execute.csr_read_data_out_reg[0] ;
 wire \execute.csr_read_data_out_reg[10] ;
 wire \execute.csr_read_data_out_reg[11] ;
 wire \execute.csr_read_data_out_reg[12] ;
 wire \execute.csr_read_data_out_reg[13] ;
 wire \execute.csr_read_data_out_reg[14] ;
 wire \execute.csr_read_data_out_reg[15] ;
 wire \execute.csr_read_data_out_reg[16] ;
 wire \execute.csr_read_data_out_reg[17] ;
 wire \execute.csr_read_data_out_reg[18] ;
 wire \execute.csr_read_data_out_reg[19] ;
 wire \execute.csr_read_data_out_reg[1] ;
 wire \execute.csr_read_data_out_reg[20] ;
 wire \execute.csr_read_data_out_reg[21] ;
 wire \execute.csr_read_data_out_reg[22] ;
 wire \execute.csr_read_data_out_reg[23] ;
 wire \execute.csr_read_data_out_reg[24] ;
 wire \execute.csr_read_data_out_reg[25] ;
 wire \execute.csr_read_data_out_reg[26] ;
 wire \execute.csr_read_data_out_reg[27] ;
 wire \execute.csr_read_data_out_reg[28] ;
 wire \execute.csr_read_data_out_reg[29] ;
 wire \execute.csr_read_data_out_reg[2] ;
 wire \execute.csr_read_data_out_reg[30] ;
 wire \execute.csr_read_data_out_reg[31] ;
 wire \execute.csr_read_data_out_reg[3] ;
 wire \execute.csr_read_data_out_reg[4] ;
 wire \execute.csr_read_data_out_reg[5] ;
 wire \execute.csr_read_data_out_reg[6] ;
 wire \execute.csr_read_data_out_reg[7] ;
 wire \execute.csr_read_data_out_reg[8] ;
 wire \execute.csr_read_data_out_reg[9] ;
 wire \execute.csr_write_address_out_reg[0] ;
 wire \execute.csr_write_address_out_reg[10] ;
 wire \execute.csr_write_address_out_reg[11] ;
 wire \execute.csr_write_address_out_reg[1] ;
 wire \execute.csr_write_address_out_reg[2] ;
 wire \execute.csr_write_address_out_reg[3] ;
 wire \execute.csr_write_address_out_reg[4] ;
 wire \execute.csr_write_address_out_reg[5] ;
 wire \execute.csr_write_address_out_reg[6] ;
 wire \execute.csr_write_address_out_reg[7] ;
 wire \execute.csr_write_address_out_reg[8] ;
 wire \execute.csr_write_address_out_reg[9] ;
 wire \execute.csr_write_data_out_reg[0] ;
 wire \execute.csr_write_data_out_reg[10] ;
 wire \execute.csr_write_data_out_reg[11] ;
 wire \execute.csr_write_data_out_reg[12] ;
 wire \execute.csr_write_data_out_reg[13] ;
 wire \execute.csr_write_data_out_reg[14] ;
 wire \execute.csr_write_data_out_reg[15] ;
 wire \execute.csr_write_data_out_reg[16] ;
 wire \execute.csr_write_data_out_reg[17] ;
 wire \execute.csr_write_data_out_reg[18] ;
 wire \execute.csr_write_data_out_reg[19] ;
 wire \execute.csr_write_data_out_reg[1] ;
 wire \execute.csr_write_data_out_reg[20] ;
 wire \execute.csr_write_data_out_reg[21] ;
 wire \execute.csr_write_data_out_reg[22] ;
 wire \execute.csr_write_data_out_reg[23] ;
 wire \execute.csr_write_data_out_reg[24] ;
 wire \execute.csr_write_data_out_reg[25] ;
 wire \execute.csr_write_data_out_reg[26] ;
 wire \execute.csr_write_data_out_reg[27] ;
 wire \execute.csr_write_data_out_reg[28] ;
 wire \execute.csr_write_data_out_reg[29] ;
 wire \execute.csr_write_data_out_reg[2] ;
 wire \execute.csr_write_data_out_reg[30] ;
 wire \execute.csr_write_data_out_reg[31] ;
 wire \execute.csr_write_data_out_reg[3] ;
 wire \execute.csr_write_data_out_reg[4] ;
 wire \execute.csr_write_data_out_reg[5] ;
 wire \execute.csr_write_data_out_reg[6] ;
 wire \execute.csr_write_data_out_reg[7] ;
 wire \execute.csr_write_data_out_reg[8] ;
 wire \execute.csr_write_data_out_reg[9] ;
 wire \execute.csr_write_enable_out_reg ;
 wire \execute.exception_out_reg ;
 wire \execute.io_mem_isbranch ;
 wire \execute.io_mem_isjump ;
 wire \execute.io_mem_memtoreg[0] ;
 wire \execute.io_mem_memtoreg[1] ;
 wire \execute.io_mem_memwrite ;
 wire \execute.io_mem_rd[0] ;
 wire \execute.io_mem_rd[1] ;
 wire \execute.io_mem_rd[2] ;
 wire \execute.io_mem_rd[3] ;
 wire \execute.io_mem_rd[4] ;
 wire \execute.io_mem_regwrite ;
 wire \execute.io_mem_zero ;
 wire \execute.io_mret_out ;
 wire \execute.io_reg_pc[0] ;
 wire \execute.io_reg_pc[10] ;
 wire \execute.io_reg_pc[11] ;
 wire \execute.io_reg_pc[12] ;
 wire \execute.io_reg_pc[13] ;
 wire \execute.io_reg_pc[14] ;
 wire \execute.io_reg_pc[15] ;
 wire \execute.io_reg_pc[16] ;
 wire \execute.io_reg_pc[17] ;
 wire \execute.io_reg_pc[18] ;
 wire \execute.io_reg_pc[19] ;
 wire \execute.io_reg_pc[1] ;
 wire \execute.io_reg_pc[20] ;
 wire \execute.io_reg_pc[21] ;
 wire \execute.io_reg_pc[22] ;
 wire \execute.io_reg_pc[23] ;
 wire \execute.io_reg_pc[24] ;
 wire \execute.io_reg_pc[25] ;
 wire \execute.io_reg_pc[26] ;
 wire \execute.io_reg_pc[27] ;
 wire \execute.io_reg_pc[28] ;
 wire \execute.io_reg_pc[29] ;
 wire \execute.io_reg_pc[2] ;
 wire \execute.io_reg_pc[30] ;
 wire \execute.io_reg_pc[31] ;
 wire \execute.io_reg_pc[3] ;
 wire \execute.io_reg_pc[4] ;
 wire \execute.io_reg_pc[5] ;
 wire \execute.io_reg_pc[6] ;
 wire \execute.io_reg_pc[7] ;
 wire \execute.io_reg_pc[8] ;
 wire \execute.io_reg_pc[9] ;
 wire \execute.io_target_pc[0] ;
 wire \execute.io_target_pc[10] ;
 wire \execute.io_target_pc[11] ;
 wire \execute.io_target_pc[12] ;
 wire \execute.io_target_pc[13] ;
 wire \execute.io_target_pc[14] ;
 wire \execute.io_target_pc[15] ;
 wire \execute.io_target_pc[16] ;
 wire \execute.io_target_pc[17] ;
 wire \execute.io_target_pc[18] ;
 wire \execute.io_target_pc[19] ;
 wire \execute.io_target_pc[1] ;
 wire \execute.io_target_pc[20] ;
 wire \execute.io_target_pc[21] ;
 wire \execute.io_target_pc[22] ;
 wire \execute.io_target_pc[23] ;
 wire \execute.io_target_pc[24] ;
 wire \execute.io_target_pc[25] ;
 wire \execute.io_target_pc[26] ;
 wire \execute.io_target_pc[27] ;
 wire \execute.io_target_pc[28] ;
 wire \execute.io_target_pc[29] ;
 wire \execute.io_target_pc[2] ;
 wire \execute.io_target_pc[30] ;
 wire \execute.io_target_pc[31] ;
 wire \execute.io_target_pc[3] ;
 wire \execute.io_target_pc[4] ;
 wire \execute.io_target_pc[5] ;
 wire \execute.io_target_pc[6] ;
 wire \execute.io_target_pc[7] ;
 wire \execute.io_target_pc[8] ;
 wire \execute.io_target_pc[9] ;
 wire \execute.io_wfi_out ;
 wire \fetch.bht.bhtTable_tag[0][0] ;
 wire \fetch.bht.bhtTable_tag[0][10] ;
 wire \fetch.bht.bhtTable_tag[0][11] ;
 wire \fetch.bht.bhtTable_tag[0][12] ;
 wire \fetch.bht.bhtTable_tag[0][13] ;
 wire \fetch.bht.bhtTable_tag[0][14] ;
 wire \fetch.bht.bhtTable_tag[0][15] ;
 wire \fetch.bht.bhtTable_tag[0][16] ;
 wire \fetch.bht.bhtTable_tag[0][17] ;
 wire \fetch.bht.bhtTable_tag[0][18] ;
 wire \fetch.bht.bhtTable_tag[0][19] ;
 wire \fetch.bht.bhtTable_tag[0][1] ;
 wire \fetch.bht.bhtTable_tag[0][20] ;
 wire \fetch.bht.bhtTable_tag[0][21] ;
 wire \fetch.bht.bhtTable_tag[0][22] ;
 wire \fetch.bht.bhtTable_tag[0][23] ;
 wire \fetch.bht.bhtTable_tag[0][24] ;
 wire \fetch.bht.bhtTable_tag[0][25] ;
 wire \fetch.bht.bhtTable_tag[0][2] ;
 wire \fetch.bht.bhtTable_tag[0][3] ;
 wire \fetch.bht.bhtTable_tag[0][4] ;
 wire \fetch.bht.bhtTable_tag[0][5] ;
 wire \fetch.bht.bhtTable_tag[0][6] ;
 wire \fetch.bht.bhtTable_tag[0][7] ;
 wire \fetch.bht.bhtTable_tag[0][8] ;
 wire \fetch.bht.bhtTable_tag[0][9] ;
 wire \fetch.bht.bhtTable_tag[10][0] ;
 wire \fetch.bht.bhtTable_tag[10][10] ;
 wire \fetch.bht.bhtTable_tag[10][11] ;
 wire \fetch.bht.bhtTable_tag[10][12] ;
 wire \fetch.bht.bhtTable_tag[10][13] ;
 wire \fetch.bht.bhtTable_tag[10][14] ;
 wire \fetch.bht.bhtTable_tag[10][15] ;
 wire \fetch.bht.bhtTable_tag[10][16] ;
 wire \fetch.bht.bhtTable_tag[10][17] ;
 wire \fetch.bht.bhtTable_tag[10][18] ;
 wire \fetch.bht.bhtTable_tag[10][19] ;
 wire \fetch.bht.bhtTable_tag[10][1] ;
 wire \fetch.bht.bhtTable_tag[10][20] ;
 wire \fetch.bht.bhtTable_tag[10][21] ;
 wire \fetch.bht.bhtTable_tag[10][22] ;
 wire \fetch.bht.bhtTable_tag[10][23] ;
 wire \fetch.bht.bhtTable_tag[10][24] ;
 wire \fetch.bht.bhtTable_tag[10][25] ;
 wire \fetch.bht.bhtTable_tag[10][2] ;
 wire \fetch.bht.bhtTable_tag[10][3] ;
 wire \fetch.bht.bhtTable_tag[10][4] ;
 wire \fetch.bht.bhtTable_tag[10][5] ;
 wire \fetch.bht.bhtTable_tag[10][6] ;
 wire \fetch.bht.bhtTable_tag[10][7] ;
 wire \fetch.bht.bhtTable_tag[10][8] ;
 wire \fetch.bht.bhtTable_tag[10][9] ;
 wire \fetch.bht.bhtTable_tag[11][0] ;
 wire \fetch.bht.bhtTable_tag[11][10] ;
 wire \fetch.bht.bhtTable_tag[11][11] ;
 wire \fetch.bht.bhtTable_tag[11][12] ;
 wire \fetch.bht.bhtTable_tag[11][13] ;
 wire \fetch.bht.bhtTable_tag[11][14] ;
 wire \fetch.bht.bhtTable_tag[11][15] ;
 wire \fetch.bht.bhtTable_tag[11][16] ;
 wire \fetch.bht.bhtTable_tag[11][17] ;
 wire \fetch.bht.bhtTable_tag[11][18] ;
 wire \fetch.bht.bhtTable_tag[11][19] ;
 wire \fetch.bht.bhtTable_tag[11][1] ;
 wire \fetch.bht.bhtTable_tag[11][20] ;
 wire \fetch.bht.bhtTable_tag[11][21] ;
 wire \fetch.bht.bhtTable_tag[11][22] ;
 wire \fetch.bht.bhtTable_tag[11][23] ;
 wire \fetch.bht.bhtTable_tag[11][24] ;
 wire \fetch.bht.bhtTable_tag[11][25] ;
 wire \fetch.bht.bhtTable_tag[11][2] ;
 wire \fetch.bht.bhtTable_tag[11][3] ;
 wire \fetch.bht.bhtTable_tag[11][4] ;
 wire \fetch.bht.bhtTable_tag[11][5] ;
 wire \fetch.bht.bhtTable_tag[11][6] ;
 wire \fetch.bht.bhtTable_tag[11][7] ;
 wire \fetch.bht.bhtTable_tag[11][8] ;
 wire \fetch.bht.bhtTable_tag[11][9] ;
 wire \fetch.bht.bhtTable_tag[12][0] ;
 wire \fetch.bht.bhtTable_tag[12][10] ;
 wire \fetch.bht.bhtTable_tag[12][11] ;
 wire \fetch.bht.bhtTable_tag[12][12] ;
 wire \fetch.bht.bhtTable_tag[12][13] ;
 wire \fetch.bht.bhtTable_tag[12][14] ;
 wire \fetch.bht.bhtTable_tag[12][15] ;
 wire \fetch.bht.bhtTable_tag[12][16] ;
 wire \fetch.bht.bhtTable_tag[12][17] ;
 wire \fetch.bht.bhtTable_tag[12][18] ;
 wire \fetch.bht.bhtTable_tag[12][19] ;
 wire \fetch.bht.bhtTable_tag[12][1] ;
 wire \fetch.bht.bhtTable_tag[12][20] ;
 wire \fetch.bht.bhtTable_tag[12][21] ;
 wire \fetch.bht.bhtTable_tag[12][22] ;
 wire \fetch.bht.bhtTable_tag[12][23] ;
 wire \fetch.bht.bhtTable_tag[12][24] ;
 wire \fetch.bht.bhtTable_tag[12][25] ;
 wire \fetch.bht.bhtTable_tag[12][2] ;
 wire \fetch.bht.bhtTable_tag[12][3] ;
 wire \fetch.bht.bhtTable_tag[12][4] ;
 wire \fetch.bht.bhtTable_tag[12][5] ;
 wire \fetch.bht.bhtTable_tag[12][6] ;
 wire \fetch.bht.bhtTable_tag[12][7] ;
 wire \fetch.bht.bhtTable_tag[12][8] ;
 wire \fetch.bht.bhtTable_tag[12][9] ;
 wire \fetch.bht.bhtTable_tag[13][0] ;
 wire \fetch.bht.bhtTable_tag[13][10] ;
 wire \fetch.bht.bhtTable_tag[13][11] ;
 wire \fetch.bht.bhtTable_tag[13][12] ;
 wire \fetch.bht.bhtTable_tag[13][13] ;
 wire \fetch.bht.bhtTable_tag[13][14] ;
 wire \fetch.bht.bhtTable_tag[13][15] ;
 wire \fetch.bht.bhtTable_tag[13][16] ;
 wire \fetch.bht.bhtTable_tag[13][17] ;
 wire \fetch.bht.bhtTable_tag[13][18] ;
 wire \fetch.bht.bhtTable_tag[13][19] ;
 wire \fetch.bht.bhtTable_tag[13][1] ;
 wire \fetch.bht.bhtTable_tag[13][20] ;
 wire \fetch.bht.bhtTable_tag[13][21] ;
 wire \fetch.bht.bhtTable_tag[13][22] ;
 wire \fetch.bht.bhtTable_tag[13][23] ;
 wire \fetch.bht.bhtTable_tag[13][24] ;
 wire \fetch.bht.bhtTable_tag[13][25] ;
 wire \fetch.bht.bhtTable_tag[13][2] ;
 wire \fetch.bht.bhtTable_tag[13][3] ;
 wire \fetch.bht.bhtTable_tag[13][4] ;
 wire \fetch.bht.bhtTable_tag[13][5] ;
 wire \fetch.bht.bhtTable_tag[13][6] ;
 wire \fetch.bht.bhtTable_tag[13][7] ;
 wire \fetch.bht.bhtTable_tag[13][8] ;
 wire \fetch.bht.bhtTable_tag[13][9] ;
 wire \fetch.bht.bhtTable_tag[14][0] ;
 wire \fetch.bht.bhtTable_tag[14][10] ;
 wire \fetch.bht.bhtTable_tag[14][11] ;
 wire \fetch.bht.bhtTable_tag[14][12] ;
 wire \fetch.bht.bhtTable_tag[14][13] ;
 wire \fetch.bht.bhtTable_tag[14][14] ;
 wire \fetch.bht.bhtTable_tag[14][15] ;
 wire \fetch.bht.bhtTable_tag[14][16] ;
 wire \fetch.bht.bhtTable_tag[14][17] ;
 wire \fetch.bht.bhtTable_tag[14][18] ;
 wire \fetch.bht.bhtTable_tag[14][19] ;
 wire \fetch.bht.bhtTable_tag[14][1] ;
 wire \fetch.bht.bhtTable_tag[14][20] ;
 wire \fetch.bht.bhtTable_tag[14][21] ;
 wire \fetch.bht.bhtTable_tag[14][22] ;
 wire \fetch.bht.bhtTable_tag[14][23] ;
 wire \fetch.bht.bhtTable_tag[14][24] ;
 wire \fetch.bht.bhtTable_tag[14][25] ;
 wire \fetch.bht.bhtTable_tag[14][2] ;
 wire \fetch.bht.bhtTable_tag[14][3] ;
 wire \fetch.bht.bhtTable_tag[14][4] ;
 wire \fetch.bht.bhtTable_tag[14][5] ;
 wire \fetch.bht.bhtTable_tag[14][6] ;
 wire \fetch.bht.bhtTable_tag[14][7] ;
 wire \fetch.bht.bhtTable_tag[14][8] ;
 wire \fetch.bht.bhtTable_tag[14][9] ;
 wire \fetch.bht.bhtTable_tag[15][0] ;
 wire \fetch.bht.bhtTable_tag[15][10] ;
 wire \fetch.bht.bhtTable_tag[15][11] ;
 wire \fetch.bht.bhtTable_tag[15][12] ;
 wire \fetch.bht.bhtTable_tag[15][13] ;
 wire \fetch.bht.bhtTable_tag[15][14] ;
 wire \fetch.bht.bhtTable_tag[15][15] ;
 wire \fetch.bht.bhtTable_tag[15][16] ;
 wire \fetch.bht.bhtTable_tag[15][17] ;
 wire \fetch.bht.bhtTable_tag[15][18] ;
 wire \fetch.bht.bhtTable_tag[15][19] ;
 wire \fetch.bht.bhtTable_tag[15][1] ;
 wire \fetch.bht.bhtTable_tag[15][20] ;
 wire \fetch.bht.bhtTable_tag[15][21] ;
 wire \fetch.bht.bhtTable_tag[15][22] ;
 wire \fetch.bht.bhtTable_tag[15][23] ;
 wire \fetch.bht.bhtTable_tag[15][24] ;
 wire \fetch.bht.bhtTable_tag[15][25] ;
 wire \fetch.bht.bhtTable_tag[15][2] ;
 wire \fetch.bht.bhtTable_tag[15][3] ;
 wire \fetch.bht.bhtTable_tag[15][4] ;
 wire \fetch.bht.bhtTable_tag[15][5] ;
 wire \fetch.bht.bhtTable_tag[15][6] ;
 wire \fetch.bht.bhtTable_tag[15][7] ;
 wire \fetch.bht.bhtTable_tag[15][8] ;
 wire \fetch.bht.bhtTable_tag[15][9] ;
 wire \fetch.bht.bhtTable_tag[1][0] ;
 wire \fetch.bht.bhtTable_tag[1][10] ;
 wire \fetch.bht.bhtTable_tag[1][11] ;
 wire \fetch.bht.bhtTable_tag[1][12] ;
 wire \fetch.bht.bhtTable_tag[1][13] ;
 wire \fetch.bht.bhtTable_tag[1][14] ;
 wire \fetch.bht.bhtTable_tag[1][15] ;
 wire \fetch.bht.bhtTable_tag[1][16] ;
 wire \fetch.bht.bhtTable_tag[1][17] ;
 wire \fetch.bht.bhtTable_tag[1][18] ;
 wire \fetch.bht.bhtTable_tag[1][19] ;
 wire \fetch.bht.bhtTable_tag[1][1] ;
 wire \fetch.bht.bhtTable_tag[1][20] ;
 wire \fetch.bht.bhtTable_tag[1][21] ;
 wire \fetch.bht.bhtTable_tag[1][22] ;
 wire \fetch.bht.bhtTable_tag[1][23] ;
 wire \fetch.bht.bhtTable_tag[1][24] ;
 wire \fetch.bht.bhtTable_tag[1][25] ;
 wire \fetch.bht.bhtTable_tag[1][2] ;
 wire \fetch.bht.bhtTable_tag[1][3] ;
 wire \fetch.bht.bhtTable_tag[1][4] ;
 wire \fetch.bht.bhtTable_tag[1][5] ;
 wire \fetch.bht.bhtTable_tag[1][6] ;
 wire \fetch.bht.bhtTable_tag[1][7] ;
 wire \fetch.bht.bhtTable_tag[1][8] ;
 wire \fetch.bht.bhtTable_tag[1][9] ;
 wire \fetch.bht.bhtTable_tag[2][0] ;
 wire \fetch.bht.bhtTable_tag[2][10] ;
 wire \fetch.bht.bhtTable_tag[2][11] ;
 wire \fetch.bht.bhtTable_tag[2][12] ;
 wire \fetch.bht.bhtTable_tag[2][13] ;
 wire \fetch.bht.bhtTable_tag[2][14] ;
 wire \fetch.bht.bhtTable_tag[2][15] ;
 wire \fetch.bht.bhtTable_tag[2][16] ;
 wire \fetch.bht.bhtTable_tag[2][17] ;
 wire \fetch.bht.bhtTable_tag[2][18] ;
 wire \fetch.bht.bhtTable_tag[2][19] ;
 wire \fetch.bht.bhtTable_tag[2][1] ;
 wire \fetch.bht.bhtTable_tag[2][20] ;
 wire \fetch.bht.bhtTable_tag[2][21] ;
 wire \fetch.bht.bhtTable_tag[2][22] ;
 wire \fetch.bht.bhtTable_tag[2][23] ;
 wire \fetch.bht.bhtTable_tag[2][24] ;
 wire \fetch.bht.bhtTable_tag[2][25] ;
 wire \fetch.bht.bhtTable_tag[2][2] ;
 wire \fetch.bht.bhtTable_tag[2][3] ;
 wire \fetch.bht.bhtTable_tag[2][4] ;
 wire \fetch.bht.bhtTable_tag[2][5] ;
 wire \fetch.bht.bhtTable_tag[2][6] ;
 wire \fetch.bht.bhtTable_tag[2][7] ;
 wire \fetch.bht.bhtTable_tag[2][8] ;
 wire \fetch.bht.bhtTable_tag[2][9] ;
 wire \fetch.bht.bhtTable_tag[3][0] ;
 wire \fetch.bht.bhtTable_tag[3][10] ;
 wire \fetch.bht.bhtTable_tag[3][11] ;
 wire \fetch.bht.bhtTable_tag[3][12] ;
 wire \fetch.bht.bhtTable_tag[3][13] ;
 wire \fetch.bht.bhtTable_tag[3][14] ;
 wire \fetch.bht.bhtTable_tag[3][15] ;
 wire \fetch.bht.bhtTable_tag[3][16] ;
 wire \fetch.bht.bhtTable_tag[3][17] ;
 wire \fetch.bht.bhtTable_tag[3][18] ;
 wire \fetch.bht.bhtTable_tag[3][19] ;
 wire \fetch.bht.bhtTable_tag[3][1] ;
 wire \fetch.bht.bhtTable_tag[3][20] ;
 wire \fetch.bht.bhtTable_tag[3][21] ;
 wire \fetch.bht.bhtTable_tag[3][22] ;
 wire \fetch.bht.bhtTable_tag[3][23] ;
 wire \fetch.bht.bhtTable_tag[3][24] ;
 wire \fetch.bht.bhtTable_tag[3][25] ;
 wire \fetch.bht.bhtTable_tag[3][2] ;
 wire \fetch.bht.bhtTable_tag[3][3] ;
 wire \fetch.bht.bhtTable_tag[3][4] ;
 wire \fetch.bht.bhtTable_tag[3][5] ;
 wire \fetch.bht.bhtTable_tag[3][6] ;
 wire \fetch.bht.bhtTable_tag[3][7] ;
 wire \fetch.bht.bhtTable_tag[3][8] ;
 wire \fetch.bht.bhtTable_tag[3][9] ;
 wire \fetch.bht.bhtTable_tag[4][0] ;
 wire \fetch.bht.bhtTable_tag[4][10] ;
 wire \fetch.bht.bhtTable_tag[4][11] ;
 wire \fetch.bht.bhtTable_tag[4][12] ;
 wire \fetch.bht.bhtTable_tag[4][13] ;
 wire \fetch.bht.bhtTable_tag[4][14] ;
 wire \fetch.bht.bhtTable_tag[4][15] ;
 wire \fetch.bht.bhtTable_tag[4][16] ;
 wire \fetch.bht.bhtTable_tag[4][17] ;
 wire \fetch.bht.bhtTable_tag[4][18] ;
 wire \fetch.bht.bhtTable_tag[4][19] ;
 wire \fetch.bht.bhtTable_tag[4][1] ;
 wire \fetch.bht.bhtTable_tag[4][20] ;
 wire \fetch.bht.bhtTable_tag[4][21] ;
 wire \fetch.bht.bhtTable_tag[4][22] ;
 wire \fetch.bht.bhtTable_tag[4][23] ;
 wire \fetch.bht.bhtTable_tag[4][24] ;
 wire \fetch.bht.bhtTable_tag[4][25] ;
 wire \fetch.bht.bhtTable_tag[4][2] ;
 wire \fetch.bht.bhtTable_tag[4][3] ;
 wire \fetch.bht.bhtTable_tag[4][4] ;
 wire \fetch.bht.bhtTable_tag[4][5] ;
 wire \fetch.bht.bhtTable_tag[4][6] ;
 wire \fetch.bht.bhtTable_tag[4][7] ;
 wire \fetch.bht.bhtTable_tag[4][8] ;
 wire \fetch.bht.bhtTable_tag[4][9] ;
 wire \fetch.bht.bhtTable_tag[5][0] ;
 wire \fetch.bht.bhtTable_tag[5][10] ;
 wire \fetch.bht.bhtTable_tag[5][11] ;
 wire \fetch.bht.bhtTable_tag[5][12] ;
 wire \fetch.bht.bhtTable_tag[5][13] ;
 wire \fetch.bht.bhtTable_tag[5][14] ;
 wire \fetch.bht.bhtTable_tag[5][15] ;
 wire \fetch.bht.bhtTable_tag[5][16] ;
 wire \fetch.bht.bhtTable_tag[5][17] ;
 wire \fetch.bht.bhtTable_tag[5][18] ;
 wire \fetch.bht.bhtTable_tag[5][19] ;
 wire \fetch.bht.bhtTable_tag[5][1] ;
 wire \fetch.bht.bhtTable_tag[5][20] ;
 wire \fetch.bht.bhtTable_tag[5][21] ;
 wire \fetch.bht.bhtTable_tag[5][22] ;
 wire \fetch.bht.bhtTable_tag[5][23] ;
 wire \fetch.bht.bhtTable_tag[5][24] ;
 wire \fetch.bht.bhtTable_tag[5][25] ;
 wire \fetch.bht.bhtTable_tag[5][2] ;
 wire \fetch.bht.bhtTable_tag[5][3] ;
 wire \fetch.bht.bhtTable_tag[5][4] ;
 wire \fetch.bht.bhtTable_tag[5][5] ;
 wire \fetch.bht.bhtTable_tag[5][6] ;
 wire \fetch.bht.bhtTable_tag[5][7] ;
 wire \fetch.bht.bhtTable_tag[5][8] ;
 wire \fetch.bht.bhtTable_tag[5][9] ;
 wire \fetch.bht.bhtTable_tag[6][0] ;
 wire \fetch.bht.bhtTable_tag[6][10] ;
 wire \fetch.bht.bhtTable_tag[6][11] ;
 wire \fetch.bht.bhtTable_tag[6][12] ;
 wire \fetch.bht.bhtTable_tag[6][13] ;
 wire \fetch.bht.bhtTable_tag[6][14] ;
 wire \fetch.bht.bhtTable_tag[6][15] ;
 wire \fetch.bht.bhtTable_tag[6][16] ;
 wire \fetch.bht.bhtTable_tag[6][17] ;
 wire \fetch.bht.bhtTable_tag[6][18] ;
 wire \fetch.bht.bhtTable_tag[6][19] ;
 wire \fetch.bht.bhtTable_tag[6][1] ;
 wire \fetch.bht.bhtTable_tag[6][20] ;
 wire \fetch.bht.bhtTable_tag[6][21] ;
 wire \fetch.bht.bhtTable_tag[6][22] ;
 wire \fetch.bht.bhtTable_tag[6][23] ;
 wire \fetch.bht.bhtTable_tag[6][24] ;
 wire \fetch.bht.bhtTable_tag[6][25] ;
 wire \fetch.bht.bhtTable_tag[6][2] ;
 wire \fetch.bht.bhtTable_tag[6][3] ;
 wire \fetch.bht.bhtTable_tag[6][4] ;
 wire \fetch.bht.bhtTable_tag[6][5] ;
 wire \fetch.bht.bhtTable_tag[6][6] ;
 wire \fetch.bht.bhtTable_tag[6][7] ;
 wire \fetch.bht.bhtTable_tag[6][8] ;
 wire \fetch.bht.bhtTable_tag[6][9] ;
 wire \fetch.bht.bhtTable_tag[7][0] ;
 wire \fetch.bht.bhtTable_tag[7][10] ;
 wire \fetch.bht.bhtTable_tag[7][11] ;
 wire \fetch.bht.bhtTable_tag[7][12] ;
 wire \fetch.bht.bhtTable_tag[7][13] ;
 wire \fetch.bht.bhtTable_tag[7][14] ;
 wire \fetch.bht.bhtTable_tag[7][15] ;
 wire \fetch.bht.bhtTable_tag[7][16] ;
 wire \fetch.bht.bhtTable_tag[7][17] ;
 wire \fetch.bht.bhtTable_tag[7][18] ;
 wire \fetch.bht.bhtTable_tag[7][19] ;
 wire \fetch.bht.bhtTable_tag[7][1] ;
 wire \fetch.bht.bhtTable_tag[7][20] ;
 wire \fetch.bht.bhtTable_tag[7][21] ;
 wire \fetch.bht.bhtTable_tag[7][22] ;
 wire \fetch.bht.bhtTable_tag[7][23] ;
 wire \fetch.bht.bhtTable_tag[7][24] ;
 wire \fetch.bht.bhtTable_tag[7][25] ;
 wire \fetch.bht.bhtTable_tag[7][2] ;
 wire \fetch.bht.bhtTable_tag[7][3] ;
 wire \fetch.bht.bhtTable_tag[7][4] ;
 wire \fetch.bht.bhtTable_tag[7][5] ;
 wire \fetch.bht.bhtTable_tag[7][6] ;
 wire \fetch.bht.bhtTable_tag[7][7] ;
 wire \fetch.bht.bhtTable_tag[7][8] ;
 wire \fetch.bht.bhtTable_tag[7][9] ;
 wire \fetch.bht.bhtTable_tag[8][0] ;
 wire \fetch.bht.bhtTable_tag[8][10] ;
 wire \fetch.bht.bhtTable_tag[8][11] ;
 wire \fetch.bht.bhtTable_tag[8][12] ;
 wire \fetch.bht.bhtTable_tag[8][13] ;
 wire \fetch.bht.bhtTable_tag[8][14] ;
 wire \fetch.bht.bhtTable_tag[8][15] ;
 wire \fetch.bht.bhtTable_tag[8][16] ;
 wire \fetch.bht.bhtTable_tag[8][17] ;
 wire \fetch.bht.bhtTable_tag[8][18] ;
 wire \fetch.bht.bhtTable_tag[8][19] ;
 wire \fetch.bht.bhtTable_tag[8][1] ;
 wire \fetch.bht.bhtTable_tag[8][20] ;
 wire \fetch.bht.bhtTable_tag[8][21] ;
 wire \fetch.bht.bhtTable_tag[8][22] ;
 wire \fetch.bht.bhtTable_tag[8][23] ;
 wire \fetch.bht.bhtTable_tag[8][24] ;
 wire \fetch.bht.bhtTable_tag[8][25] ;
 wire \fetch.bht.bhtTable_tag[8][2] ;
 wire \fetch.bht.bhtTable_tag[8][3] ;
 wire \fetch.bht.bhtTable_tag[8][4] ;
 wire \fetch.bht.bhtTable_tag[8][5] ;
 wire \fetch.bht.bhtTable_tag[8][6] ;
 wire \fetch.bht.bhtTable_tag[8][7] ;
 wire \fetch.bht.bhtTable_tag[8][8] ;
 wire \fetch.bht.bhtTable_tag[8][9] ;
 wire \fetch.bht.bhtTable_tag[9][0] ;
 wire \fetch.bht.bhtTable_tag[9][10] ;
 wire \fetch.bht.bhtTable_tag[9][11] ;
 wire \fetch.bht.bhtTable_tag[9][12] ;
 wire \fetch.bht.bhtTable_tag[9][13] ;
 wire \fetch.bht.bhtTable_tag[9][14] ;
 wire \fetch.bht.bhtTable_tag[9][15] ;
 wire \fetch.bht.bhtTable_tag[9][16] ;
 wire \fetch.bht.bhtTable_tag[9][17] ;
 wire \fetch.bht.bhtTable_tag[9][18] ;
 wire \fetch.bht.bhtTable_tag[9][19] ;
 wire \fetch.bht.bhtTable_tag[9][1] ;
 wire \fetch.bht.bhtTable_tag[9][20] ;
 wire \fetch.bht.bhtTable_tag[9][21] ;
 wire \fetch.bht.bhtTable_tag[9][22] ;
 wire \fetch.bht.bhtTable_tag[9][23] ;
 wire \fetch.bht.bhtTable_tag[9][24] ;
 wire \fetch.bht.bhtTable_tag[9][25] ;
 wire \fetch.bht.bhtTable_tag[9][2] ;
 wire \fetch.bht.bhtTable_tag[9][3] ;
 wire \fetch.bht.bhtTable_tag[9][4] ;
 wire \fetch.bht.bhtTable_tag[9][5] ;
 wire \fetch.bht.bhtTable_tag[9][6] ;
 wire \fetch.bht.bhtTable_tag[9][7] ;
 wire \fetch.bht.bhtTable_tag[9][8] ;
 wire \fetch.bht.bhtTable_tag[9][9] ;
 wire \fetch.bht.bhtTable_tag_MPORT_en ;
 wire \fetch.bht.bhtTable_target_pc[0][0] ;
 wire \fetch.bht.bhtTable_target_pc[0][10] ;
 wire \fetch.bht.bhtTable_target_pc[0][11] ;
 wire \fetch.bht.bhtTable_target_pc[0][12] ;
 wire \fetch.bht.bhtTable_target_pc[0][13] ;
 wire \fetch.bht.bhtTable_target_pc[0][14] ;
 wire \fetch.bht.bhtTable_target_pc[0][15] ;
 wire \fetch.bht.bhtTable_target_pc[0][16] ;
 wire \fetch.bht.bhtTable_target_pc[0][17] ;
 wire \fetch.bht.bhtTable_target_pc[0][18] ;
 wire \fetch.bht.bhtTable_target_pc[0][19] ;
 wire \fetch.bht.bhtTable_target_pc[0][1] ;
 wire \fetch.bht.bhtTable_target_pc[0][20] ;
 wire \fetch.bht.bhtTable_target_pc[0][21] ;
 wire \fetch.bht.bhtTable_target_pc[0][22] ;
 wire \fetch.bht.bhtTable_target_pc[0][23] ;
 wire \fetch.bht.bhtTable_target_pc[0][24] ;
 wire \fetch.bht.bhtTable_target_pc[0][25] ;
 wire \fetch.bht.bhtTable_target_pc[0][26] ;
 wire \fetch.bht.bhtTable_target_pc[0][27] ;
 wire \fetch.bht.bhtTable_target_pc[0][28] ;
 wire \fetch.bht.bhtTable_target_pc[0][29] ;
 wire \fetch.bht.bhtTable_target_pc[0][2] ;
 wire \fetch.bht.bhtTable_target_pc[0][30] ;
 wire \fetch.bht.bhtTable_target_pc[0][31] ;
 wire \fetch.bht.bhtTable_target_pc[0][3] ;
 wire \fetch.bht.bhtTable_target_pc[0][4] ;
 wire \fetch.bht.bhtTable_target_pc[0][5] ;
 wire \fetch.bht.bhtTable_target_pc[0][6] ;
 wire \fetch.bht.bhtTable_target_pc[0][7] ;
 wire \fetch.bht.bhtTable_target_pc[0][8] ;
 wire \fetch.bht.bhtTable_target_pc[0][9] ;
 wire \fetch.bht.bhtTable_target_pc[10][0] ;
 wire \fetch.bht.bhtTable_target_pc[10][10] ;
 wire \fetch.bht.bhtTable_target_pc[10][11] ;
 wire \fetch.bht.bhtTable_target_pc[10][12] ;
 wire \fetch.bht.bhtTable_target_pc[10][13] ;
 wire \fetch.bht.bhtTable_target_pc[10][14] ;
 wire \fetch.bht.bhtTable_target_pc[10][15] ;
 wire \fetch.bht.bhtTable_target_pc[10][16] ;
 wire \fetch.bht.bhtTable_target_pc[10][17] ;
 wire \fetch.bht.bhtTable_target_pc[10][18] ;
 wire \fetch.bht.bhtTable_target_pc[10][19] ;
 wire \fetch.bht.bhtTable_target_pc[10][1] ;
 wire \fetch.bht.bhtTable_target_pc[10][20] ;
 wire \fetch.bht.bhtTable_target_pc[10][21] ;
 wire \fetch.bht.bhtTable_target_pc[10][22] ;
 wire \fetch.bht.bhtTable_target_pc[10][23] ;
 wire \fetch.bht.bhtTable_target_pc[10][24] ;
 wire \fetch.bht.bhtTable_target_pc[10][25] ;
 wire \fetch.bht.bhtTable_target_pc[10][26] ;
 wire \fetch.bht.bhtTable_target_pc[10][27] ;
 wire \fetch.bht.bhtTable_target_pc[10][28] ;
 wire \fetch.bht.bhtTable_target_pc[10][29] ;
 wire \fetch.bht.bhtTable_target_pc[10][2] ;
 wire \fetch.bht.bhtTable_target_pc[10][30] ;
 wire \fetch.bht.bhtTable_target_pc[10][31] ;
 wire \fetch.bht.bhtTable_target_pc[10][3] ;
 wire \fetch.bht.bhtTable_target_pc[10][4] ;
 wire \fetch.bht.bhtTable_target_pc[10][5] ;
 wire \fetch.bht.bhtTable_target_pc[10][6] ;
 wire \fetch.bht.bhtTable_target_pc[10][7] ;
 wire \fetch.bht.bhtTable_target_pc[10][8] ;
 wire \fetch.bht.bhtTable_target_pc[10][9] ;
 wire \fetch.bht.bhtTable_target_pc[11][0] ;
 wire \fetch.bht.bhtTable_target_pc[11][10] ;
 wire \fetch.bht.bhtTable_target_pc[11][11] ;
 wire \fetch.bht.bhtTable_target_pc[11][12] ;
 wire \fetch.bht.bhtTable_target_pc[11][13] ;
 wire \fetch.bht.bhtTable_target_pc[11][14] ;
 wire \fetch.bht.bhtTable_target_pc[11][15] ;
 wire \fetch.bht.bhtTable_target_pc[11][16] ;
 wire \fetch.bht.bhtTable_target_pc[11][17] ;
 wire \fetch.bht.bhtTable_target_pc[11][18] ;
 wire \fetch.bht.bhtTable_target_pc[11][19] ;
 wire \fetch.bht.bhtTable_target_pc[11][1] ;
 wire \fetch.bht.bhtTable_target_pc[11][20] ;
 wire \fetch.bht.bhtTable_target_pc[11][21] ;
 wire \fetch.bht.bhtTable_target_pc[11][22] ;
 wire \fetch.bht.bhtTable_target_pc[11][23] ;
 wire \fetch.bht.bhtTable_target_pc[11][24] ;
 wire \fetch.bht.bhtTable_target_pc[11][25] ;
 wire \fetch.bht.bhtTable_target_pc[11][26] ;
 wire \fetch.bht.bhtTable_target_pc[11][27] ;
 wire \fetch.bht.bhtTable_target_pc[11][28] ;
 wire \fetch.bht.bhtTable_target_pc[11][29] ;
 wire \fetch.bht.bhtTable_target_pc[11][2] ;
 wire \fetch.bht.bhtTable_target_pc[11][30] ;
 wire \fetch.bht.bhtTable_target_pc[11][31] ;
 wire \fetch.bht.bhtTable_target_pc[11][3] ;
 wire \fetch.bht.bhtTable_target_pc[11][4] ;
 wire \fetch.bht.bhtTable_target_pc[11][5] ;
 wire \fetch.bht.bhtTable_target_pc[11][6] ;
 wire \fetch.bht.bhtTable_target_pc[11][7] ;
 wire \fetch.bht.bhtTable_target_pc[11][8] ;
 wire \fetch.bht.bhtTable_target_pc[11][9] ;
 wire \fetch.bht.bhtTable_target_pc[12][0] ;
 wire \fetch.bht.bhtTable_target_pc[12][10] ;
 wire \fetch.bht.bhtTable_target_pc[12][11] ;
 wire \fetch.bht.bhtTable_target_pc[12][12] ;
 wire \fetch.bht.bhtTable_target_pc[12][13] ;
 wire \fetch.bht.bhtTable_target_pc[12][14] ;
 wire \fetch.bht.bhtTable_target_pc[12][15] ;
 wire \fetch.bht.bhtTable_target_pc[12][16] ;
 wire \fetch.bht.bhtTable_target_pc[12][17] ;
 wire \fetch.bht.bhtTable_target_pc[12][18] ;
 wire \fetch.bht.bhtTable_target_pc[12][19] ;
 wire \fetch.bht.bhtTable_target_pc[12][1] ;
 wire \fetch.bht.bhtTable_target_pc[12][20] ;
 wire \fetch.bht.bhtTable_target_pc[12][21] ;
 wire \fetch.bht.bhtTable_target_pc[12][22] ;
 wire \fetch.bht.bhtTable_target_pc[12][23] ;
 wire \fetch.bht.bhtTable_target_pc[12][24] ;
 wire \fetch.bht.bhtTable_target_pc[12][25] ;
 wire \fetch.bht.bhtTable_target_pc[12][26] ;
 wire \fetch.bht.bhtTable_target_pc[12][27] ;
 wire \fetch.bht.bhtTable_target_pc[12][28] ;
 wire \fetch.bht.bhtTable_target_pc[12][29] ;
 wire \fetch.bht.bhtTable_target_pc[12][2] ;
 wire \fetch.bht.bhtTable_target_pc[12][30] ;
 wire \fetch.bht.bhtTable_target_pc[12][31] ;
 wire \fetch.bht.bhtTable_target_pc[12][3] ;
 wire \fetch.bht.bhtTable_target_pc[12][4] ;
 wire \fetch.bht.bhtTable_target_pc[12][5] ;
 wire \fetch.bht.bhtTable_target_pc[12][6] ;
 wire \fetch.bht.bhtTable_target_pc[12][7] ;
 wire \fetch.bht.bhtTable_target_pc[12][8] ;
 wire \fetch.bht.bhtTable_target_pc[12][9] ;
 wire \fetch.bht.bhtTable_target_pc[13][0] ;
 wire \fetch.bht.bhtTable_target_pc[13][10] ;
 wire \fetch.bht.bhtTable_target_pc[13][11] ;
 wire \fetch.bht.bhtTable_target_pc[13][12] ;
 wire \fetch.bht.bhtTable_target_pc[13][13] ;
 wire \fetch.bht.bhtTable_target_pc[13][14] ;
 wire \fetch.bht.bhtTable_target_pc[13][15] ;
 wire \fetch.bht.bhtTable_target_pc[13][16] ;
 wire \fetch.bht.bhtTable_target_pc[13][17] ;
 wire \fetch.bht.bhtTable_target_pc[13][18] ;
 wire \fetch.bht.bhtTable_target_pc[13][19] ;
 wire \fetch.bht.bhtTable_target_pc[13][1] ;
 wire \fetch.bht.bhtTable_target_pc[13][20] ;
 wire \fetch.bht.bhtTable_target_pc[13][21] ;
 wire \fetch.bht.bhtTable_target_pc[13][22] ;
 wire \fetch.bht.bhtTable_target_pc[13][23] ;
 wire \fetch.bht.bhtTable_target_pc[13][24] ;
 wire \fetch.bht.bhtTable_target_pc[13][25] ;
 wire \fetch.bht.bhtTable_target_pc[13][26] ;
 wire \fetch.bht.bhtTable_target_pc[13][27] ;
 wire \fetch.bht.bhtTable_target_pc[13][28] ;
 wire \fetch.bht.bhtTable_target_pc[13][29] ;
 wire \fetch.bht.bhtTable_target_pc[13][2] ;
 wire \fetch.bht.bhtTable_target_pc[13][30] ;
 wire \fetch.bht.bhtTable_target_pc[13][31] ;
 wire \fetch.bht.bhtTable_target_pc[13][3] ;
 wire \fetch.bht.bhtTable_target_pc[13][4] ;
 wire \fetch.bht.bhtTable_target_pc[13][5] ;
 wire \fetch.bht.bhtTable_target_pc[13][6] ;
 wire \fetch.bht.bhtTable_target_pc[13][7] ;
 wire \fetch.bht.bhtTable_target_pc[13][8] ;
 wire \fetch.bht.bhtTable_target_pc[13][9] ;
 wire \fetch.bht.bhtTable_target_pc[14][0] ;
 wire \fetch.bht.bhtTable_target_pc[14][10] ;
 wire \fetch.bht.bhtTable_target_pc[14][11] ;
 wire \fetch.bht.bhtTable_target_pc[14][12] ;
 wire \fetch.bht.bhtTable_target_pc[14][13] ;
 wire \fetch.bht.bhtTable_target_pc[14][14] ;
 wire \fetch.bht.bhtTable_target_pc[14][15] ;
 wire \fetch.bht.bhtTable_target_pc[14][16] ;
 wire \fetch.bht.bhtTable_target_pc[14][17] ;
 wire \fetch.bht.bhtTable_target_pc[14][18] ;
 wire \fetch.bht.bhtTable_target_pc[14][19] ;
 wire \fetch.bht.bhtTable_target_pc[14][1] ;
 wire \fetch.bht.bhtTable_target_pc[14][20] ;
 wire \fetch.bht.bhtTable_target_pc[14][21] ;
 wire \fetch.bht.bhtTable_target_pc[14][22] ;
 wire \fetch.bht.bhtTable_target_pc[14][23] ;
 wire \fetch.bht.bhtTable_target_pc[14][24] ;
 wire \fetch.bht.bhtTable_target_pc[14][25] ;
 wire \fetch.bht.bhtTable_target_pc[14][26] ;
 wire \fetch.bht.bhtTable_target_pc[14][27] ;
 wire \fetch.bht.bhtTable_target_pc[14][28] ;
 wire \fetch.bht.bhtTable_target_pc[14][29] ;
 wire \fetch.bht.bhtTable_target_pc[14][2] ;
 wire \fetch.bht.bhtTable_target_pc[14][30] ;
 wire \fetch.bht.bhtTable_target_pc[14][31] ;
 wire \fetch.bht.bhtTable_target_pc[14][3] ;
 wire \fetch.bht.bhtTable_target_pc[14][4] ;
 wire \fetch.bht.bhtTable_target_pc[14][5] ;
 wire \fetch.bht.bhtTable_target_pc[14][6] ;
 wire \fetch.bht.bhtTable_target_pc[14][7] ;
 wire \fetch.bht.bhtTable_target_pc[14][8] ;
 wire \fetch.bht.bhtTable_target_pc[14][9] ;
 wire \fetch.bht.bhtTable_target_pc[15][0] ;
 wire \fetch.bht.bhtTable_target_pc[15][10] ;
 wire \fetch.bht.bhtTable_target_pc[15][11] ;
 wire \fetch.bht.bhtTable_target_pc[15][12] ;
 wire \fetch.bht.bhtTable_target_pc[15][13] ;
 wire \fetch.bht.bhtTable_target_pc[15][14] ;
 wire \fetch.bht.bhtTable_target_pc[15][15] ;
 wire \fetch.bht.bhtTable_target_pc[15][16] ;
 wire \fetch.bht.bhtTable_target_pc[15][17] ;
 wire \fetch.bht.bhtTable_target_pc[15][18] ;
 wire \fetch.bht.bhtTable_target_pc[15][19] ;
 wire \fetch.bht.bhtTable_target_pc[15][1] ;
 wire \fetch.bht.bhtTable_target_pc[15][20] ;
 wire \fetch.bht.bhtTable_target_pc[15][21] ;
 wire \fetch.bht.bhtTable_target_pc[15][22] ;
 wire \fetch.bht.bhtTable_target_pc[15][23] ;
 wire \fetch.bht.bhtTable_target_pc[15][24] ;
 wire \fetch.bht.bhtTable_target_pc[15][25] ;
 wire \fetch.bht.bhtTable_target_pc[15][26] ;
 wire \fetch.bht.bhtTable_target_pc[15][27] ;
 wire \fetch.bht.bhtTable_target_pc[15][28] ;
 wire \fetch.bht.bhtTable_target_pc[15][29] ;
 wire \fetch.bht.bhtTable_target_pc[15][2] ;
 wire \fetch.bht.bhtTable_target_pc[15][30] ;
 wire \fetch.bht.bhtTable_target_pc[15][31] ;
 wire \fetch.bht.bhtTable_target_pc[15][3] ;
 wire \fetch.bht.bhtTable_target_pc[15][4] ;
 wire \fetch.bht.bhtTable_target_pc[15][5] ;
 wire \fetch.bht.bhtTable_target_pc[15][6] ;
 wire \fetch.bht.bhtTable_target_pc[15][7] ;
 wire \fetch.bht.bhtTable_target_pc[15][8] ;
 wire \fetch.bht.bhtTable_target_pc[15][9] ;
 wire \fetch.bht.bhtTable_target_pc[1][0] ;
 wire \fetch.bht.bhtTable_target_pc[1][10] ;
 wire \fetch.bht.bhtTable_target_pc[1][11] ;
 wire \fetch.bht.bhtTable_target_pc[1][12] ;
 wire \fetch.bht.bhtTable_target_pc[1][13] ;
 wire \fetch.bht.bhtTable_target_pc[1][14] ;
 wire \fetch.bht.bhtTable_target_pc[1][15] ;
 wire \fetch.bht.bhtTable_target_pc[1][16] ;
 wire \fetch.bht.bhtTable_target_pc[1][17] ;
 wire \fetch.bht.bhtTable_target_pc[1][18] ;
 wire \fetch.bht.bhtTable_target_pc[1][19] ;
 wire \fetch.bht.bhtTable_target_pc[1][1] ;
 wire \fetch.bht.bhtTable_target_pc[1][20] ;
 wire \fetch.bht.bhtTable_target_pc[1][21] ;
 wire \fetch.bht.bhtTable_target_pc[1][22] ;
 wire \fetch.bht.bhtTable_target_pc[1][23] ;
 wire \fetch.bht.bhtTable_target_pc[1][24] ;
 wire \fetch.bht.bhtTable_target_pc[1][25] ;
 wire \fetch.bht.bhtTable_target_pc[1][26] ;
 wire \fetch.bht.bhtTable_target_pc[1][27] ;
 wire \fetch.bht.bhtTable_target_pc[1][28] ;
 wire \fetch.bht.bhtTable_target_pc[1][29] ;
 wire \fetch.bht.bhtTable_target_pc[1][2] ;
 wire \fetch.bht.bhtTable_target_pc[1][30] ;
 wire \fetch.bht.bhtTable_target_pc[1][31] ;
 wire \fetch.bht.bhtTable_target_pc[1][3] ;
 wire \fetch.bht.bhtTable_target_pc[1][4] ;
 wire \fetch.bht.bhtTable_target_pc[1][5] ;
 wire \fetch.bht.bhtTable_target_pc[1][6] ;
 wire \fetch.bht.bhtTable_target_pc[1][7] ;
 wire \fetch.bht.bhtTable_target_pc[1][8] ;
 wire \fetch.bht.bhtTable_target_pc[1][9] ;
 wire \fetch.bht.bhtTable_target_pc[2][0] ;
 wire \fetch.bht.bhtTable_target_pc[2][10] ;
 wire \fetch.bht.bhtTable_target_pc[2][11] ;
 wire \fetch.bht.bhtTable_target_pc[2][12] ;
 wire \fetch.bht.bhtTable_target_pc[2][13] ;
 wire \fetch.bht.bhtTable_target_pc[2][14] ;
 wire \fetch.bht.bhtTable_target_pc[2][15] ;
 wire \fetch.bht.bhtTable_target_pc[2][16] ;
 wire \fetch.bht.bhtTable_target_pc[2][17] ;
 wire \fetch.bht.bhtTable_target_pc[2][18] ;
 wire \fetch.bht.bhtTable_target_pc[2][19] ;
 wire \fetch.bht.bhtTable_target_pc[2][1] ;
 wire \fetch.bht.bhtTable_target_pc[2][20] ;
 wire \fetch.bht.bhtTable_target_pc[2][21] ;
 wire \fetch.bht.bhtTable_target_pc[2][22] ;
 wire \fetch.bht.bhtTable_target_pc[2][23] ;
 wire \fetch.bht.bhtTable_target_pc[2][24] ;
 wire \fetch.bht.bhtTable_target_pc[2][25] ;
 wire \fetch.bht.bhtTable_target_pc[2][26] ;
 wire \fetch.bht.bhtTable_target_pc[2][27] ;
 wire \fetch.bht.bhtTable_target_pc[2][28] ;
 wire \fetch.bht.bhtTable_target_pc[2][29] ;
 wire \fetch.bht.bhtTable_target_pc[2][2] ;
 wire \fetch.bht.bhtTable_target_pc[2][30] ;
 wire \fetch.bht.bhtTable_target_pc[2][31] ;
 wire \fetch.bht.bhtTable_target_pc[2][3] ;
 wire \fetch.bht.bhtTable_target_pc[2][4] ;
 wire \fetch.bht.bhtTable_target_pc[2][5] ;
 wire \fetch.bht.bhtTable_target_pc[2][6] ;
 wire \fetch.bht.bhtTable_target_pc[2][7] ;
 wire \fetch.bht.bhtTable_target_pc[2][8] ;
 wire \fetch.bht.bhtTable_target_pc[2][9] ;
 wire \fetch.bht.bhtTable_target_pc[3][0] ;
 wire \fetch.bht.bhtTable_target_pc[3][10] ;
 wire \fetch.bht.bhtTable_target_pc[3][11] ;
 wire \fetch.bht.bhtTable_target_pc[3][12] ;
 wire \fetch.bht.bhtTable_target_pc[3][13] ;
 wire \fetch.bht.bhtTable_target_pc[3][14] ;
 wire \fetch.bht.bhtTable_target_pc[3][15] ;
 wire \fetch.bht.bhtTable_target_pc[3][16] ;
 wire \fetch.bht.bhtTable_target_pc[3][17] ;
 wire \fetch.bht.bhtTable_target_pc[3][18] ;
 wire \fetch.bht.bhtTable_target_pc[3][19] ;
 wire \fetch.bht.bhtTable_target_pc[3][1] ;
 wire \fetch.bht.bhtTable_target_pc[3][20] ;
 wire \fetch.bht.bhtTable_target_pc[3][21] ;
 wire \fetch.bht.bhtTable_target_pc[3][22] ;
 wire \fetch.bht.bhtTable_target_pc[3][23] ;
 wire \fetch.bht.bhtTable_target_pc[3][24] ;
 wire \fetch.bht.bhtTable_target_pc[3][25] ;
 wire \fetch.bht.bhtTable_target_pc[3][26] ;
 wire \fetch.bht.bhtTable_target_pc[3][27] ;
 wire \fetch.bht.bhtTable_target_pc[3][28] ;
 wire \fetch.bht.bhtTable_target_pc[3][29] ;
 wire \fetch.bht.bhtTable_target_pc[3][2] ;
 wire \fetch.bht.bhtTable_target_pc[3][30] ;
 wire \fetch.bht.bhtTable_target_pc[3][31] ;
 wire \fetch.bht.bhtTable_target_pc[3][3] ;
 wire \fetch.bht.bhtTable_target_pc[3][4] ;
 wire \fetch.bht.bhtTable_target_pc[3][5] ;
 wire \fetch.bht.bhtTable_target_pc[3][6] ;
 wire \fetch.bht.bhtTable_target_pc[3][7] ;
 wire \fetch.bht.bhtTable_target_pc[3][8] ;
 wire \fetch.bht.bhtTable_target_pc[3][9] ;
 wire \fetch.bht.bhtTable_target_pc[4][0] ;
 wire \fetch.bht.bhtTable_target_pc[4][10] ;
 wire \fetch.bht.bhtTable_target_pc[4][11] ;
 wire \fetch.bht.bhtTable_target_pc[4][12] ;
 wire \fetch.bht.bhtTable_target_pc[4][13] ;
 wire \fetch.bht.bhtTable_target_pc[4][14] ;
 wire \fetch.bht.bhtTable_target_pc[4][15] ;
 wire \fetch.bht.bhtTable_target_pc[4][16] ;
 wire \fetch.bht.bhtTable_target_pc[4][17] ;
 wire \fetch.bht.bhtTable_target_pc[4][18] ;
 wire \fetch.bht.bhtTable_target_pc[4][19] ;
 wire \fetch.bht.bhtTable_target_pc[4][1] ;
 wire \fetch.bht.bhtTable_target_pc[4][20] ;
 wire \fetch.bht.bhtTable_target_pc[4][21] ;
 wire \fetch.bht.bhtTable_target_pc[4][22] ;
 wire \fetch.bht.bhtTable_target_pc[4][23] ;
 wire \fetch.bht.bhtTable_target_pc[4][24] ;
 wire \fetch.bht.bhtTable_target_pc[4][25] ;
 wire \fetch.bht.bhtTable_target_pc[4][26] ;
 wire \fetch.bht.bhtTable_target_pc[4][27] ;
 wire \fetch.bht.bhtTable_target_pc[4][28] ;
 wire \fetch.bht.bhtTable_target_pc[4][29] ;
 wire \fetch.bht.bhtTable_target_pc[4][2] ;
 wire \fetch.bht.bhtTable_target_pc[4][30] ;
 wire \fetch.bht.bhtTable_target_pc[4][31] ;
 wire \fetch.bht.bhtTable_target_pc[4][3] ;
 wire \fetch.bht.bhtTable_target_pc[4][4] ;
 wire \fetch.bht.bhtTable_target_pc[4][5] ;
 wire \fetch.bht.bhtTable_target_pc[4][6] ;
 wire \fetch.bht.bhtTable_target_pc[4][7] ;
 wire \fetch.bht.bhtTable_target_pc[4][8] ;
 wire \fetch.bht.bhtTable_target_pc[4][9] ;
 wire \fetch.bht.bhtTable_target_pc[5][0] ;
 wire \fetch.bht.bhtTable_target_pc[5][10] ;
 wire \fetch.bht.bhtTable_target_pc[5][11] ;
 wire \fetch.bht.bhtTable_target_pc[5][12] ;
 wire \fetch.bht.bhtTable_target_pc[5][13] ;
 wire \fetch.bht.bhtTable_target_pc[5][14] ;
 wire \fetch.bht.bhtTable_target_pc[5][15] ;
 wire \fetch.bht.bhtTable_target_pc[5][16] ;
 wire \fetch.bht.bhtTable_target_pc[5][17] ;
 wire \fetch.bht.bhtTable_target_pc[5][18] ;
 wire \fetch.bht.bhtTable_target_pc[5][19] ;
 wire \fetch.bht.bhtTable_target_pc[5][1] ;
 wire \fetch.bht.bhtTable_target_pc[5][20] ;
 wire \fetch.bht.bhtTable_target_pc[5][21] ;
 wire \fetch.bht.bhtTable_target_pc[5][22] ;
 wire \fetch.bht.bhtTable_target_pc[5][23] ;
 wire \fetch.bht.bhtTable_target_pc[5][24] ;
 wire \fetch.bht.bhtTable_target_pc[5][25] ;
 wire \fetch.bht.bhtTable_target_pc[5][26] ;
 wire \fetch.bht.bhtTable_target_pc[5][27] ;
 wire \fetch.bht.bhtTable_target_pc[5][28] ;
 wire \fetch.bht.bhtTable_target_pc[5][29] ;
 wire \fetch.bht.bhtTable_target_pc[5][2] ;
 wire \fetch.bht.bhtTable_target_pc[5][30] ;
 wire \fetch.bht.bhtTable_target_pc[5][31] ;
 wire \fetch.bht.bhtTable_target_pc[5][3] ;
 wire \fetch.bht.bhtTable_target_pc[5][4] ;
 wire \fetch.bht.bhtTable_target_pc[5][5] ;
 wire \fetch.bht.bhtTable_target_pc[5][6] ;
 wire \fetch.bht.bhtTable_target_pc[5][7] ;
 wire \fetch.bht.bhtTable_target_pc[5][8] ;
 wire \fetch.bht.bhtTable_target_pc[5][9] ;
 wire \fetch.bht.bhtTable_target_pc[6][0] ;
 wire \fetch.bht.bhtTable_target_pc[6][10] ;
 wire \fetch.bht.bhtTable_target_pc[6][11] ;
 wire \fetch.bht.bhtTable_target_pc[6][12] ;
 wire \fetch.bht.bhtTable_target_pc[6][13] ;
 wire \fetch.bht.bhtTable_target_pc[6][14] ;
 wire \fetch.bht.bhtTable_target_pc[6][15] ;
 wire \fetch.bht.bhtTable_target_pc[6][16] ;
 wire \fetch.bht.bhtTable_target_pc[6][17] ;
 wire \fetch.bht.bhtTable_target_pc[6][18] ;
 wire \fetch.bht.bhtTable_target_pc[6][19] ;
 wire \fetch.bht.bhtTable_target_pc[6][1] ;
 wire \fetch.bht.bhtTable_target_pc[6][20] ;
 wire \fetch.bht.bhtTable_target_pc[6][21] ;
 wire \fetch.bht.bhtTable_target_pc[6][22] ;
 wire \fetch.bht.bhtTable_target_pc[6][23] ;
 wire \fetch.bht.bhtTable_target_pc[6][24] ;
 wire \fetch.bht.bhtTable_target_pc[6][25] ;
 wire \fetch.bht.bhtTable_target_pc[6][26] ;
 wire \fetch.bht.bhtTable_target_pc[6][27] ;
 wire \fetch.bht.bhtTable_target_pc[6][28] ;
 wire \fetch.bht.bhtTable_target_pc[6][29] ;
 wire \fetch.bht.bhtTable_target_pc[6][2] ;
 wire \fetch.bht.bhtTable_target_pc[6][30] ;
 wire \fetch.bht.bhtTable_target_pc[6][31] ;
 wire \fetch.bht.bhtTable_target_pc[6][3] ;
 wire \fetch.bht.bhtTable_target_pc[6][4] ;
 wire \fetch.bht.bhtTable_target_pc[6][5] ;
 wire \fetch.bht.bhtTable_target_pc[6][6] ;
 wire \fetch.bht.bhtTable_target_pc[6][7] ;
 wire \fetch.bht.bhtTable_target_pc[6][8] ;
 wire \fetch.bht.bhtTable_target_pc[6][9] ;
 wire \fetch.bht.bhtTable_target_pc[7][0] ;
 wire \fetch.bht.bhtTable_target_pc[7][10] ;
 wire \fetch.bht.bhtTable_target_pc[7][11] ;
 wire \fetch.bht.bhtTable_target_pc[7][12] ;
 wire \fetch.bht.bhtTable_target_pc[7][13] ;
 wire \fetch.bht.bhtTable_target_pc[7][14] ;
 wire \fetch.bht.bhtTable_target_pc[7][15] ;
 wire \fetch.bht.bhtTable_target_pc[7][16] ;
 wire \fetch.bht.bhtTable_target_pc[7][17] ;
 wire \fetch.bht.bhtTable_target_pc[7][18] ;
 wire \fetch.bht.bhtTable_target_pc[7][19] ;
 wire \fetch.bht.bhtTable_target_pc[7][1] ;
 wire \fetch.bht.bhtTable_target_pc[7][20] ;
 wire \fetch.bht.bhtTable_target_pc[7][21] ;
 wire \fetch.bht.bhtTable_target_pc[7][22] ;
 wire \fetch.bht.bhtTable_target_pc[7][23] ;
 wire \fetch.bht.bhtTable_target_pc[7][24] ;
 wire \fetch.bht.bhtTable_target_pc[7][25] ;
 wire \fetch.bht.bhtTable_target_pc[7][26] ;
 wire \fetch.bht.bhtTable_target_pc[7][27] ;
 wire \fetch.bht.bhtTable_target_pc[7][28] ;
 wire \fetch.bht.bhtTable_target_pc[7][29] ;
 wire \fetch.bht.bhtTable_target_pc[7][2] ;
 wire \fetch.bht.bhtTable_target_pc[7][30] ;
 wire \fetch.bht.bhtTable_target_pc[7][31] ;
 wire \fetch.bht.bhtTable_target_pc[7][3] ;
 wire \fetch.bht.bhtTable_target_pc[7][4] ;
 wire \fetch.bht.bhtTable_target_pc[7][5] ;
 wire \fetch.bht.bhtTable_target_pc[7][6] ;
 wire \fetch.bht.bhtTable_target_pc[7][7] ;
 wire \fetch.bht.bhtTable_target_pc[7][8] ;
 wire \fetch.bht.bhtTable_target_pc[7][9] ;
 wire \fetch.bht.bhtTable_target_pc[8][0] ;
 wire \fetch.bht.bhtTable_target_pc[8][10] ;
 wire \fetch.bht.bhtTable_target_pc[8][11] ;
 wire \fetch.bht.bhtTable_target_pc[8][12] ;
 wire \fetch.bht.bhtTable_target_pc[8][13] ;
 wire \fetch.bht.bhtTable_target_pc[8][14] ;
 wire \fetch.bht.bhtTable_target_pc[8][15] ;
 wire \fetch.bht.bhtTable_target_pc[8][16] ;
 wire \fetch.bht.bhtTable_target_pc[8][17] ;
 wire \fetch.bht.bhtTable_target_pc[8][18] ;
 wire \fetch.bht.bhtTable_target_pc[8][19] ;
 wire \fetch.bht.bhtTable_target_pc[8][1] ;
 wire \fetch.bht.bhtTable_target_pc[8][20] ;
 wire \fetch.bht.bhtTable_target_pc[8][21] ;
 wire \fetch.bht.bhtTable_target_pc[8][22] ;
 wire \fetch.bht.bhtTable_target_pc[8][23] ;
 wire \fetch.bht.bhtTable_target_pc[8][24] ;
 wire \fetch.bht.bhtTable_target_pc[8][25] ;
 wire \fetch.bht.bhtTable_target_pc[8][26] ;
 wire \fetch.bht.bhtTable_target_pc[8][27] ;
 wire \fetch.bht.bhtTable_target_pc[8][28] ;
 wire \fetch.bht.bhtTable_target_pc[8][29] ;
 wire \fetch.bht.bhtTable_target_pc[8][2] ;
 wire \fetch.bht.bhtTable_target_pc[8][30] ;
 wire \fetch.bht.bhtTable_target_pc[8][31] ;
 wire \fetch.bht.bhtTable_target_pc[8][3] ;
 wire \fetch.bht.bhtTable_target_pc[8][4] ;
 wire \fetch.bht.bhtTable_target_pc[8][5] ;
 wire \fetch.bht.bhtTable_target_pc[8][6] ;
 wire \fetch.bht.bhtTable_target_pc[8][7] ;
 wire \fetch.bht.bhtTable_target_pc[8][8] ;
 wire \fetch.bht.bhtTable_target_pc[8][9] ;
 wire \fetch.bht.bhtTable_target_pc[9][0] ;
 wire \fetch.bht.bhtTable_target_pc[9][10] ;
 wire \fetch.bht.bhtTable_target_pc[9][11] ;
 wire \fetch.bht.bhtTable_target_pc[9][12] ;
 wire \fetch.bht.bhtTable_target_pc[9][13] ;
 wire \fetch.bht.bhtTable_target_pc[9][14] ;
 wire \fetch.bht.bhtTable_target_pc[9][15] ;
 wire \fetch.bht.bhtTable_target_pc[9][16] ;
 wire \fetch.bht.bhtTable_target_pc[9][17] ;
 wire \fetch.bht.bhtTable_target_pc[9][18] ;
 wire \fetch.bht.bhtTable_target_pc[9][19] ;
 wire \fetch.bht.bhtTable_target_pc[9][1] ;
 wire \fetch.bht.bhtTable_target_pc[9][20] ;
 wire \fetch.bht.bhtTable_target_pc[9][21] ;
 wire \fetch.bht.bhtTable_target_pc[9][22] ;
 wire \fetch.bht.bhtTable_target_pc[9][23] ;
 wire \fetch.bht.bhtTable_target_pc[9][24] ;
 wire \fetch.bht.bhtTable_target_pc[9][25] ;
 wire \fetch.bht.bhtTable_target_pc[9][26] ;
 wire \fetch.bht.bhtTable_target_pc[9][27] ;
 wire \fetch.bht.bhtTable_target_pc[9][28] ;
 wire \fetch.bht.bhtTable_target_pc[9][29] ;
 wire \fetch.bht.bhtTable_target_pc[9][2] ;
 wire \fetch.bht.bhtTable_target_pc[9][30] ;
 wire \fetch.bht.bhtTable_target_pc[9][31] ;
 wire \fetch.bht.bhtTable_target_pc[9][3] ;
 wire \fetch.bht.bhtTable_target_pc[9][4] ;
 wire \fetch.bht.bhtTable_target_pc[9][5] ;
 wire \fetch.bht.bhtTable_target_pc[9][6] ;
 wire \fetch.bht.bhtTable_target_pc[9][7] ;
 wire \fetch.bht.bhtTable_target_pc[9][8] ;
 wire \fetch.bht.bhtTable_target_pc[9][9] ;
 wire \fetch.bht.bhtTable_valid[0] ;
 wire \fetch.bht.bhtTable_valid[10] ;
 wire \fetch.bht.bhtTable_valid[11] ;
 wire \fetch.bht.bhtTable_valid[12] ;
 wire \fetch.bht.bhtTable_valid[13] ;
 wire \fetch.bht.bhtTable_valid[14] ;
 wire \fetch.bht.bhtTable_valid[15] ;
 wire \fetch.bht.bhtTable_valid[1] ;
 wire \fetch.bht.bhtTable_valid[2] ;
 wire \fetch.bht.bhtTable_valid[3] ;
 wire \fetch.bht.bhtTable_valid[4] ;
 wire \fetch.bht.bhtTable_valid[5] ;
 wire \fetch.bht.bhtTable_valid[6] ;
 wire \fetch.bht.bhtTable_valid[7] ;
 wire \fetch.bht.bhtTable_valid[8] ;
 wire \fetch.bht.bhtTable_valid[9] ;
 wire \fetch.btb.btbTable[0][0] ;
 wire \fetch.btb.btbTable[0][1] ;
 wire \fetch.btb.btbTable[10][0] ;
 wire \fetch.btb.btbTable[10][1] ;
 wire \fetch.btb.btbTable[11][0] ;
 wire \fetch.btb.btbTable[11][1] ;
 wire \fetch.btb.btbTable[12][0] ;
 wire \fetch.btb.btbTable[12][1] ;
 wire \fetch.btb.btbTable[13][0] ;
 wire \fetch.btb.btbTable[13][1] ;
 wire \fetch.btb.btbTable[14][0] ;
 wire \fetch.btb.btbTable[14][1] ;
 wire \fetch.btb.btbTable[15][0] ;
 wire \fetch.btb.btbTable[15][1] ;
 wire \fetch.btb.btbTable[1][0] ;
 wire \fetch.btb.btbTable[1][1] ;
 wire \fetch.btb.btbTable[2][0] ;
 wire \fetch.btb.btbTable[2][1] ;
 wire \fetch.btb.btbTable[3][0] ;
 wire \fetch.btb.btbTable[3][1] ;
 wire \fetch.btb.btbTable[4][0] ;
 wire \fetch.btb.btbTable[4][1] ;
 wire \fetch.btb.btbTable[5][0] ;
 wire \fetch.btb.btbTable[5][1] ;
 wire \fetch.btb.btbTable[6][0] ;
 wire \fetch.btb.btbTable[6][1] ;
 wire \fetch.btb.btbTable[7][0] ;
 wire \fetch.btb.btbTable[7][1] ;
 wire \fetch.btb.btbTable[8][0] ;
 wire \fetch.btb.btbTable[8][1] ;
 wire \fetch.btb.btbTable[9][0] ;
 wire \fetch.btb.btbTable[9][1] ;
 wire \fetch.btb.io_branch ;
 wire \memory.csr_read_data_out_reg[0] ;
 wire \memory.csr_read_data_out_reg[10] ;
 wire \memory.csr_read_data_out_reg[11] ;
 wire \memory.csr_read_data_out_reg[12] ;
 wire \memory.csr_read_data_out_reg[13] ;
 wire \memory.csr_read_data_out_reg[14] ;
 wire \memory.csr_read_data_out_reg[15] ;
 wire \memory.csr_read_data_out_reg[16] ;
 wire \memory.csr_read_data_out_reg[17] ;
 wire \memory.csr_read_data_out_reg[18] ;
 wire \memory.csr_read_data_out_reg[19] ;
 wire \memory.csr_read_data_out_reg[1] ;
 wire \memory.csr_read_data_out_reg[20] ;
 wire \memory.csr_read_data_out_reg[21] ;
 wire \memory.csr_read_data_out_reg[22] ;
 wire \memory.csr_read_data_out_reg[23] ;
 wire \memory.csr_read_data_out_reg[24] ;
 wire \memory.csr_read_data_out_reg[25] ;
 wire \memory.csr_read_data_out_reg[26] ;
 wire \memory.csr_read_data_out_reg[27] ;
 wire \memory.csr_read_data_out_reg[28] ;
 wire \memory.csr_read_data_out_reg[29] ;
 wire \memory.csr_read_data_out_reg[2] ;
 wire \memory.csr_read_data_out_reg[30] ;
 wire \memory.csr_read_data_out_reg[31] ;
 wire \memory.csr_read_data_out_reg[3] ;
 wire \memory.csr_read_data_out_reg[4] ;
 wire \memory.csr_read_data_out_reg[5] ;
 wire \memory.csr_read_data_out_reg[6] ;
 wire \memory.csr_read_data_out_reg[7] ;
 wire \memory.csr_read_data_out_reg[8] ;
 wire \memory.csr_read_data_out_reg[9] ;
 wire \memory.io_wb_aluresult[0] ;
 wire \memory.io_wb_aluresult[10] ;
 wire \memory.io_wb_aluresult[11] ;
 wire \memory.io_wb_aluresult[12] ;
 wire \memory.io_wb_aluresult[13] ;
 wire \memory.io_wb_aluresult[14] ;
 wire \memory.io_wb_aluresult[15] ;
 wire \memory.io_wb_aluresult[16] ;
 wire \memory.io_wb_aluresult[17] ;
 wire \memory.io_wb_aluresult[18] ;
 wire \memory.io_wb_aluresult[19] ;
 wire \memory.io_wb_aluresult[1] ;
 wire \memory.io_wb_aluresult[20] ;
 wire \memory.io_wb_aluresult[21] ;
 wire \memory.io_wb_aluresult[22] ;
 wire \memory.io_wb_aluresult[23] ;
 wire \memory.io_wb_aluresult[24] ;
 wire \memory.io_wb_aluresult[25] ;
 wire \memory.io_wb_aluresult[26] ;
 wire \memory.io_wb_aluresult[27] ;
 wire \memory.io_wb_aluresult[28] ;
 wire \memory.io_wb_aluresult[29] ;
 wire \memory.io_wb_aluresult[2] ;
 wire \memory.io_wb_aluresult[30] ;
 wire \memory.io_wb_aluresult[31] ;
 wire \memory.io_wb_aluresult[3] ;
 wire \memory.io_wb_aluresult[4] ;
 wire \memory.io_wb_aluresult[5] ;
 wire \memory.io_wb_aluresult[6] ;
 wire \memory.io_wb_aluresult[7] ;
 wire \memory.io_wb_aluresult[8] ;
 wire \memory.io_wb_aluresult[9] ;
 wire \memory.io_wb_memtoreg[0] ;
 wire \memory.io_wb_memtoreg[1] ;
 wire \memory.io_wb_readdata[0] ;
 wire \memory.io_wb_readdata[10] ;
 wire \memory.io_wb_readdata[11] ;
 wire \memory.io_wb_readdata[12] ;
 wire \memory.io_wb_readdata[13] ;
 wire \memory.io_wb_readdata[14] ;
 wire \memory.io_wb_readdata[15] ;
 wire \memory.io_wb_readdata[16] ;
 wire \memory.io_wb_readdata[17] ;
 wire \memory.io_wb_readdata[18] ;
 wire \memory.io_wb_readdata[19] ;
 wire \memory.io_wb_readdata[1] ;
 wire \memory.io_wb_readdata[20] ;
 wire \memory.io_wb_readdata[21] ;
 wire \memory.io_wb_readdata[22] ;
 wire \memory.io_wb_readdata[23] ;
 wire \memory.io_wb_readdata[24] ;
 wire \memory.io_wb_readdata[25] ;
 wire \memory.io_wb_readdata[26] ;
 wire \memory.io_wb_readdata[27] ;
 wire \memory.io_wb_readdata[28] ;
 wire \memory.io_wb_readdata[29] ;
 wire \memory.io_wb_readdata[2] ;
 wire \memory.io_wb_readdata[30] ;
 wire \memory.io_wb_readdata[31] ;
 wire \memory.io_wb_readdata[3] ;
 wire \memory.io_wb_readdata[4] ;
 wire \memory.io_wb_readdata[5] ;
 wire \memory.io_wb_readdata[6] ;
 wire \memory.io_wb_readdata[7] ;
 wire \memory.io_wb_readdata[8] ;
 wire \memory.io_wb_readdata[9] ;
 wire \memory.io_wb_reg_pc[0] ;
 wire \memory.io_wb_reg_pc[10] ;
 wire \memory.io_wb_reg_pc[11] ;
 wire \memory.io_wb_reg_pc[12] ;
 wire \memory.io_wb_reg_pc[13] ;
 wire \memory.io_wb_reg_pc[14] ;
 wire \memory.io_wb_reg_pc[15] ;
 wire \memory.io_wb_reg_pc[16] ;
 wire \memory.io_wb_reg_pc[17] ;
 wire \memory.io_wb_reg_pc[18] ;
 wire \memory.io_wb_reg_pc[19] ;
 wire \memory.io_wb_reg_pc[1] ;
 wire \memory.io_wb_reg_pc[20] ;
 wire \memory.io_wb_reg_pc[21] ;
 wire \memory.io_wb_reg_pc[22] ;
 wire \memory.io_wb_reg_pc[23] ;
 wire \memory.io_wb_reg_pc[24] ;
 wire \memory.io_wb_reg_pc[25] ;
 wire \memory.io_wb_reg_pc[26] ;
 wire \memory.io_wb_reg_pc[27] ;
 wire \memory.io_wb_reg_pc[28] ;
 wire \memory.io_wb_reg_pc[29] ;
 wire \memory.io_wb_reg_pc[2] ;
 wire \memory.io_wb_reg_pc[30] ;
 wire \memory.io_wb_reg_pc[31] ;
 wire \memory.io_wb_reg_pc[3] ;
 wire \memory.io_wb_reg_pc[4] ;
 wire \memory.io_wb_reg_pc[5] ;
 wire \memory.io_wb_reg_pc[6] ;
 wire \memory.io_wb_reg_pc[7] ;
 wire \memory.io_wb_reg_pc[8] ;
 wire \memory.io_wb_reg_pc[9] ;

 sky130_fd_sc_hd__buf_1 _13497_ (.A(\csr.io_mem_pc[4] ),
    .X(_09879_));
 sky130_fd_sc_hd__buf_1 _13498_ (.A(_09879_),
    .X(_09880_));
 sky130_fd_sc_hd__buf_1 _13499_ (.A(_09880_),
    .X(_09881_));
 sky130_fd_sc_hd__buf_1 _13500_ (.A(\csr.io_mem_pc[5] ),
    .X(_09882_));
 sky130_fd_sc_hd__buf_1 _13501_ (.A(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__buf_1 _13502_ (.A(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__buf_1 _13503_ (.A(\fetch.bht.bhtTable_tag_MPORT_en ),
    .X(_09885_));
 sky130_fd_sc_hd__and2b_2 _13504_ (.A_N(\csr.io_mem_pc[2] ),
    .B(\csr.io_mem_pc[3] ),
    .X(_09886_));
 sky130_fd_sc_hd__buf_1 _13505_ (.A(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__a41o_2 _13506_ (.A1(_09881_),
    .A2(_09884_),
    .A3(_09885_),
    .A4(_09887_),
    .B1(\fetch.bht.bhtTable_valid[14] ),
    .X(_00009_));
 sky130_fd_sc_hd__buf_1 _13507_ (.A(\csr.io_mem_pc[3] ),
    .X(_09888_));
 sky130_fd_sc_hd__and2b_2 _13508_ (.A_N(_09888_),
    .B(\csr.io_mem_pc[2] ),
    .X(_09889_));
 sky130_fd_sc_hd__buf_1 _13509_ (.A(_09889_),
    .X(_09890_));
 sky130_fd_sc_hd__a41o_2 _13510_ (.A1(_09881_),
    .A2(_09884_),
    .A3(_09885_),
    .A4(_09890_),
    .B1(\fetch.bht.bhtTable_valid[13] ),
    .X(_00008_));
 sky130_fd_sc_hd__buf_1 _13511_ (.A(\csr.io_mem_pc[2] ),
    .X(_09891_));
 sky130_fd_sc_hd__nor2_2 _13512_ (.A(_09891_),
    .B(_09888_),
    .Y(_09892_));
 sky130_fd_sc_hd__a41o_2 _13513_ (.A1(_09881_),
    .A2(_09884_),
    .A3(_09885_),
    .A4(_09892_),
    .B1(\fetch.bht.bhtTable_valid[12] ),
    .X(_00007_));
 sky130_fd_sc_hd__and2_2 _13514_ (.A(\csr.io_mem_pc[2] ),
    .B(\csr.io_mem_pc[3] ),
    .X(_09893_));
 sky130_fd_sc_hd__buf_1 _13515_ (.A(_09893_),
    .X(_09894_));
 sky130_fd_sc_hd__and4b_2 _13516_ (.A_N(_09879_),
    .B(_09882_),
    .C(\fetch.bht.bhtTable_tag_MPORT_en ),
    .D(_09894_),
    .X(_09895_));
 sky130_fd_sc_hd__buf_1 _13517_ (.A(_09895_),
    .X(_09896_));
 sky130_fd_sc_hd__buf_1 _13518_ (.A(_09896_),
    .X(_09897_));
 sky130_fd_sc_hd__buf_1 _13519_ (.A(_09897_),
    .X(_09898_));
 sky130_fd_sc_hd__or2_2 _13520_ (.A(\fetch.bht.bhtTable_valid[11] ),
    .B(_09898_),
    .X(_09899_));
 sky130_fd_sc_hd__buf_1 _13521_ (.A(_09899_),
    .X(_00006_));
 sky130_fd_sc_hd__inv_2 _13522_ (.A(\fetch.bht.bhtTable_tag_MPORT_en ),
    .Y(_09900_));
 sky130_fd_sc_hd__or4bb_2 _13523_ (.A(_09900_),
    .B(_09880_),
    .C_N(_09883_),
    .D_N(_09887_),
    .X(_09901_));
 sky130_fd_sc_hd__buf_1 _13524_ (.A(_09901_),
    .X(_09902_));
 sky130_fd_sc_hd__buf_1 _13525_ (.A(_09902_),
    .X(_09903_));
 sky130_fd_sc_hd__or2b_2 _13526_ (.A(\fetch.bht.bhtTable_valid[10] ),
    .B_N(_09903_),
    .X(_09904_));
 sky130_fd_sc_hd__buf_1 _13527_ (.A(_09904_),
    .X(_00005_));
 sky130_fd_sc_hd__or4bb_2 _13528_ (.A(_09900_),
    .B(_09880_),
    .C_N(_09883_),
    .D_N(_09890_),
    .X(_09905_));
 sky130_fd_sc_hd__buf_1 _13529_ (.A(_09905_),
    .X(_09906_));
 sky130_fd_sc_hd__buf_1 _13530_ (.A(_09906_),
    .X(_09907_));
 sky130_fd_sc_hd__or2b_2 _13531_ (.A(\fetch.bht.bhtTable_valid[9] ),
    .B_N(_09907_),
    .X(_09908_));
 sky130_fd_sc_hd__buf_1 _13532_ (.A(_09908_),
    .X(_00019_));
 sky130_fd_sc_hd__and4b_2 _13533_ (.A_N(_09879_),
    .B(_09882_),
    .C(\fetch.bht.bhtTable_tag_MPORT_en ),
    .D(_09892_),
    .X(_09909_));
 sky130_fd_sc_hd__buf_1 _13534_ (.A(_09909_),
    .X(_09910_));
 sky130_fd_sc_hd__buf_1 _13535_ (.A(_09910_),
    .X(_09911_));
 sky130_fd_sc_hd__buf_1 _13536_ (.A(_09911_),
    .X(_09912_));
 sky130_fd_sc_hd__or2_2 _13537_ (.A(\fetch.bht.bhtTable_valid[8] ),
    .B(_09912_),
    .X(_09913_));
 sky130_fd_sc_hd__buf_1 _13538_ (.A(_09913_),
    .X(_00018_));
 sky130_fd_sc_hd__buf_1 _13539_ (.A(_09885_),
    .X(_09914_));
 sky130_fd_sc_hd__and2b_2 _13540_ (.A_N(\csr.io_mem_pc[5] ),
    .B(_09879_),
    .X(_09915_));
 sky130_fd_sc_hd__buf_1 _13541_ (.A(_09915_),
    .X(_09916_));
 sky130_fd_sc_hd__a31o_2 _13542_ (.A1(_09914_),
    .A2(_09894_),
    .A3(_09916_),
    .B1(\fetch.bht.bhtTable_valid[7] ),
    .X(_00017_));
 sky130_fd_sc_hd__a31o_2 _13543_ (.A1(_09914_),
    .A2(_09887_),
    .A3(_09916_),
    .B1(\fetch.bht.bhtTable_valid[6] ),
    .X(_00016_));
 sky130_fd_sc_hd__a31o_2 _13544_ (.A1(_09914_),
    .A2(_09890_),
    .A3(_09916_),
    .B1(\fetch.bht.bhtTable_valid[5] ),
    .X(_00015_));
 sky130_fd_sc_hd__a31o_2 _13545_ (.A1(_09914_),
    .A2(_09892_),
    .A3(_09916_),
    .B1(\fetch.bht.bhtTable_valid[4] ),
    .X(_00014_));
 sky130_fd_sc_hd__nor2_2 _13546_ (.A(_09879_),
    .B(_09882_),
    .Y(_09917_));
 sky130_fd_sc_hd__a31o_2 _13547_ (.A1(_09914_),
    .A2(_09894_),
    .A3(_09917_),
    .B1(\fetch.bht.bhtTable_valid[3] ),
    .X(_00013_));
 sky130_fd_sc_hd__a31o_2 _13548_ (.A1(_09914_),
    .A2(_09887_),
    .A3(_09917_),
    .B1(\fetch.bht.bhtTable_valid[2] ),
    .X(_00012_));
 sky130_fd_sc_hd__a31o_2 _13549_ (.A1(_09914_),
    .A2(_09890_),
    .A3(_09917_),
    .B1(\fetch.bht.bhtTable_valid[1] ),
    .X(_00011_));
 sky130_fd_sc_hd__a31o_2 _13550_ (.A1(_09914_),
    .A2(_09892_),
    .A3(_09917_),
    .B1(\fetch.bht.bhtTable_valid[0] ),
    .X(_00004_));
 sky130_fd_sc_hd__nor2_2 _13551_ (.A(\execute.io_mem_rd[0] ),
    .B(\execute.io_mem_rd[1] ),
    .Y(_09918_));
 sky130_fd_sc_hd__nor2_2 _13552_ (.A(\execute.io_mem_rd[2] ),
    .B(\execute.io_mem_rd[3] ),
    .Y(_09919_));
 sky130_fd_sc_hd__inv_2 _13553_ (.A(\execute.io_mem_rd[4] ),
    .Y(_09920_));
 sky130_fd_sc_hd__nand3_2 _13554_ (.A(_09918_),
    .B(_09919_),
    .C(_09920_),
    .Y(_09921_));
 sky130_fd_sc_hd__o22a_2 _13555_ (.A1(io_memory_address[0]),
    .A2(io_memory_address[1]),
    .B1(io_memory_read),
    .B2(\execute.io_mem_memwrite ),
    .X(_09922_));
 sky130_fd_sc_hd__and3_2 _13556_ (.A(\csr.meie ),
    .B(\csr.ie ),
    .C(io_meip),
    .X(_09923_));
 sky130_fd_sc_hd__a31o_2 _13557_ (.A1(\csr.msie ),
    .A2(\csr.msip ),
    .A3(\csr.ie ),
    .B1(_09923_),
    .X(_09924_));
 sky130_fd_sc_hd__a311o_2 _13558_ (.A1(\csr.mtie ),
    .A2(\csr.ie ),
    .A3(\csr.mtip ),
    .B1(\execute.exception_out_reg ),
    .C1(_09924_),
    .X(_09925_));
 sky130_fd_sc_hd__a211oi_2 _13559_ (.A1(io_memory_read),
    .A2(_09921_),
    .B1(_09922_),
    .C1(_09925_),
    .Y(_09926_));
 sky130_fd_sc_hd__and2b_2 _13560_ (.A_N(_09926_),
    .B(\execute.io_mem_memwrite ),
    .X(_09927_));
 sky130_fd_sc_hd__buf_1 _13561_ (.A(_09927_),
    .X(io_memory_write));
 sky130_fd_sc_hd__and3_2 _13562_ (.A(\csr.io_mem_pc[4] ),
    .B(\csr.io_mem_pc[2] ),
    .C(\csr.io_mem_pc[3] ),
    .X(_09928_));
 sky130_fd_sc_hd__a31o_2 _13563_ (.A1(_09884_),
    .A2(_09914_),
    .A3(_09928_),
    .B1(\fetch.bht.bhtTable_valid[15] ),
    .X(_00010_));
 sky130_fd_sc_hd__buf_1 _13564_ (.A(\decode.io_wb_rd[2] ),
    .X(_09929_));
 sky130_fd_sc_hd__buf_1 _13565_ (.A(_09929_),
    .X(_09930_));
 sky130_fd_sc_hd__inv_2 _13566_ (.A(\decode.io_wb_rd[1] ),
    .Y(_09931_));
 sky130_fd_sc_hd__nor2_2 _13567_ (.A(\decode.io_wb_rd[0] ),
    .B(_09931_),
    .Y(_09932_));
 sky130_fd_sc_hd__and2_2 _13568_ (.A(\decode.io_wb_rd[4] ),
    .B(\decode.io_wb_regwrite ),
    .X(_09933_));
 sky130_fd_sc_hd__inv_2 _13569_ (.A(\decode.io_wb_rd[3] ),
    .Y(_09934_));
 sky130_fd_sc_hd__buf_1 _13570_ (.A(_09934_),
    .X(_09935_));
 sky130_fd_sc_hd__and4_2 _13571_ (.A(_09930_),
    .B(_09932_),
    .C(_09933_),
    .D(_09935_),
    .X(_09936_));
 sky130_fd_sc_hd__buf_1 _13572_ (.A(_09936_),
    .X(_09937_));
 sky130_fd_sc_hd__buf_1 _13573_ (.A(_09937_),
    .X(_09938_));
 sky130_fd_sc_hd__buf_1 _13574_ (.A(\memory.io_wb_memtoreg[1] ),
    .X(_09939_));
 sky130_fd_sc_hd__buf_1 _13575_ (.A(\memory.io_wb_memtoreg[0] ),
    .X(_09940_));
 sky130_fd_sc_hd__nand2_2 _13576_ (.A(_09939_),
    .B(_09940_),
    .Y(_09941_));
 sky130_fd_sc_hd__buf_1 _13577_ (.A(_09941_),
    .X(_09942_));
 sky130_fd_sc_hd__buf_1 _13578_ (.A(_09939_),
    .X(_09943_));
 sky130_fd_sc_hd__a21o_2 _13579_ (.A1(_09939_),
    .A2(\memory.io_wb_aluresult[0] ),
    .B1(_09940_),
    .X(_09944_));
 sky130_fd_sc_hd__o21ai_2 _13580_ (.A1(_09943_),
    .A2(\memory.io_wb_readdata[0] ),
    .B1(_09944_),
    .Y(_09945_));
 sky130_fd_sc_hd__nand2b_2 _13581_ (.A_N(_09939_),
    .B(_09940_),
    .Y(_09946_));
 sky130_fd_sc_hd__nand2b_2 _13582_ (.A_N(_09940_),
    .B(_09939_),
    .Y(_09947_));
 sky130_fd_sc_hd__nand3_2 _13583_ (.A(_09946_),
    .B(_09947_),
    .C(\memory.io_wb_reg_pc[0] ),
    .Y(_09948_));
 sky130_fd_sc_hd__a2bb2o_2 _13584_ (.A1_N(\memory.csr_read_data_out_reg[0] ),
    .A2_N(_09942_),
    .B1(_09945_),
    .B2(_09948_),
    .X(_09949_));
 sky130_fd_sc_hd__buf_1 _13585_ (.A(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__buf_1 _13586_ (.A(_09937_),
    .X(_09951_));
 sky130_fd_sc_hd__nand2_2 _13587_ (.A(_09950_),
    .B(_09951_),
    .Y(_09952_));
 sky130_fd_sc_hd__inv_2 _13588_ (.A(reset),
    .Y(_09953_));
 sky130_fd_sc_hd__buf_1 _13589_ (.A(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__buf_1 _13590_ (.A(_09954_),
    .X(_09955_));
 sky130_fd_sc_hd__buf_1 _13591_ (.A(_09955_),
    .X(_09956_));
 sky130_fd_sc_hd__buf_1 _13592_ (.A(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__o211a_2 _13593_ (.A1(\decode.regfile.registers_22[0] ),
    .A2(_09938_),
    .B1(_09952_),
    .C1(_09957_),
    .X(_00020_));
 sky130_fd_sc_hd__a21o_2 _13594_ (.A1(\memory.io_wb_memtoreg[1] ),
    .A2(\memory.io_wb_aluresult[1] ),
    .B1(\memory.io_wb_memtoreg[0] ),
    .X(_09958_));
 sky130_fd_sc_hd__o21a_2 _13595_ (.A1(\memory.io_wb_memtoreg[1] ),
    .A2(\memory.io_wb_readdata[1] ),
    .B1(_09958_),
    .X(_09959_));
 sky130_fd_sc_hd__and2_2 _13596_ (.A(\memory.io_wb_memtoreg[1] ),
    .B(\memory.io_wb_memtoreg[0] ),
    .X(_09960_));
 sky130_fd_sc_hd__nor2_2 _13597_ (.A(\memory.io_wb_memtoreg[1] ),
    .B(\memory.io_wb_memtoreg[0] ),
    .Y(_09961_));
 sky130_fd_sc_hd__o21a_2 _13598_ (.A1(_09960_),
    .A2(_09961_),
    .B1(\memory.io_wb_reg_pc[1] ),
    .X(_09962_));
 sky130_fd_sc_hd__o22ai_2 _13599_ (.A1(\memory.csr_read_data_out_reg[1] ),
    .A2(_09941_),
    .B1(_09959_),
    .B2(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__buf_1 _13600_ (.A(_09963_),
    .X(_09964_));
 sky130_fd_sc_hd__nand2_2 _13601_ (.A(_09964_),
    .B(_09951_),
    .Y(_09965_));
 sky130_fd_sc_hd__o211a_2 _13602_ (.A1(\decode.regfile.registers_22[1] ),
    .A2(_09938_),
    .B1(_09965_),
    .C1(_09957_),
    .X(_00021_));
 sky130_fd_sc_hd__a21o_2 _13603_ (.A1(_09939_),
    .A2(\memory.io_wb_aluresult[2] ),
    .B1(_09940_),
    .X(_09966_));
 sky130_fd_sc_hd__o21ai_2 _13604_ (.A1(_09939_),
    .A2(\memory.io_wb_readdata[2] ),
    .B1(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__o21ai_2 _13605_ (.A1(_09960_),
    .A2(_09961_),
    .B1(\memory.io_wb_reg_pc[2] ),
    .Y(_09968_));
 sky130_fd_sc_hd__a2bb2o_2 _13606_ (.A1_N(\memory.csr_read_data_out_reg[2] ),
    .A2_N(_09942_),
    .B1(_09967_),
    .B2(_09968_),
    .X(_09969_));
 sky130_fd_sc_hd__buf_1 _13607_ (.A(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__nand2_2 _13608_ (.A(_09970_),
    .B(_09951_),
    .Y(_09971_));
 sky130_fd_sc_hd__o211a_2 _13609_ (.A1(\decode.regfile.registers_22[2] ),
    .A2(_09938_),
    .B1(_09971_),
    .C1(_09957_),
    .X(_00022_));
 sky130_fd_sc_hd__and3b_2 _13610_ (.A_N(_09939_),
    .B(_09940_),
    .C(\memory.io_wb_readdata[3] ),
    .X(_09972_));
 sky130_fd_sc_hd__a221o_2 _13611_ (.A1(_09939_),
    .A2(\memory.io_wb_aluresult[3] ),
    .B1(_09961_),
    .B2(\memory.io_wb_reg_pc[3] ),
    .C1(_09960_),
    .X(_09973_));
 sky130_fd_sc_hd__o22ai_2 _13612_ (.A1(\memory.csr_read_data_out_reg[3] ),
    .A2(_09941_),
    .B1(_09972_),
    .B2(_09973_),
    .Y(_09974_));
 sky130_fd_sc_hd__buf_1 _13613_ (.A(_09974_),
    .X(_09975_));
 sky130_fd_sc_hd__nand2_2 _13614_ (.A(_09975_),
    .B(_09951_),
    .Y(_09976_));
 sky130_fd_sc_hd__o211a_2 _13615_ (.A1(\decode.regfile.registers_22[3] ),
    .A2(_09938_),
    .B1(_09976_),
    .C1(_09957_),
    .X(_00023_));
 sky130_fd_sc_hd__buf_1 _13616_ (.A(_09960_),
    .X(_09977_));
 sky130_fd_sc_hd__buf_1 _13617_ (.A(_09961_),
    .X(_09978_));
 sky130_fd_sc_hd__o21ai_2 _13618_ (.A1(_09977_),
    .A2(_09978_),
    .B1(\memory.io_wb_reg_pc[4] ),
    .Y(_09979_));
 sky130_fd_sc_hd__and2b_2 _13619_ (.A_N(\memory.io_wb_memtoreg[1] ),
    .B(_09940_),
    .X(_09980_));
 sky130_fd_sc_hd__buf_1 _13620_ (.A(_09980_),
    .X(_09981_));
 sky130_fd_sc_hd__a221oi_2 _13621_ (.A1(_09943_),
    .A2(\memory.io_wb_aluresult[4] ),
    .B1(_09981_),
    .B2(\memory.io_wb_readdata[4] ),
    .C1(_09977_),
    .Y(_09982_));
 sky130_fd_sc_hd__a2bb2o_2 _13622_ (.A1_N(\memory.csr_read_data_out_reg[4] ),
    .A2_N(_09942_),
    .B1(_09979_),
    .B2(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__buf_1 _13623_ (.A(_09983_),
    .X(_09984_));
 sky130_fd_sc_hd__nand2_2 _13624_ (.A(_09984_),
    .B(_09951_),
    .Y(_09985_));
 sky130_fd_sc_hd__o211a_2 _13625_ (.A1(\decode.regfile.registers_22[4] ),
    .A2(_09938_),
    .B1(_09985_),
    .C1(_09957_),
    .X(_00024_));
 sky130_fd_sc_hd__buf_1 _13626_ (.A(_09942_),
    .X(_09986_));
 sky130_fd_sc_hd__buf_1 _13627_ (.A(_09986_),
    .X(_09987_));
 sky130_fd_sc_hd__buf_1 _13628_ (.A(_09987_),
    .X(_09988_));
 sky130_fd_sc_hd__buf_1 _13629_ (.A(_09988_),
    .X(_09989_));
 sky130_fd_sc_hd__a22o_2 _13630_ (.A1(_09943_),
    .A2(\memory.io_wb_aluresult[5] ),
    .B1(_09980_),
    .B2(\memory.io_wb_readdata[5] ),
    .X(_09990_));
 sky130_fd_sc_hd__a211o_2 _13631_ (.A1(\memory.io_wb_reg_pc[5] ),
    .A2(_09978_),
    .B1(_09977_),
    .C1(_09990_),
    .X(_09991_));
 sky130_fd_sc_hd__o21ai_2 _13632_ (.A1(\memory.csr_read_data_out_reg[5] ),
    .A2(_09989_),
    .B1(_09991_),
    .Y(_09992_));
 sky130_fd_sc_hd__buf_1 _13633_ (.A(_09992_),
    .X(_09993_));
 sky130_fd_sc_hd__nand2_2 _13634_ (.A(_09993_),
    .B(_09951_),
    .Y(_09994_));
 sky130_fd_sc_hd__o211a_2 _13635_ (.A1(\decode.regfile.registers_22[5] ),
    .A2(_09938_),
    .B1(_09994_),
    .C1(_09957_),
    .X(_00025_));
 sky130_fd_sc_hd__buf_1 _13636_ (.A(_09977_),
    .X(_09995_));
 sky130_fd_sc_hd__a22o_2 _13637_ (.A1(_09943_),
    .A2(\memory.io_wb_aluresult[6] ),
    .B1(_09981_),
    .B2(\memory.io_wb_readdata[6] ),
    .X(_09996_));
 sky130_fd_sc_hd__a211o_2 _13638_ (.A1(\memory.io_wb_reg_pc[6] ),
    .A2(_09978_),
    .B1(_09995_),
    .C1(_09996_),
    .X(_09997_));
 sky130_fd_sc_hd__o21ai_2 _13639_ (.A1(\memory.csr_read_data_out_reg[6] ),
    .A2(_09989_),
    .B1(_09997_),
    .Y(_09998_));
 sky130_fd_sc_hd__buf_1 _13640_ (.A(_09998_),
    .X(_09999_));
 sky130_fd_sc_hd__nand2_2 _13641_ (.A(_09999_),
    .B(_09951_),
    .Y(_10000_));
 sky130_fd_sc_hd__o211a_2 _13642_ (.A1(\decode.regfile.registers_22[6] ),
    .A2(_09938_),
    .B1(_10000_),
    .C1(_09957_),
    .X(_00026_));
 sky130_fd_sc_hd__buf_1 _13643_ (.A(_09978_),
    .X(_10001_));
 sky130_fd_sc_hd__and2_2 _13644_ (.A(\memory.io_wb_reg_pc[7] ),
    .B(_10001_),
    .X(_10002_));
 sky130_fd_sc_hd__buf_1 _13645_ (.A(_09943_),
    .X(_10003_));
 sky130_fd_sc_hd__buf_1 _13646_ (.A(_09981_),
    .X(_10004_));
 sky130_fd_sc_hd__buf_1 _13647_ (.A(_09977_),
    .X(_10005_));
 sky130_fd_sc_hd__a221o_2 _13648_ (.A1(_10003_),
    .A2(\memory.io_wb_aluresult[7] ),
    .B1(_10004_),
    .B2(\memory.io_wb_readdata[7] ),
    .C1(_10005_),
    .X(_10006_));
 sky130_fd_sc_hd__o22ai_2 _13649_ (.A1(\memory.csr_read_data_out_reg[7] ),
    .A2(_09989_),
    .B1(_10002_),
    .B2(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__buf_1 _13650_ (.A(_10007_),
    .X(_10008_));
 sky130_fd_sc_hd__nand2_2 _13651_ (.A(_10008_),
    .B(_09951_),
    .Y(_10009_));
 sky130_fd_sc_hd__o211a_2 _13652_ (.A1(\decode.regfile.registers_22[7] ),
    .A2(_09938_),
    .B1(_10009_),
    .C1(_09957_),
    .X(_00027_));
 sky130_fd_sc_hd__buf_1 _13653_ (.A(_09942_),
    .X(_10010_));
 sky130_fd_sc_hd__o21ai_2 _13654_ (.A1(_09995_),
    .A2(_09978_),
    .B1(\memory.io_wb_reg_pc[8] ),
    .Y(_10011_));
 sky130_fd_sc_hd__buf_1 _13655_ (.A(_09943_),
    .X(_10012_));
 sky130_fd_sc_hd__a221oi_2 _13656_ (.A1(_10012_),
    .A2(\memory.io_wb_aluresult[8] ),
    .B1(_09981_),
    .B2(\memory.io_wb_readdata[8] ),
    .C1(_09995_),
    .Y(_10013_));
 sky130_fd_sc_hd__a2bb2o_2 _13657_ (.A1_N(\memory.csr_read_data_out_reg[8] ),
    .A2_N(_10010_),
    .B1(_10011_),
    .B2(_10013_),
    .X(_10014_));
 sky130_fd_sc_hd__buf_1 _13658_ (.A(_10014_),
    .X(_10015_));
 sky130_fd_sc_hd__buf_1 _13659_ (.A(_09937_),
    .X(_10016_));
 sky130_fd_sc_hd__nand2_2 _13660_ (.A(_10015_),
    .B(_10016_),
    .Y(_10017_));
 sky130_fd_sc_hd__buf_1 _13661_ (.A(_09954_),
    .X(_10018_));
 sky130_fd_sc_hd__buf_1 _13662_ (.A(_10018_),
    .X(_10019_));
 sky130_fd_sc_hd__buf_1 _13663_ (.A(_10019_),
    .X(_10020_));
 sky130_fd_sc_hd__o211a_2 _13664_ (.A1(\decode.regfile.registers_22[8] ),
    .A2(_09938_),
    .B1(_10017_),
    .C1(_10020_),
    .X(_00028_));
 sky130_fd_sc_hd__buf_1 _13665_ (.A(_09940_),
    .X(_10021_));
 sky130_fd_sc_hd__and3b_2 _13666_ (.A_N(_10012_),
    .B(_10021_),
    .C(\memory.io_wb_readdata[9] ),
    .X(_10022_));
 sky130_fd_sc_hd__a221o_2 _13667_ (.A1(_10012_),
    .A2(\memory.io_wb_aluresult[9] ),
    .B1(_09978_),
    .B2(\memory.io_wb_reg_pc[9] ),
    .C1(_09995_),
    .X(_10023_));
 sky130_fd_sc_hd__o22ai_2 _13668_ (.A1(\memory.csr_read_data_out_reg[9] ),
    .A2(_09988_),
    .B1(_10022_),
    .B2(_10023_),
    .Y(_10024_));
 sky130_fd_sc_hd__buf_1 _13669_ (.A(_10024_),
    .X(_10025_));
 sky130_fd_sc_hd__nand2_2 _13670_ (.A(_10025_),
    .B(_10016_),
    .Y(_10026_));
 sky130_fd_sc_hd__o211a_2 _13671_ (.A1(\decode.regfile.registers_22[9] ),
    .A2(_09938_),
    .B1(_10026_),
    .C1(_10020_),
    .X(_00029_));
 sky130_fd_sc_hd__buf_1 _13672_ (.A(_09937_),
    .X(_10027_));
 sky130_fd_sc_hd__and3_2 _13673_ (.A(_09946_),
    .B(_09947_),
    .C(\memory.io_wb_reg_pc[10] ),
    .X(_10028_));
 sky130_fd_sc_hd__a221o_2 _13674_ (.A1(_10012_),
    .A2(\memory.io_wb_aluresult[10] ),
    .B1(_09981_),
    .B2(\memory.io_wb_readdata[10] ),
    .C1(_09977_),
    .X(_10029_));
 sky130_fd_sc_hd__o22ai_2 _13675_ (.A1(\memory.csr_read_data_out_reg[10] ),
    .A2(_09988_),
    .B1(_10028_),
    .B2(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__buf_1 _13676_ (.A(_10030_),
    .X(_10031_));
 sky130_fd_sc_hd__nand2_2 _13677_ (.A(_10031_),
    .B(_10016_),
    .Y(_10032_));
 sky130_fd_sc_hd__o211a_2 _13678_ (.A1(\decode.regfile.registers_22[10] ),
    .A2(_10027_),
    .B1(_10032_),
    .C1(_10020_),
    .X(_00030_));
 sky130_fd_sc_hd__and3b_2 _13679_ (.A_N(_10012_),
    .B(_10021_),
    .C(\memory.io_wb_readdata[11] ),
    .X(_10033_));
 sky130_fd_sc_hd__a221o_2 _13680_ (.A1(_10012_),
    .A2(\memory.io_wb_aluresult[11] ),
    .B1(_09978_),
    .B2(\memory.io_wb_reg_pc[11] ),
    .C1(_09977_),
    .X(_10034_));
 sky130_fd_sc_hd__o22ai_2 _13681_ (.A1(\memory.csr_read_data_out_reg[11] ),
    .A2(_09988_),
    .B1(_10033_),
    .B2(_10034_),
    .Y(_10035_));
 sky130_fd_sc_hd__buf_1 _13682_ (.A(_10035_),
    .X(_10036_));
 sky130_fd_sc_hd__nand2_2 _13683_ (.A(_10036_),
    .B(_10016_),
    .Y(_10037_));
 sky130_fd_sc_hd__o211a_2 _13684_ (.A1(\decode.regfile.registers_22[11] ),
    .A2(_10027_),
    .B1(_10037_),
    .C1(_10020_),
    .X(_00031_));
 sky130_fd_sc_hd__a21o_2 _13685_ (.A1(_09939_),
    .A2(\memory.io_wb_aluresult[12] ),
    .B1(_09940_),
    .X(_10038_));
 sky130_fd_sc_hd__o21ai_2 _13686_ (.A1(_09943_),
    .A2(\memory.io_wb_readdata[12] ),
    .B1(_10038_),
    .Y(_10039_));
 sky130_fd_sc_hd__o21ai_2 _13687_ (.A1(_09977_),
    .A2(_09978_),
    .B1(\memory.io_wb_reg_pc[12] ),
    .Y(_10040_));
 sky130_fd_sc_hd__a2bb2o_2 _13688_ (.A1_N(\memory.csr_read_data_out_reg[12] ),
    .A2_N(_09989_),
    .B1(_10039_),
    .B2(_10040_),
    .X(_10041_));
 sky130_fd_sc_hd__buf_1 _13689_ (.A(_10041_),
    .X(_10042_));
 sky130_fd_sc_hd__nand2_2 _13690_ (.A(_10042_),
    .B(_10016_),
    .Y(_10043_));
 sky130_fd_sc_hd__o211a_2 _13691_ (.A1(\decode.regfile.registers_22[12] ),
    .A2(_10027_),
    .B1(_10043_),
    .C1(_10020_),
    .X(_00032_));
 sky130_fd_sc_hd__o21ai_2 _13692_ (.A1(_09977_),
    .A2(_09978_),
    .B1(\memory.io_wb_reg_pc[13] ),
    .Y(_10044_));
 sky130_fd_sc_hd__a22oi_2 _13693_ (.A1(_09943_),
    .A2(\memory.io_wb_aluresult[13] ),
    .B1(_09981_),
    .B2(\memory.io_wb_readdata[13] ),
    .Y(_10045_));
 sky130_fd_sc_hd__nor2_2 _13694_ (.A(\memory.csr_read_data_out_reg[13] ),
    .B(_09942_),
    .Y(_10046_));
 sky130_fd_sc_hd__a31o_2 _13695_ (.A1(_09989_),
    .A2(_10044_),
    .A3(_10045_),
    .B1(_10046_),
    .X(_10047_));
 sky130_fd_sc_hd__buf_1 _13696_ (.A(_10047_),
    .X(_10048_));
 sky130_fd_sc_hd__nand2_2 _13697_ (.A(_10048_),
    .B(_10016_),
    .Y(_10049_));
 sky130_fd_sc_hd__o211a_2 _13698_ (.A1(\decode.regfile.registers_22[13] ),
    .A2(_10027_),
    .B1(_10049_),
    .C1(_10020_),
    .X(_00033_));
 sky130_fd_sc_hd__o21a_2 _13699_ (.A1(_10021_),
    .A2(\memory.io_wb_aluresult[14] ),
    .B1(_10012_),
    .X(_10050_));
 sky130_fd_sc_hd__a221oi_2 _13700_ (.A1(_10021_),
    .A2(\memory.io_wb_readdata[14] ),
    .B1(_10001_),
    .B2(\memory.io_wb_reg_pc[14] ),
    .C1(_10050_),
    .Y(_10051_));
 sky130_fd_sc_hd__o21bai_2 _13701_ (.A1(\memory.csr_read_data_out_reg[14] ),
    .A2(_09989_),
    .B1_N(_10051_),
    .Y(_10052_));
 sky130_fd_sc_hd__buf_1 _13702_ (.A(_10052_),
    .X(_10053_));
 sky130_fd_sc_hd__nand2_2 _13703_ (.A(_10053_),
    .B(_10016_),
    .Y(_10054_));
 sky130_fd_sc_hd__o211a_2 _13704_ (.A1(\decode.regfile.registers_22[14] ),
    .A2(_10027_),
    .B1(_10054_),
    .C1(_10020_),
    .X(_00034_));
 sky130_fd_sc_hd__nand2_2 _13705_ (.A(\memory.io_wb_readdata[15] ),
    .B(_09981_),
    .Y(_10055_));
 sky130_fd_sc_hd__a221oi_2 _13706_ (.A1(_10012_),
    .A2(\memory.io_wb_aluresult[15] ),
    .B1(_09978_),
    .B2(\memory.io_wb_reg_pc[15] ),
    .C1(_09995_),
    .Y(_10056_));
 sky130_fd_sc_hd__a2bb2o_2 _13707_ (.A1_N(\memory.csr_read_data_out_reg[15] ),
    .A2_N(_09989_),
    .B1(_10055_),
    .B2(_10056_),
    .X(_10057_));
 sky130_fd_sc_hd__buf_1 _13708_ (.A(_10057_),
    .X(_10058_));
 sky130_fd_sc_hd__nand2_2 _13709_ (.A(_10058_),
    .B(_10016_),
    .Y(_10059_));
 sky130_fd_sc_hd__o211a_2 _13710_ (.A1(\decode.regfile.registers_22[15] ),
    .A2(_10027_),
    .B1(_10059_),
    .C1(_10020_),
    .X(_00035_));
 sky130_fd_sc_hd__buf_1 _13711_ (.A(_10003_),
    .X(_10060_));
 sky130_fd_sc_hd__and3b_2 _13712_ (.A_N(_10060_),
    .B(_10021_),
    .C(\memory.io_wb_readdata[16] ),
    .X(_10061_));
 sky130_fd_sc_hd__a221o_2 _13713_ (.A1(_10003_),
    .A2(\memory.io_wb_aluresult[16] ),
    .B1(_10001_),
    .B2(\memory.io_wb_reg_pc[16] ),
    .C1(_10005_),
    .X(_10062_));
 sky130_fd_sc_hd__o22ai_2 _13714_ (.A1(\memory.csr_read_data_out_reg[16] ),
    .A2(_09987_),
    .B1(_10061_),
    .B2(_10062_),
    .Y(_10063_));
 sky130_fd_sc_hd__buf_1 _13715_ (.A(_10063_),
    .X(_10064_));
 sky130_fd_sc_hd__nand2_2 _13716_ (.A(_10064_),
    .B(_10016_),
    .Y(_10065_));
 sky130_fd_sc_hd__o211a_2 _13717_ (.A1(\decode.regfile.registers_22[16] ),
    .A2(_10027_),
    .B1(_10065_),
    .C1(_10020_),
    .X(_00036_));
 sky130_fd_sc_hd__or3b_2 _13718_ (.A(_10012_),
    .B(_10021_),
    .C_N(\memory.io_wb_reg_pc[17] ),
    .X(_10066_));
 sky130_fd_sc_hd__a221oi_2 _13719_ (.A1(_10003_),
    .A2(\memory.io_wb_aluresult[17] ),
    .B1(_10004_),
    .B2(\memory.io_wb_readdata[17] ),
    .C1(_09995_),
    .Y(_10067_));
 sky130_fd_sc_hd__a2bb2o_2 _13720_ (.A1_N(\memory.csr_read_data_out_reg[17] ),
    .A2_N(_09986_),
    .B1(_10066_),
    .B2(_10067_),
    .X(_10068_));
 sky130_fd_sc_hd__buf_1 _13721_ (.A(_10068_),
    .X(_10069_));
 sky130_fd_sc_hd__nand2_2 _13722_ (.A(_10069_),
    .B(_10016_),
    .Y(_10070_));
 sky130_fd_sc_hd__o211a_2 _13723_ (.A1(\decode.regfile.registers_22[17] ),
    .A2(_10027_),
    .B1(_10070_),
    .C1(_10020_),
    .X(_00037_));
 sky130_fd_sc_hd__o21ai_2 _13724_ (.A1(_10005_),
    .A2(_10001_),
    .B1(\memory.io_wb_reg_pc[18] ),
    .Y(_10071_));
 sky130_fd_sc_hd__a221oi_2 _13725_ (.A1(_10003_),
    .A2(\memory.io_wb_aluresult[18] ),
    .B1(_10004_),
    .B2(\memory.io_wb_readdata[18] ),
    .C1(_10005_),
    .Y(_10072_));
 sky130_fd_sc_hd__a2bb2o_2 _13726_ (.A1_N(\memory.csr_read_data_out_reg[18] ),
    .A2_N(_09986_),
    .B1(_10071_),
    .B2(_10072_),
    .X(_10073_));
 sky130_fd_sc_hd__buf_1 _13727_ (.A(_10073_),
    .X(_10074_));
 sky130_fd_sc_hd__buf_1 _13728_ (.A(_09937_),
    .X(_10075_));
 sky130_fd_sc_hd__nand2_2 _13729_ (.A(_10074_),
    .B(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__buf_1 _13730_ (.A(_10019_),
    .X(_10077_));
 sky130_fd_sc_hd__o211a_2 _13731_ (.A1(\decode.regfile.registers_22[18] ),
    .A2(_10027_),
    .B1(_10076_),
    .C1(_10077_),
    .X(_00038_));
 sky130_fd_sc_hd__and3b_2 _13732_ (.A_N(_10003_),
    .B(_10021_),
    .C(\memory.io_wb_readdata[19] ),
    .X(_10078_));
 sky130_fd_sc_hd__a221o_2 _13733_ (.A1(_10003_),
    .A2(\memory.io_wb_aluresult[19] ),
    .B1(_10001_),
    .B2(\memory.io_wb_reg_pc[19] ),
    .C1(_09995_),
    .X(_10079_));
 sky130_fd_sc_hd__o22ai_2 _13734_ (.A1(\memory.csr_read_data_out_reg[19] ),
    .A2(_09986_),
    .B1(_10078_),
    .B2(_10079_),
    .Y(_10080_));
 sky130_fd_sc_hd__buf_1 _13735_ (.A(_10080_),
    .X(_10081_));
 sky130_fd_sc_hd__nand2_2 _13736_ (.A(_10081_),
    .B(_10075_),
    .Y(_10082_));
 sky130_fd_sc_hd__o211a_2 _13737_ (.A1(\decode.regfile.registers_22[19] ),
    .A2(_10027_),
    .B1(_10082_),
    .C1(_10077_),
    .X(_00039_));
 sky130_fd_sc_hd__buf_1 _13738_ (.A(_09937_),
    .X(_10083_));
 sky130_fd_sc_hd__a221o_2 _13739_ (.A1(_09943_),
    .A2(\memory.io_wb_aluresult[20] ),
    .B1(_09981_),
    .B2(\memory.io_wb_readdata[20] ),
    .C1(_09977_),
    .X(_10084_));
 sky130_fd_sc_hd__a31o_2 _13740_ (.A1(\memory.io_wb_reg_pc[20] ),
    .A2(_09946_),
    .A3(_09947_),
    .B1(_10084_),
    .X(_10085_));
 sky130_fd_sc_hd__o21ai_2 _13741_ (.A1(\memory.csr_read_data_out_reg[20] ),
    .A2(_10010_),
    .B1(_10085_),
    .Y(_10086_));
 sky130_fd_sc_hd__buf_1 _13742_ (.A(_10086_),
    .X(_10087_));
 sky130_fd_sc_hd__nand2_2 _13743_ (.A(_10087_),
    .B(_10075_),
    .Y(_10088_));
 sky130_fd_sc_hd__o211a_2 _13744_ (.A1(\decode.regfile.registers_22[20] ),
    .A2(_10083_),
    .B1(_10088_),
    .C1(_10077_),
    .X(_00040_));
 sky130_fd_sc_hd__or3b_2 _13745_ (.A(_09943_),
    .B(_09940_),
    .C_N(\memory.io_wb_reg_pc[21] ),
    .X(_10089_));
 sky130_fd_sc_hd__a221oi_2 _13746_ (.A1(_10012_),
    .A2(\memory.io_wb_aluresult[21] ),
    .B1(_09981_),
    .B2(\memory.io_wb_readdata[21] ),
    .C1(_09995_),
    .Y(_10090_));
 sky130_fd_sc_hd__a2bb2o_2 _13747_ (.A1_N(\memory.csr_read_data_out_reg[21] ),
    .A2_N(_09987_),
    .B1(_10089_),
    .B2(_10090_),
    .X(_10091_));
 sky130_fd_sc_hd__buf_1 _13748_ (.A(_10091_),
    .X(_10092_));
 sky130_fd_sc_hd__nand2_2 _13749_ (.A(_10092_),
    .B(_10075_),
    .Y(_10093_));
 sky130_fd_sc_hd__o211a_2 _13750_ (.A1(\decode.regfile.registers_22[21] ),
    .A2(_10083_),
    .B1(_10093_),
    .C1(_10077_),
    .X(_00041_));
 sky130_fd_sc_hd__a221o_2 _13751_ (.A1(_10003_),
    .A2(\memory.io_wb_aluresult[22] ),
    .B1(_09981_),
    .B2(\memory.io_wb_readdata[22] ),
    .C1(_09995_),
    .X(_10094_));
 sky130_fd_sc_hd__a31o_2 _13752_ (.A1(\memory.io_wb_reg_pc[22] ),
    .A2(_09946_),
    .A3(_09947_),
    .B1(_10094_),
    .X(_10095_));
 sky130_fd_sc_hd__o21ai_2 _13753_ (.A1(\memory.csr_read_data_out_reg[22] ),
    .A2(_09989_),
    .B1(_10095_),
    .Y(_10096_));
 sky130_fd_sc_hd__buf_1 _13754_ (.A(_10096_),
    .X(_10097_));
 sky130_fd_sc_hd__nand2_2 _13755_ (.A(_10097_),
    .B(_10075_),
    .Y(_10098_));
 sky130_fd_sc_hd__o211a_2 _13756_ (.A1(\decode.regfile.registers_22[22] ),
    .A2(_10083_),
    .B1(_10098_),
    .C1(_10077_),
    .X(_00042_));
 sky130_fd_sc_hd__and3b_2 _13757_ (.A_N(_10003_),
    .B(_10021_),
    .C(\memory.io_wb_readdata[23] ),
    .X(_10099_));
 sky130_fd_sc_hd__a221o_2 _13758_ (.A1(_10003_),
    .A2(\memory.io_wb_aluresult[23] ),
    .B1(_10001_),
    .B2(\memory.io_wb_reg_pc[23] ),
    .C1(_09995_),
    .X(_10100_));
 sky130_fd_sc_hd__o22ai_2 _13759_ (.A1(\memory.csr_read_data_out_reg[23] ),
    .A2(_09986_),
    .B1(_10099_),
    .B2(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__buf_1 _13760_ (.A(_10101_),
    .X(_10102_));
 sky130_fd_sc_hd__nand2_2 _13761_ (.A(_10102_),
    .B(_10075_),
    .Y(_10103_));
 sky130_fd_sc_hd__o211a_2 _13762_ (.A1(\decode.regfile.registers_22[23] ),
    .A2(_10083_),
    .B1(_10103_),
    .C1(_10077_),
    .X(_00043_));
 sky130_fd_sc_hd__and2_2 _13763_ (.A(\memory.io_wb_reg_pc[24] ),
    .B(_10001_),
    .X(_10104_));
 sky130_fd_sc_hd__a221o_2 _13764_ (.A1(_10060_),
    .A2(\memory.io_wb_aluresult[24] ),
    .B1(_10004_),
    .B2(\memory.io_wb_readdata[24] ),
    .C1(_10005_),
    .X(_10105_));
 sky130_fd_sc_hd__o22ai_2 _13765_ (.A1(\memory.csr_read_data_out_reg[24] ),
    .A2(_09988_),
    .B1(_10104_),
    .B2(_10105_),
    .Y(_10106_));
 sky130_fd_sc_hd__buf_1 _13766_ (.A(_10106_),
    .X(_10107_));
 sky130_fd_sc_hd__nand2_2 _13767_ (.A(_10107_),
    .B(_10075_),
    .Y(_10108_));
 sky130_fd_sc_hd__o211a_2 _13768_ (.A1(\decode.regfile.registers_22[24] ),
    .A2(_10083_),
    .B1(_10108_),
    .C1(_10077_),
    .X(_00044_));
 sky130_fd_sc_hd__a22o_2 _13769_ (.A1(_10060_),
    .A2(\memory.io_wb_aluresult[25] ),
    .B1(_10004_),
    .B2(\memory.io_wb_readdata[25] ),
    .X(_10109_));
 sky130_fd_sc_hd__a211o_2 _13770_ (.A1(\memory.io_wb_reg_pc[25] ),
    .A2(_10001_),
    .B1(_10005_),
    .C1(_10109_),
    .X(_10110_));
 sky130_fd_sc_hd__o21ai_2 _13771_ (.A1(\memory.csr_read_data_out_reg[25] ),
    .A2(_09989_),
    .B1(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__buf_1 _13772_ (.A(_10111_),
    .X(_10112_));
 sky130_fd_sc_hd__nand2_2 _13773_ (.A(_10112_),
    .B(_10075_),
    .Y(_10113_));
 sky130_fd_sc_hd__o211a_2 _13774_ (.A1(\decode.regfile.registers_22[25] ),
    .A2(_10083_),
    .B1(_10113_),
    .C1(_10077_),
    .X(_00045_));
 sky130_fd_sc_hd__a221o_2 _13775_ (.A1(_10060_),
    .A2(\memory.io_wb_aluresult[26] ),
    .B1(_10004_),
    .B2(\memory.io_wb_readdata[26] ),
    .C1(_10005_),
    .X(_10114_));
 sky130_fd_sc_hd__a31o_2 _13776_ (.A1(\memory.io_wb_reg_pc[26] ),
    .A2(_09946_),
    .A3(_09947_),
    .B1(_10114_),
    .X(_10115_));
 sky130_fd_sc_hd__o21ai_2 _13777_ (.A1(\memory.csr_read_data_out_reg[26] ),
    .A2(_09987_),
    .B1(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__buf_1 _13778_ (.A(_10116_),
    .X(_10117_));
 sky130_fd_sc_hd__nand2_2 _13779_ (.A(_10117_),
    .B(_10075_),
    .Y(_10118_));
 sky130_fd_sc_hd__o211a_2 _13780_ (.A1(\decode.regfile.registers_22[26] ),
    .A2(_10083_),
    .B1(_10118_),
    .C1(_10077_),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_2 _13781_ (.A1(_10060_),
    .A2(\memory.io_wb_aluresult[27] ),
    .B1(_10004_),
    .B2(\memory.io_wb_readdata[27] ),
    .X(_10119_));
 sky130_fd_sc_hd__a211o_2 _13782_ (.A1(\memory.io_wb_reg_pc[27] ),
    .A2(_10001_),
    .B1(_10005_),
    .C1(_10119_),
    .X(_10120_));
 sky130_fd_sc_hd__o21ai_2 _13783_ (.A1(\memory.csr_read_data_out_reg[27] ),
    .A2(_09987_),
    .B1(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__buf_1 _13784_ (.A(_10121_),
    .X(_10122_));
 sky130_fd_sc_hd__nand2_2 _13785_ (.A(_10122_),
    .B(_10075_),
    .Y(_10123_));
 sky130_fd_sc_hd__o211a_2 _13786_ (.A1(\decode.regfile.registers_22[27] ),
    .A2(_10083_),
    .B1(_10123_),
    .C1(_10077_),
    .X(_00047_));
 sky130_fd_sc_hd__a21o_2 _13787_ (.A1(_10060_),
    .A2(\memory.io_wb_aluresult[28] ),
    .B1(_10021_),
    .X(_10124_));
 sky130_fd_sc_hd__o21a_2 _13788_ (.A1(_10060_),
    .A2(\memory.io_wb_readdata[28] ),
    .B1(_10124_),
    .X(_10125_));
 sky130_fd_sc_hd__a31o_2 _13789_ (.A1(\memory.io_wb_reg_pc[28] ),
    .A2(_09946_),
    .A3(_09947_),
    .B1(_10125_),
    .X(_10126_));
 sky130_fd_sc_hd__o21ai_2 _13790_ (.A1(\memory.csr_read_data_out_reg[28] ),
    .A2(_09988_),
    .B1(_10126_),
    .Y(_10127_));
 sky130_fd_sc_hd__buf_1 _13791_ (.A(_10127_),
    .X(_10128_));
 sky130_fd_sc_hd__nand2_2 _13792_ (.A(_10128_),
    .B(_09937_),
    .Y(_10129_));
 sky130_fd_sc_hd__buf_1 _13793_ (.A(_09954_),
    .X(_10130_));
 sky130_fd_sc_hd__buf_1 _13794_ (.A(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__buf_1 _13795_ (.A(_10131_),
    .X(_10132_));
 sky130_fd_sc_hd__o211a_2 _13796_ (.A1(\decode.regfile.registers_22[28] ),
    .A2(_10083_),
    .B1(_10129_),
    .C1(_10132_),
    .X(_00048_));
 sky130_fd_sc_hd__a221o_2 _13797_ (.A1(_10060_),
    .A2(\memory.io_wb_aluresult[29] ),
    .B1(_10004_),
    .B2(\memory.io_wb_readdata[29] ),
    .C1(_10005_),
    .X(_10133_));
 sky130_fd_sc_hd__a31o_2 _13798_ (.A1(\memory.io_wb_reg_pc[29] ),
    .A2(_09946_),
    .A3(_09947_),
    .B1(_10133_),
    .X(_10134_));
 sky130_fd_sc_hd__o21ai_2 _13799_ (.A1(\memory.csr_read_data_out_reg[29] ),
    .A2(_09988_),
    .B1(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__buf_1 _13800_ (.A(_10135_),
    .X(_10136_));
 sky130_fd_sc_hd__nand2_2 _13801_ (.A(_10136_),
    .B(_09937_),
    .Y(_10137_));
 sky130_fd_sc_hd__o211a_2 _13802_ (.A1(\decode.regfile.registers_22[29] ),
    .A2(_10083_),
    .B1(_10137_),
    .C1(_10132_),
    .X(_00049_));
 sky130_fd_sc_hd__and2b_2 _13803_ (.A_N(_10021_),
    .B(\memory.io_wb_reg_pc[30] ),
    .X(_10138_));
 sky130_fd_sc_hd__o22a_2 _13804_ (.A1(_10060_),
    .A2(_10138_),
    .B1(_09947_),
    .B2(\memory.io_wb_aluresult[30] ),
    .X(_10139_));
 sky130_fd_sc_hd__a21o_2 _13805_ (.A1(\memory.io_wb_readdata[30] ),
    .A2(_10004_),
    .B1(_10139_),
    .X(_10140_));
 sky130_fd_sc_hd__o21ai_2 _13806_ (.A1(\memory.csr_read_data_out_reg[30] ),
    .A2(_09989_),
    .B1(_10140_),
    .Y(_10141_));
 sky130_fd_sc_hd__buf_1 _13807_ (.A(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__nand2_2 _13808_ (.A(_10142_),
    .B(_09937_),
    .Y(_10143_));
 sky130_fd_sc_hd__o211a_2 _13809_ (.A1(\decode.regfile.registers_22[30] ),
    .A2(_09951_),
    .B1(_10143_),
    .C1(_10132_),
    .X(_00050_));
 sky130_fd_sc_hd__and2_2 _13810_ (.A(\memory.io_wb_reg_pc[31] ),
    .B(_10001_),
    .X(_10144_));
 sky130_fd_sc_hd__a221o_2 _13811_ (.A1(_10060_),
    .A2(\memory.io_wb_aluresult[31] ),
    .B1(_10004_),
    .B2(\memory.io_wb_readdata[31] ),
    .C1(_10005_),
    .X(_10145_));
 sky130_fd_sc_hd__o22ai_2 _13812_ (.A1(\memory.csr_read_data_out_reg[31] ),
    .A2(_09988_),
    .B1(_10144_),
    .B2(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__buf_1 _13813_ (.A(_10146_),
    .X(_10147_));
 sky130_fd_sc_hd__nand2_2 _13814_ (.A(_10147_),
    .B(_09937_),
    .Y(_10148_));
 sky130_fd_sc_hd__o211a_2 _13815_ (.A1(\decode.regfile.registers_22[31] ),
    .A2(_09951_),
    .B1(_10148_),
    .C1(_10132_),
    .X(_00051_));
 sky130_fd_sc_hd__buf_1 _13816_ (.A(_09933_),
    .X(_10149_));
 sky130_fd_sc_hd__and2_2 _13817_ (.A(\decode.io_wb_rd[0] ),
    .B(\decode.io_wb_rd[1] ),
    .X(_10150_));
 sky130_fd_sc_hd__and4_2 _13818_ (.A(_09930_),
    .B(_10149_),
    .C(_10150_),
    .D(_09935_),
    .X(_10151_));
 sky130_fd_sc_hd__buf_1 _13819_ (.A(_10151_),
    .X(_10152_));
 sky130_fd_sc_hd__buf_1 _13820_ (.A(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__buf_1 _13821_ (.A(_10152_),
    .X(_10154_));
 sky130_fd_sc_hd__nand2_2 _13822_ (.A(_09950_),
    .B(_10154_),
    .Y(_10155_));
 sky130_fd_sc_hd__o211a_2 _13823_ (.A1(\decode.regfile.registers_23[0] ),
    .A2(_10153_),
    .B1(_10155_),
    .C1(_10132_),
    .X(_00052_));
 sky130_fd_sc_hd__nand2_2 _13824_ (.A(_09964_),
    .B(_10154_),
    .Y(_10156_));
 sky130_fd_sc_hd__o211a_2 _13825_ (.A1(\decode.regfile.registers_23[1] ),
    .A2(_10153_),
    .B1(_10156_),
    .C1(_10132_),
    .X(_00053_));
 sky130_fd_sc_hd__nand2_2 _13826_ (.A(_09970_),
    .B(_10154_),
    .Y(_10157_));
 sky130_fd_sc_hd__o211a_2 _13827_ (.A1(\decode.regfile.registers_23[2] ),
    .A2(_10153_),
    .B1(_10157_),
    .C1(_10132_),
    .X(_00054_));
 sky130_fd_sc_hd__nand2_2 _13828_ (.A(_09975_),
    .B(_10154_),
    .Y(_10158_));
 sky130_fd_sc_hd__o211a_2 _13829_ (.A1(\decode.regfile.registers_23[3] ),
    .A2(_10153_),
    .B1(_10158_),
    .C1(_10132_),
    .X(_00055_));
 sky130_fd_sc_hd__nand2_2 _13830_ (.A(_09984_),
    .B(_10154_),
    .Y(_10159_));
 sky130_fd_sc_hd__o211a_2 _13831_ (.A1(\decode.regfile.registers_23[4] ),
    .A2(_10153_),
    .B1(_10159_),
    .C1(_10132_),
    .X(_00056_));
 sky130_fd_sc_hd__nand2_2 _13832_ (.A(_09993_),
    .B(_10154_),
    .Y(_10160_));
 sky130_fd_sc_hd__o211a_2 _13833_ (.A1(\decode.regfile.registers_23[5] ),
    .A2(_10153_),
    .B1(_10160_),
    .C1(_10132_),
    .X(_00057_));
 sky130_fd_sc_hd__nand2_2 _13834_ (.A(_09999_),
    .B(_10154_),
    .Y(_10161_));
 sky130_fd_sc_hd__buf_1 _13835_ (.A(_10131_),
    .X(_10162_));
 sky130_fd_sc_hd__o211a_2 _13836_ (.A1(\decode.regfile.registers_23[6] ),
    .A2(_10153_),
    .B1(_10161_),
    .C1(_10162_),
    .X(_00058_));
 sky130_fd_sc_hd__nand2_2 _13837_ (.A(_10008_),
    .B(_10154_),
    .Y(_10163_));
 sky130_fd_sc_hd__o211a_2 _13838_ (.A1(\decode.regfile.registers_23[7] ),
    .A2(_10153_),
    .B1(_10163_),
    .C1(_10162_),
    .X(_00059_));
 sky130_fd_sc_hd__buf_1 _13839_ (.A(_10152_),
    .X(_10164_));
 sky130_fd_sc_hd__nand2_2 _13840_ (.A(_10015_),
    .B(_10164_),
    .Y(_10165_));
 sky130_fd_sc_hd__o211a_2 _13841_ (.A1(\decode.regfile.registers_23[8] ),
    .A2(_10153_),
    .B1(_10165_),
    .C1(_10162_),
    .X(_00060_));
 sky130_fd_sc_hd__nand2_2 _13842_ (.A(_10025_),
    .B(_10164_),
    .Y(_10166_));
 sky130_fd_sc_hd__o211a_2 _13843_ (.A1(\decode.regfile.registers_23[9] ),
    .A2(_10153_),
    .B1(_10166_),
    .C1(_10162_),
    .X(_00061_));
 sky130_fd_sc_hd__buf_1 _13844_ (.A(_10152_),
    .X(_10167_));
 sky130_fd_sc_hd__nand2_2 _13845_ (.A(_10031_),
    .B(_10164_),
    .Y(_10168_));
 sky130_fd_sc_hd__o211a_2 _13846_ (.A1(\decode.regfile.registers_23[10] ),
    .A2(_10167_),
    .B1(_10168_),
    .C1(_10162_),
    .X(_00062_));
 sky130_fd_sc_hd__nand2_2 _13847_ (.A(_10036_),
    .B(_10164_),
    .Y(_10169_));
 sky130_fd_sc_hd__o211a_2 _13848_ (.A1(\decode.regfile.registers_23[11] ),
    .A2(_10167_),
    .B1(_10169_),
    .C1(_10162_),
    .X(_00063_));
 sky130_fd_sc_hd__nand2_2 _13849_ (.A(_10042_),
    .B(_10164_),
    .Y(_10170_));
 sky130_fd_sc_hd__o211a_2 _13850_ (.A1(\decode.regfile.registers_23[12] ),
    .A2(_10167_),
    .B1(_10170_),
    .C1(_10162_),
    .X(_00064_));
 sky130_fd_sc_hd__nand2_2 _13851_ (.A(_10048_),
    .B(_10164_),
    .Y(_10171_));
 sky130_fd_sc_hd__o211a_2 _13852_ (.A1(\decode.regfile.registers_23[13] ),
    .A2(_10167_),
    .B1(_10171_),
    .C1(_10162_),
    .X(_00065_));
 sky130_fd_sc_hd__nand2_2 _13853_ (.A(_10053_),
    .B(_10164_),
    .Y(_10172_));
 sky130_fd_sc_hd__o211a_2 _13854_ (.A1(\decode.regfile.registers_23[14] ),
    .A2(_10167_),
    .B1(_10172_),
    .C1(_10162_),
    .X(_00066_));
 sky130_fd_sc_hd__nand2_2 _13855_ (.A(_10058_),
    .B(_10164_),
    .Y(_10173_));
 sky130_fd_sc_hd__o211a_2 _13856_ (.A1(\decode.regfile.registers_23[15] ),
    .A2(_10167_),
    .B1(_10173_),
    .C1(_10162_),
    .X(_00067_));
 sky130_fd_sc_hd__nand2_2 _13857_ (.A(_10064_),
    .B(_10164_),
    .Y(_10174_));
 sky130_fd_sc_hd__buf_1 _13858_ (.A(_10131_),
    .X(_10175_));
 sky130_fd_sc_hd__o211a_2 _13859_ (.A1(\decode.regfile.registers_23[16] ),
    .A2(_10167_),
    .B1(_10174_),
    .C1(_10175_),
    .X(_00068_));
 sky130_fd_sc_hd__nand2_2 _13860_ (.A(_10069_),
    .B(_10164_),
    .Y(_10176_));
 sky130_fd_sc_hd__o211a_2 _13861_ (.A1(\decode.regfile.registers_23[17] ),
    .A2(_10167_),
    .B1(_10176_),
    .C1(_10175_),
    .X(_00069_));
 sky130_fd_sc_hd__buf_1 _13862_ (.A(_10152_),
    .X(_10177_));
 sky130_fd_sc_hd__nand2_2 _13863_ (.A(_10074_),
    .B(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__o211a_2 _13864_ (.A1(\decode.regfile.registers_23[18] ),
    .A2(_10167_),
    .B1(_10178_),
    .C1(_10175_),
    .X(_00070_));
 sky130_fd_sc_hd__nand2_2 _13865_ (.A(_10081_),
    .B(_10177_),
    .Y(_10179_));
 sky130_fd_sc_hd__o211a_2 _13866_ (.A1(\decode.regfile.registers_23[19] ),
    .A2(_10167_),
    .B1(_10179_),
    .C1(_10175_),
    .X(_00071_));
 sky130_fd_sc_hd__buf_1 _13867_ (.A(_10152_),
    .X(_10180_));
 sky130_fd_sc_hd__nand2_2 _13868_ (.A(_10087_),
    .B(_10177_),
    .Y(_10181_));
 sky130_fd_sc_hd__o211a_2 _13869_ (.A1(\decode.regfile.registers_23[20] ),
    .A2(_10180_),
    .B1(_10181_),
    .C1(_10175_),
    .X(_00072_));
 sky130_fd_sc_hd__nand2_2 _13870_ (.A(_10092_),
    .B(_10177_),
    .Y(_10182_));
 sky130_fd_sc_hd__o211a_2 _13871_ (.A1(\decode.regfile.registers_23[21] ),
    .A2(_10180_),
    .B1(_10182_),
    .C1(_10175_),
    .X(_00073_));
 sky130_fd_sc_hd__nand2_2 _13872_ (.A(_10097_),
    .B(_10177_),
    .Y(_10183_));
 sky130_fd_sc_hd__o211a_2 _13873_ (.A1(\decode.regfile.registers_23[22] ),
    .A2(_10180_),
    .B1(_10183_),
    .C1(_10175_),
    .X(_00074_));
 sky130_fd_sc_hd__nand2_2 _13874_ (.A(_10102_),
    .B(_10177_),
    .Y(_10184_));
 sky130_fd_sc_hd__o211a_2 _13875_ (.A1(\decode.regfile.registers_23[23] ),
    .A2(_10180_),
    .B1(_10184_),
    .C1(_10175_),
    .X(_00075_));
 sky130_fd_sc_hd__nand2_2 _13876_ (.A(_10107_),
    .B(_10177_),
    .Y(_10185_));
 sky130_fd_sc_hd__o211a_2 _13877_ (.A1(\decode.regfile.registers_23[24] ),
    .A2(_10180_),
    .B1(_10185_),
    .C1(_10175_),
    .X(_00076_));
 sky130_fd_sc_hd__nand2_2 _13878_ (.A(_10112_),
    .B(_10177_),
    .Y(_10186_));
 sky130_fd_sc_hd__o211a_2 _13879_ (.A1(\decode.regfile.registers_23[25] ),
    .A2(_10180_),
    .B1(_10186_),
    .C1(_10175_),
    .X(_00077_));
 sky130_fd_sc_hd__nand2_2 _13880_ (.A(_10117_),
    .B(_10177_),
    .Y(_10187_));
 sky130_fd_sc_hd__buf_1 _13881_ (.A(_10131_),
    .X(_10188_));
 sky130_fd_sc_hd__o211a_2 _13882_ (.A1(\decode.regfile.registers_23[26] ),
    .A2(_10180_),
    .B1(_10187_),
    .C1(_10188_),
    .X(_00078_));
 sky130_fd_sc_hd__nand2_2 _13883_ (.A(_10122_),
    .B(_10177_),
    .Y(_10189_));
 sky130_fd_sc_hd__o211a_2 _13884_ (.A1(\decode.regfile.registers_23[27] ),
    .A2(_10180_),
    .B1(_10189_),
    .C1(_10188_),
    .X(_00079_));
 sky130_fd_sc_hd__nand2_2 _13885_ (.A(_10128_),
    .B(_10152_),
    .Y(_10190_));
 sky130_fd_sc_hd__o211a_2 _13886_ (.A1(\decode.regfile.registers_23[28] ),
    .A2(_10180_),
    .B1(_10190_),
    .C1(_10188_),
    .X(_00080_));
 sky130_fd_sc_hd__nand2_2 _13887_ (.A(_10136_),
    .B(_10152_),
    .Y(_10191_));
 sky130_fd_sc_hd__o211a_2 _13888_ (.A1(\decode.regfile.registers_23[29] ),
    .A2(_10180_),
    .B1(_10191_),
    .C1(_10188_),
    .X(_00081_));
 sky130_fd_sc_hd__nand2_2 _13889_ (.A(_10142_),
    .B(_10152_),
    .Y(_10192_));
 sky130_fd_sc_hd__o211a_2 _13890_ (.A1(\decode.regfile.registers_23[30] ),
    .A2(_10154_),
    .B1(_10192_),
    .C1(_10188_),
    .X(_00082_));
 sky130_fd_sc_hd__nand2_2 _13891_ (.A(_10147_),
    .B(_10152_),
    .Y(_10193_));
 sky130_fd_sc_hd__o211a_2 _13892_ (.A1(\decode.regfile.registers_23[31] ),
    .A2(_10154_),
    .B1(_10193_),
    .C1(_10188_),
    .X(_00083_));
 sky130_fd_sc_hd__buf_1 _13893_ (.A(\decode.io_wb_rd[3] ),
    .X(_10194_));
 sky130_fd_sc_hd__buf_1 _13894_ (.A(_10194_),
    .X(_10195_));
 sky130_fd_sc_hd__nor2_2 _13895_ (.A(\decode.io_wb_rd[0] ),
    .B(\decode.io_wb_rd[1] ),
    .Y(_10196_));
 sky130_fd_sc_hd__and4b_2 _13896_ (.A_N(_09930_),
    .B(_10195_),
    .C(_10149_),
    .D(_10196_),
    .X(_10197_));
 sky130_fd_sc_hd__buf_1 _13897_ (.A(_10197_),
    .X(_10198_));
 sky130_fd_sc_hd__buf_1 _13898_ (.A(_10198_),
    .X(_10199_));
 sky130_fd_sc_hd__buf_1 _13899_ (.A(_10198_),
    .X(_10200_));
 sky130_fd_sc_hd__nand2_2 _13900_ (.A(_09950_),
    .B(_10200_),
    .Y(_10201_));
 sky130_fd_sc_hd__o211a_2 _13901_ (.A1(\decode.regfile.registers_24[0] ),
    .A2(_10199_),
    .B1(_10201_),
    .C1(_10188_),
    .X(_00084_));
 sky130_fd_sc_hd__nand2_2 _13902_ (.A(_09964_),
    .B(_10200_),
    .Y(_10202_));
 sky130_fd_sc_hd__o211a_2 _13903_ (.A1(\decode.regfile.registers_24[1] ),
    .A2(_10199_),
    .B1(_10202_),
    .C1(_10188_),
    .X(_00085_));
 sky130_fd_sc_hd__nand2_2 _13904_ (.A(_09970_),
    .B(_10200_),
    .Y(_10203_));
 sky130_fd_sc_hd__o211a_2 _13905_ (.A1(\decode.regfile.registers_24[2] ),
    .A2(_10199_),
    .B1(_10203_),
    .C1(_10188_),
    .X(_00086_));
 sky130_fd_sc_hd__nand2_2 _13906_ (.A(_09975_),
    .B(_10200_),
    .Y(_10204_));
 sky130_fd_sc_hd__o211a_2 _13907_ (.A1(\decode.regfile.registers_24[3] ),
    .A2(_10199_),
    .B1(_10204_),
    .C1(_10188_),
    .X(_00087_));
 sky130_fd_sc_hd__nand2_2 _13908_ (.A(_09984_),
    .B(_10200_),
    .Y(_10205_));
 sky130_fd_sc_hd__buf_1 _13909_ (.A(_10131_),
    .X(_10206_));
 sky130_fd_sc_hd__o211a_2 _13910_ (.A1(\decode.regfile.registers_24[4] ),
    .A2(_10199_),
    .B1(_10205_),
    .C1(_10206_),
    .X(_00088_));
 sky130_fd_sc_hd__nand2_2 _13911_ (.A(_09993_),
    .B(_10200_),
    .Y(_10207_));
 sky130_fd_sc_hd__o211a_2 _13912_ (.A1(\decode.regfile.registers_24[5] ),
    .A2(_10199_),
    .B1(_10207_),
    .C1(_10206_),
    .X(_00089_));
 sky130_fd_sc_hd__nand2_2 _13913_ (.A(_09999_),
    .B(_10200_),
    .Y(_10208_));
 sky130_fd_sc_hd__o211a_2 _13914_ (.A1(\decode.regfile.registers_24[6] ),
    .A2(_10199_),
    .B1(_10208_),
    .C1(_10206_),
    .X(_00090_));
 sky130_fd_sc_hd__nand2_2 _13915_ (.A(_10008_),
    .B(_10200_),
    .Y(_10209_));
 sky130_fd_sc_hd__o211a_2 _13916_ (.A1(\decode.regfile.registers_24[7] ),
    .A2(_10199_),
    .B1(_10209_),
    .C1(_10206_),
    .X(_00091_));
 sky130_fd_sc_hd__buf_1 _13917_ (.A(_10198_),
    .X(_10210_));
 sky130_fd_sc_hd__nand2_2 _13918_ (.A(_10015_),
    .B(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__o211a_2 _13919_ (.A1(\decode.regfile.registers_24[8] ),
    .A2(_10199_),
    .B1(_10211_),
    .C1(_10206_),
    .X(_00092_));
 sky130_fd_sc_hd__nand2_2 _13920_ (.A(_10025_),
    .B(_10210_),
    .Y(_10212_));
 sky130_fd_sc_hd__o211a_2 _13921_ (.A1(\decode.regfile.registers_24[9] ),
    .A2(_10199_),
    .B1(_10212_),
    .C1(_10206_),
    .X(_00093_));
 sky130_fd_sc_hd__buf_1 _13922_ (.A(_10198_),
    .X(_10213_));
 sky130_fd_sc_hd__nand2_2 _13923_ (.A(_10031_),
    .B(_10210_),
    .Y(_10214_));
 sky130_fd_sc_hd__o211a_2 _13924_ (.A1(\decode.regfile.registers_24[10] ),
    .A2(_10213_),
    .B1(_10214_),
    .C1(_10206_),
    .X(_00094_));
 sky130_fd_sc_hd__nand2_2 _13925_ (.A(_10036_),
    .B(_10210_),
    .Y(_10215_));
 sky130_fd_sc_hd__o211a_2 _13926_ (.A1(\decode.regfile.registers_24[11] ),
    .A2(_10213_),
    .B1(_10215_),
    .C1(_10206_),
    .X(_00095_));
 sky130_fd_sc_hd__nand2_2 _13927_ (.A(_10042_),
    .B(_10210_),
    .Y(_10216_));
 sky130_fd_sc_hd__o211a_2 _13928_ (.A1(\decode.regfile.registers_24[12] ),
    .A2(_10213_),
    .B1(_10216_),
    .C1(_10206_),
    .X(_00096_));
 sky130_fd_sc_hd__nand2_2 _13929_ (.A(_10048_),
    .B(_10210_),
    .Y(_10217_));
 sky130_fd_sc_hd__o211a_2 _13930_ (.A1(\decode.regfile.registers_24[13] ),
    .A2(_10213_),
    .B1(_10217_),
    .C1(_10206_),
    .X(_00097_));
 sky130_fd_sc_hd__nand2_2 _13931_ (.A(_10053_),
    .B(_10210_),
    .Y(_10218_));
 sky130_fd_sc_hd__buf_1 _13932_ (.A(_10131_),
    .X(_10219_));
 sky130_fd_sc_hd__o211a_2 _13933_ (.A1(\decode.regfile.registers_24[14] ),
    .A2(_10213_),
    .B1(_10218_),
    .C1(_10219_),
    .X(_00098_));
 sky130_fd_sc_hd__nand2_2 _13934_ (.A(_10058_),
    .B(_10210_),
    .Y(_10220_));
 sky130_fd_sc_hd__o211a_2 _13935_ (.A1(\decode.regfile.registers_24[15] ),
    .A2(_10213_),
    .B1(_10220_),
    .C1(_10219_),
    .X(_00099_));
 sky130_fd_sc_hd__nand2_2 _13936_ (.A(_10064_),
    .B(_10210_),
    .Y(_10221_));
 sky130_fd_sc_hd__o211a_2 _13937_ (.A1(\decode.regfile.registers_24[16] ),
    .A2(_10213_),
    .B1(_10221_),
    .C1(_10219_),
    .X(_00100_));
 sky130_fd_sc_hd__nand2_2 _13938_ (.A(_10069_),
    .B(_10210_),
    .Y(_10222_));
 sky130_fd_sc_hd__o211a_2 _13939_ (.A1(\decode.regfile.registers_24[17] ),
    .A2(_10213_),
    .B1(_10222_),
    .C1(_10219_),
    .X(_00101_));
 sky130_fd_sc_hd__buf_1 _13940_ (.A(_10198_),
    .X(_10223_));
 sky130_fd_sc_hd__nand2_2 _13941_ (.A(_10074_),
    .B(_10223_),
    .Y(_10224_));
 sky130_fd_sc_hd__o211a_2 _13942_ (.A1(\decode.regfile.registers_24[18] ),
    .A2(_10213_),
    .B1(_10224_),
    .C1(_10219_),
    .X(_00102_));
 sky130_fd_sc_hd__nand2_2 _13943_ (.A(_10081_),
    .B(_10223_),
    .Y(_10225_));
 sky130_fd_sc_hd__o211a_2 _13944_ (.A1(\decode.regfile.registers_24[19] ),
    .A2(_10213_),
    .B1(_10225_),
    .C1(_10219_),
    .X(_00103_));
 sky130_fd_sc_hd__buf_1 _13945_ (.A(_10198_),
    .X(_10226_));
 sky130_fd_sc_hd__nand2_2 _13946_ (.A(_10087_),
    .B(_10223_),
    .Y(_10227_));
 sky130_fd_sc_hd__o211a_2 _13947_ (.A1(\decode.regfile.registers_24[20] ),
    .A2(_10226_),
    .B1(_10227_),
    .C1(_10219_),
    .X(_00104_));
 sky130_fd_sc_hd__nand2_2 _13948_ (.A(_10092_),
    .B(_10223_),
    .Y(_10228_));
 sky130_fd_sc_hd__o211a_2 _13949_ (.A1(\decode.regfile.registers_24[21] ),
    .A2(_10226_),
    .B1(_10228_),
    .C1(_10219_),
    .X(_00105_));
 sky130_fd_sc_hd__nand2_2 _13950_ (.A(_10097_),
    .B(_10223_),
    .Y(_10229_));
 sky130_fd_sc_hd__o211a_2 _13951_ (.A1(\decode.regfile.registers_24[22] ),
    .A2(_10226_),
    .B1(_10229_),
    .C1(_10219_),
    .X(_00106_));
 sky130_fd_sc_hd__nand2_2 _13952_ (.A(_10102_),
    .B(_10223_),
    .Y(_10230_));
 sky130_fd_sc_hd__o211a_2 _13953_ (.A1(\decode.regfile.registers_24[23] ),
    .A2(_10226_),
    .B1(_10230_),
    .C1(_10219_),
    .X(_00107_));
 sky130_fd_sc_hd__nand2_2 _13954_ (.A(_10107_),
    .B(_10223_),
    .Y(_10231_));
 sky130_fd_sc_hd__buf_1 _13955_ (.A(_10131_),
    .X(_10232_));
 sky130_fd_sc_hd__o211a_2 _13956_ (.A1(\decode.regfile.registers_24[24] ),
    .A2(_10226_),
    .B1(_10231_),
    .C1(_10232_),
    .X(_00108_));
 sky130_fd_sc_hd__nand2_2 _13957_ (.A(_10112_),
    .B(_10223_),
    .Y(_10233_));
 sky130_fd_sc_hd__o211a_2 _13958_ (.A1(\decode.regfile.registers_24[25] ),
    .A2(_10226_),
    .B1(_10233_),
    .C1(_10232_),
    .X(_00109_));
 sky130_fd_sc_hd__nand2_2 _13959_ (.A(_10117_),
    .B(_10223_),
    .Y(_10234_));
 sky130_fd_sc_hd__o211a_2 _13960_ (.A1(\decode.regfile.registers_24[26] ),
    .A2(_10226_),
    .B1(_10234_),
    .C1(_10232_),
    .X(_00110_));
 sky130_fd_sc_hd__nand2_2 _13961_ (.A(_10122_),
    .B(_10223_),
    .Y(_10235_));
 sky130_fd_sc_hd__o211a_2 _13962_ (.A1(\decode.regfile.registers_24[27] ),
    .A2(_10226_),
    .B1(_10235_),
    .C1(_10232_),
    .X(_00111_));
 sky130_fd_sc_hd__nand2_2 _13963_ (.A(_10128_),
    .B(_10198_),
    .Y(_10236_));
 sky130_fd_sc_hd__o211a_2 _13964_ (.A1(\decode.regfile.registers_24[28] ),
    .A2(_10226_),
    .B1(_10236_),
    .C1(_10232_),
    .X(_00112_));
 sky130_fd_sc_hd__nand2_2 _13965_ (.A(_10136_),
    .B(_10198_),
    .Y(_10237_));
 sky130_fd_sc_hd__o211a_2 _13966_ (.A1(\decode.regfile.registers_24[29] ),
    .A2(_10226_),
    .B1(_10237_),
    .C1(_10232_),
    .X(_00113_));
 sky130_fd_sc_hd__nand2_2 _13967_ (.A(_10142_),
    .B(_10198_),
    .Y(_10238_));
 sky130_fd_sc_hd__o211a_2 _13968_ (.A1(\decode.regfile.registers_24[30] ),
    .A2(_10200_),
    .B1(_10238_),
    .C1(_10232_),
    .X(_00114_));
 sky130_fd_sc_hd__nand2_2 _13969_ (.A(_10147_),
    .B(_10198_),
    .Y(_10239_));
 sky130_fd_sc_hd__o211a_2 _13970_ (.A1(\decode.regfile.registers_24[31] ),
    .A2(_10200_),
    .B1(_10239_),
    .C1(_10232_),
    .X(_00115_));
 sky130_fd_sc_hd__and2_2 _13971_ (.A(_09931_),
    .B(\decode.io_wb_rd[0] ),
    .X(_10240_));
 sky130_fd_sc_hd__and4b_2 _13972_ (.A_N(_09930_),
    .B(_10194_),
    .C(_09933_),
    .D(_10240_),
    .X(_10241_));
 sky130_fd_sc_hd__buf_1 _13973_ (.A(_10241_),
    .X(_10242_));
 sky130_fd_sc_hd__buf_1 _13974_ (.A(_10242_),
    .X(_10243_));
 sky130_fd_sc_hd__buf_1 _13975_ (.A(_10242_),
    .X(_10244_));
 sky130_fd_sc_hd__buf_1 _13976_ (.A(_09949_),
    .X(_10245_));
 sky130_fd_sc_hd__nand2_2 _13977_ (.A(_10244_),
    .B(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__o211a_2 _13978_ (.A1(\decode.regfile.registers_25[0] ),
    .A2(_10243_),
    .B1(_10246_),
    .C1(_10232_),
    .X(_00116_));
 sky130_fd_sc_hd__nand2_2 _13979_ (.A(_10244_),
    .B(_09963_),
    .Y(_10247_));
 sky130_fd_sc_hd__o211a_2 _13980_ (.A1(\decode.regfile.registers_25[1] ),
    .A2(_10243_),
    .B1(_10247_),
    .C1(_10232_),
    .X(_00117_));
 sky130_fd_sc_hd__nand2_2 _13981_ (.A(_09970_),
    .B(_10244_),
    .Y(_10248_));
 sky130_fd_sc_hd__buf_1 _13982_ (.A(_10131_),
    .X(_10249_));
 sky130_fd_sc_hd__o211a_2 _13983_ (.A1(\decode.regfile.registers_25[2] ),
    .A2(_10243_),
    .B1(_10248_),
    .C1(_10249_),
    .X(_00118_));
 sky130_fd_sc_hd__nand2_2 _13984_ (.A(_09975_),
    .B(_10244_),
    .Y(_10250_));
 sky130_fd_sc_hd__o211a_2 _13985_ (.A1(\decode.regfile.registers_25[3] ),
    .A2(_10243_),
    .B1(_10250_),
    .C1(_10249_),
    .X(_00119_));
 sky130_fd_sc_hd__nand2_2 _13986_ (.A(_09984_),
    .B(_10244_),
    .Y(_10251_));
 sky130_fd_sc_hd__o211a_2 _13987_ (.A1(\decode.regfile.registers_25[4] ),
    .A2(_10243_),
    .B1(_10251_),
    .C1(_10249_),
    .X(_00120_));
 sky130_fd_sc_hd__nand2_2 _13988_ (.A(_09993_),
    .B(_10244_),
    .Y(_10252_));
 sky130_fd_sc_hd__o211a_2 _13989_ (.A1(\decode.regfile.registers_25[5] ),
    .A2(_10243_),
    .B1(_10252_),
    .C1(_10249_),
    .X(_00121_));
 sky130_fd_sc_hd__nand2_2 _13990_ (.A(_09999_),
    .B(_10244_),
    .Y(_10253_));
 sky130_fd_sc_hd__o211a_2 _13991_ (.A1(\decode.regfile.registers_25[6] ),
    .A2(_10243_),
    .B1(_10253_),
    .C1(_10249_),
    .X(_00122_));
 sky130_fd_sc_hd__nand2_2 _13992_ (.A(_10008_),
    .B(_10244_),
    .Y(_10254_));
 sky130_fd_sc_hd__o211a_2 _13993_ (.A1(\decode.regfile.registers_25[7] ),
    .A2(_10243_),
    .B1(_10254_),
    .C1(_10249_),
    .X(_00123_));
 sky130_fd_sc_hd__buf_1 _13994_ (.A(_10242_),
    .X(_10255_));
 sky130_fd_sc_hd__nand2_2 _13995_ (.A(_10015_),
    .B(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__o211a_2 _13996_ (.A1(\decode.regfile.registers_25[8] ),
    .A2(_10243_),
    .B1(_10256_),
    .C1(_10249_),
    .X(_00124_));
 sky130_fd_sc_hd__nand2_2 _13997_ (.A(_10025_),
    .B(_10255_),
    .Y(_10257_));
 sky130_fd_sc_hd__o211a_2 _13998_ (.A1(\decode.regfile.registers_25[9] ),
    .A2(_10243_),
    .B1(_10257_),
    .C1(_10249_),
    .X(_00125_));
 sky130_fd_sc_hd__buf_1 _13999_ (.A(_10242_),
    .X(_10258_));
 sky130_fd_sc_hd__nand2_2 _14000_ (.A(_10031_),
    .B(_10255_),
    .Y(_10259_));
 sky130_fd_sc_hd__o211a_2 _14001_ (.A1(\decode.regfile.registers_25[10] ),
    .A2(_10258_),
    .B1(_10259_),
    .C1(_10249_),
    .X(_00126_));
 sky130_fd_sc_hd__nand2_2 _14002_ (.A(_10036_),
    .B(_10255_),
    .Y(_10260_));
 sky130_fd_sc_hd__o211a_2 _14003_ (.A1(\decode.regfile.registers_25[11] ),
    .A2(_10258_),
    .B1(_10260_),
    .C1(_10249_),
    .X(_00127_));
 sky130_fd_sc_hd__nand2_2 _14004_ (.A(_10042_),
    .B(_10255_),
    .Y(_10261_));
 sky130_fd_sc_hd__buf_1 _14005_ (.A(_10131_),
    .X(_10262_));
 sky130_fd_sc_hd__o211a_2 _14006_ (.A1(\decode.regfile.registers_25[12] ),
    .A2(_10258_),
    .B1(_10261_),
    .C1(_10262_),
    .X(_00128_));
 sky130_fd_sc_hd__nand2_2 _14007_ (.A(_10048_),
    .B(_10255_),
    .Y(_10263_));
 sky130_fd_sc_hd__o211a_2 _14008_ (.A1(\decode.regfile.registers_25[13] ),
    .A2(_10258_),
    .B1(_10263_),
    .C1(_10262_),
    .X(_00129_));
 sky130_fd_sc_hd__nand2_2 _14009_ (.A(_10053_),
    .B(_10255_),
    .Y(_10264_));
 sky130_fd_sc_hd__o211a_2 _14010_ (.A1(\decode.regfile.registers_25[14] ),
    .A2(_10258_),
    .B1(_10264_),
    .C1(_10262_),
    .X(_00130_));
 sky130_fd_sc_hd__nand2_2 _14011_ (.A(_10058_),
    .B(_10255_),
    .Y(_10265_));
 sky130_fd_sc_hd__o211a_2 _14012_ (.A1(\decode.regfile.registers_25[15] ),
    .A2(_10258_),
    .B1(_10265_),
    .C1(_10262_),
    .X(_00131_));
 sky130_fd_sc_hd__nand2_2 _14013_ (.A(_10064_),
    .B(_10255_),
    .Y(_10266_));
 sky130_fd_sc_hd__o211a_2 _14014_ (.A1(\decode.regfile.registers_25[16] ),
    .A2(_10258_),
    .B1(_10266_),
    .C1(_10262_),
    .X(_00132_));
 sky130_fd_sc_hd__nand2_2 _14015_ (.A(_10069_),
    .B(_10255_),
    .Y(_10267_));
 sky130_fd_sc_hd__o211a_2 _14016_ (.A1(\decode.regfile.registers_25[17] ),
    .A2(_10258_),
    .B1(_10267_),
    .C1(_10262_),
    .X(_00133_));
 sky130_fd_sc_hd__buf_1 _14017_ (.A(_10242_),
    .X(_10268_));
 sky130_fd_sc_hd__nand2_2 _14018_ (.A(_10074_),
    .B(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__o211a_2 _14019_ (.A1(\decode.regfile.registers_25[18] ),
    .A2(_10258_),
    .B1(_10269_),
    .C1(_10262_),
    .X(_00134_));
 sky130_fd_sc_hd__nand2_2 _14020_ (.A(_10081_),
    .B(_10268_),
    .Y(_10270_));
 sky130_fd_sc_hd__o211a_2 _14021_ (.A1(\decode.regfile.registers_25[19] ),
    .A2(_10258_),
    .B1(_10270_),
    .C1(_10262_),
    .X(_00135_));
 sky130_fd_sc_hd__buf_1 _14022_ (.A(_10242_),
    .X(_10271_));
 sky130_fd_sc_hd__nand2_2 _14023_ (.A(_10087_),
    .B(_10268_),
    .Y(_10272_));
 sky130_fd_sc_hd__o211a_2 _14024_ (.A1(\decode.regfile.registers_25[20] ),
    .A2(_10271_),
    .B1(_10272_),
    .C1(_10262_),
    .X(_00136_));
 sky130_fd_sc_hd__nand2_2 _14025_ (.A(_10092_),
    .B(_10268_),
    .Y(_10273_));
 sky130_fd_sc_hd__o211a_2 _14026_ (.A1(\decode.regfile.registers_25[21] ),
    .A2(_10271_),
    .B1(_10273_),
    .C1(_10262_),
    .X(_00137_));
 sky130_fd_sc_hd__nand2_2 _14027_ (.A(_10097_),
    .B(_10268_),
    .Y(_10274_));
 sky130_fd_sc_hd__buf_1 _14028_ (.A(_10131_),
    .X(_10275_));
 sky130_fd_sc_hd__o211a_2 _14029_ (.A1(\decode.regfile.registers_25[22] ),
    .A2(_10271_),
    .B1(_10274_),
    .C1(_10275_),
    .X(_00138_));
 sky130_fd_sc_hd__nand2_2 _14030_ (.A(_10102_),
    .B(_10268_),
    .Y(_10276_));
 sky130_fd_sc_hd__o211a_2 _14031_ (.A1(\decode.regfile.registers_25[23] ),
    .A2(_10271_),
    .B1(_10276_),
    .C1(_10275_),
    .X(_00139_));
 sky130_fd_sc_hd__nand2_2 _14032_ (.A(_10107_),
    .B(_10268_),
    .Y(_10277_));
 sky130_fd_sc_hd__o211a_2 _14033_ (.A1(\decode.regfile.registers_25[24] ),
    .A2(_10271_),
    .B1(_10277_),
    .C1(_10275_),
    .X(_00140_));
 sky130_fd_sc_hd__nand2_2 _14034_ (.A(_10112_),
    .B(_10268_),
    .Y(_10278_));
 sky130_fd_sc_hd__o211a_2 _14035_ (.A1(\decode.regfile.registers_25[25] ),
    .A2(_10271_),
    .B1(_10278_),
    .C1(_10275_),
    .X(_00141_));
 sky130_fd_sc_hd__nand2_2 _14036_ (.A(_10117_),
    .B(_10268_),
    .Y(_10279_));
 sky130_fd_sc_hd__o211a_2 _14037_ (.A1(\decode.regfile.registers_25[26] ),
    .A2(_10271_),
    .B1(_10279_),
    .C1(_10275_),
    .X(_00142_));
 sky130_fd_sc_hd__nand2_2 _14038_ (.A(_10122_),
    .B(_10268_),
    .Y(_10280_));
 sky130_fd_sc_hd__o211a_2 _14039_ (.A1(\decode.regfile.registers_25[27] ),
    .A2(_10271_),
    .B1(_10280_),
    .C1(_10275_),
    .X(_00143_));
 sky130_fd_sc_hd__nand2_2 _14040_ (.A(_10128_),
    .B(_10242_),
    .Y(_10281_));
 sky130_fd_sc_hd__o211a_2 _14041_ (.A1(\decode.regfile.registers_25[28] ),
    .A2(_10271_),
    .B1(_10281_),
    .C1(_10275_),
    .X(_00144_));
 sky130_fd_sc_hd__nand2_2 _14042_ (.A(_10136_),
    .B(_10242_),
    .Y(_10282_));
 sky130_fd_sc_hd__o211a_2 _14043_ (.A1(\decode.regfile.registers_25[29] ),
    .A2(_10271_),
    .B1(_10282_),
    .C1(_10275_),
    .X(_00145_));
 sky130_fd_sc_hd__nand2_2 _14044_ (.A(_10142_),
    .B(_10242_),
    .Y(_10283_));
 sky130_fd_sc_hd__o211a_2 _14045_ (.A1(\decode.regfile.registers_25[30] ),
    .A2(_10244_),
    .B1(_10283_),
    .C1(_10275_),
    .X(_00146_));
 sky130_fd_sc_hd__nand2_2 _14046_ (.A(_10147_),
    .B(_10242_),
    .Y(_10284_));
 sky130_fd_sc_hd__o211a_2 _14047_ (.A1(\decode.regfile.registers_25[31] ),
    .A2(_10244_),
    .B1(_10284_),
    .C1(_10275_),
    .X(_00147_));
 sky130_fd_sc_hd__and4b_2 _14048_ (.A_N(_09930_),
    .B(_10195_),
    .C(_09932_),
    .D(_09933_),
    .X(_10285_));
 sky130_fd_sc_hd__buf_1 _14049_ (.A(_10285_),
    .X(_10286_));
 sky130_fd_sc_hd__buf_1 _14050_ (.A(_10286_),
    .X(_10287_));
 sky130_fd_sc_hd__buf_1 _14051_ (.A(_10286_),
    .X(_10288_));
 sky130_fd_sc_hd__nand2_2 _14052_ (.A(_09950_),
    .B(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__buf_1 _14053_ (.A(_10130_),
    .X(_10290_));
 sky130_fd_sc_hd__buf_1 _14054_ (.A(_10290_),
    .X(_10291_));
 sky130_fd_sc_hd__o211a_2 _14055_ (.A1(\decode.regfile.registers_26[0] ),
    .A2(_10287_),
    .B1(_10289_),
    .C1(_10291_),
    .X(_00148_));
 sky130_fd_sc_hd__nand2_2 _14056_ (.A(_09964_),
    .B(_10288_),
    .Y(_10292_));
 sky130_fd_sc_hd__o211a_2 _14057_ (.A1(\decode.regfile.registers_26[1] ),
    .A2(_10287_),
    .B1(_10292_),
    .C1(_10291_),
    .X(_00149_));
 sky130_fd_sc_hd__nand2_2 _14058_ (.A(_09970_),
    .B(_10288_),
    .Y(_10293_));
 sky130_fd_sc_hd__o211a_2 _14059_ (.A1(\decode.regfile.registers_26[2] ),
    .A2(_10287_),
    .B1(_10293_),
    .C1(_10291_),
    .X(_00150_));
 sky130_fd_sc_hd__nand2_2 _14060_ (.A(_09975_),
    .B(_10288_),
    .Y(_10294_));
 sky130_fd_sc_hd__o211a_2 _14061_ (.A1(\decode.regfile.registers_26[3] ),
    .A2(_10287_),
    .B1(_10294_),
    .C1(_10291_),
    .X(_00151_));
 sky130_fd_sc_hd__nand2_2 _14062_ (.A(_09984_),
    .B(_10288_),
    .Y(_10295_));
 sky130_fd_sc_hd__o211a_2 _14063_ (.A1(\decode.regfile.registers_26[4] ),
    .A2(_10287_),
    .B1(_10295_),
    .C1(_10291_),
    .X(_00152_));
 sky130_fd_sc_hd__nand2_2 _14064_ (.A(_09993_),
    .B(_10288_),
    .Y(_10296_));
 sky130_fd_sc_hd__o211a_2 _14065_ (.A1(\decode.regfile.registers_26[5] ),
    .A2(_10287_),
    .B1(_10296_),
    .C1(_10291_),
    .X(_00153_));
 sky130_fd_sc_hd__nand2_2 _14066_ (.A(_09999_),
    .B(_10288_),
    .Y(_10297_));
 sky130_fd_sc_hd__o211a_2 _14067_ (.A1(\decode.regfile.registers_26[6] ),
    .A2(_10287_),
    .B1(_10297_),
    .C1(_10291_),
    .X(_00154_));
 sky130_fd_sc_hd__nand2_2 _14068_ (.A(_10008_),
    .B(_10288_),
    .Y(_10298_));
 sky130_fd_sc_hd__o211a_2 _14069_ (.A1(\decode.regfile.registers_26[7] ),
    .A2(_10287_),
    .B1(_10298_),
    .C1(_10291_),
    .X(_00155_));
 sky130_fd_sc_hd__buf_1 _14070_ (.A(_10286_),
    .X(_10299_));
 sky130_fd_sc_hd__nand2_2 _14071_ (.A(_10015_),
    .B(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__o211a_2 _14072_ (.A1(\decode.regfile.registers_26[8] ),
    .A2(_10287_),
    .B1(_10300_),
    .C1(_10291_),
    .X(_00156_));
 sky130_fd_sc_hd__nand2_2 _14073_ (.A(_10025_),
    .B(_10299_),
    .Y(_10301_));
 sky130_fd_sc_hd__o211a_2 _14074_ (.A1(\decode.regfile.registers_26[9] ),
    .A2(_10287_),
    .B1(_10301_),
    .C1(_10291_),
    .X(_00157_));
 sky130_fd_sc_hd__buf_1 _14075_ (.A(_10286_),
    .X(_10302_));
 sky130_fd_sc_hd__nand2_2 _14076_ (.A(_10031_),
    .B(_10299_),
    .Y(_10303_));
 sky130_fd_sc_hd__buf_1 _14077_ (.A(_10290_),
    .X(_10304_));
 sky130_fd_sc_hd__o211a_2 _14078_ (.A1(\decode.regfile.registers_26[10] ),
    .A2(_10302_),
    .B1(_10303_),
    .C1(_10304_),
    .X(_00158_));
 sky130_fd_sc_hd__nand2_2 _14079_ (.A(_10036_),
    .B(_10299_),
    .Y(_10305_));
 sky130_fd_sc_hd__o211a_2 _14080_ (.A1(\decode.regfile.registers_26[11] ),
    .A2(_10302_),
    .B1(_10305_),
    .C1(_10304_),
    .X(_00159_));
 sky130_fd_sc_hd__nand2_2 _14081_ (.A(_10042_),
    .B(_10299_),
    .Y(_10306_));
 sky130_fd_sc_hd__o211a_2 _14082_ (.A1(\decode.regfile.registers_26[12] ),
    .A2(_10302_),
    .B1(_10306_),
    .C1(_10304_),
    .X(_00160_));
 sky130_fd_sc_hd__nand2_2 _14083_ (.A(_10048_),
    .B(_10299_),
    .Y(_10307_));
 sky130_fd_sc_hd__o211a_2 _14084_ (.A1(\decode.regfile.registers_26[13] ),
    .A2(_10302_),
    .B1(_10307_),
    .C1(_10304_),
    .X(_00161_));
 sky130_fd_sc_hd__nand2_2 _14085_ (.A(_10053_),
    .B(_10299_),
    .Y(_10308_));
 sky130_fd_sc_hd__o211a_2 _14086_ (.A1(\decode.regfile.registers_26[14] ),
    .A2(_10302_),
    .B1(_10308_),
    .C1(_10304_),
    .X(_00162_));
 sky130_fd_sc_hd__nand2_2 _14087_ (.A(_10058_),
    .B(_10299_),
    .Y(_10309_));
 sky130_fd_sc_hd__o211a_2 _14088_ (.A1(\decode.regfile.registers_26[15] ),
    .A2(_10302_),
    .B1(_10309_),
    .C1(_10304_),
    .X(_00163_));
 sky130_fd_sc_hd__nand2_2 _14089_ (.A(_10064_),
    .B(_10299_),
    .Y(_10310_));
 sky130_fd_sc_hd__o211a_2 _14090_ (.A1(\decode.regfile.registers_26[16] ),
    .A2(_10302_),
    .B1(_10310_),
    .C1(_10304_),
    .X(_00164_));
 sky130_fd_sc_hd__nand2_2 _14091_ (.A(_10069_),
    .B(_10299_),
    .Y(_10311_));
 sky130_fd_sc_hd__o211a_2 _14092_ (.A1(\decode.regfile.registers_26[17] ),
    .A2(_10302_),
    .B1(_10311_),
    .C1(_10304_),
    .X(_00165_));
 sky130_fd_sc_hd__buf_1 _14093_ (.A(_10286_),
    .X(_10312_));
 sky130_fd_sc_hd__nand2_2 _14094_ (.A(_10074_),
    .B(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__o211a_2 _14095_ (.A1(\decode.regfile.registers_26[18] ),
    .A2(_10302_),
    .B1(_10313_),
    .C1(_10304_),
    .X(_00166_));
 sky130_fd_sc_hd__nand2_2 _14096_ (.A(_10081_),
    .B(_10312_),
    .Y(_10314_));
 sky130_fd_sc_hd__o211a_2 _14097_ (.A1(\decode.regfile.registers_26[19] ),
    .A2(_10302_),
    .B1(_10314_),
    .C1(_10304_),
    .X(_00167_));
 sky130_fd_sc_hd__buf_1 _14098_ (.A(_10286_),
    .X(_10315_));
 sky130_fd_sc_hd__nand2_2 _14099_ (.A(_10087_),
    .B(_10312_),
    .Y(_10316_));
 sky130_fd_sc_hd__buf_1 _14100_ (.A(_10290_),
    .X(_10317_));
 sky130_fd_sc_hd__o211a_2 _14101_ (.A1(\decode.regfile.registers_26[20] ),
    .A2(_10315_),
    .B1(_10316_),
    .C1(_10317_),
    .X(_00168_));
 sky130_fd_sc_hd__nand2_2 _14102_ (.A(_10092_),
    .B(_10312_),
    .Y(_10318_));
 sky130_fd_sc_hd__o211a_2 _14103_ (.A1(\decode.regfile.registers_26[21] ),
    .A2(_10315_),
    .B1(_10318_),
    .C1(_10317_),
    .X(_00169_));
 sky130_fd_sc_hd__nand2_2 _14104_ (.A(_10097_),
    .B(_10312_),
    .Y(_10319_));
 sky130_fd_sc_hd__o211a_2 _14105_ (.A1(\decode.regfile.registers_26[22] ),
    .A2(_10315_),
    .B1(_10319_),
    .C1(_10317_),
    .X(_00170_));
 sky130_fd_sc_hd__nand2_2 _14106_ (.A(_10102_),
    .B(_10312_),
    .Y(_10320_));
 sky130_fd_sc_hd__o211a_2 _14107_ (.A1(\decode.regfile.registers_26[23] ),
    .A2(_10315_),
    .B1(_10320_),
    .C1(_10317_),
    .X(_00171_));
 sky130_fd_sc_hd__nand2_2 _14108_ (.A(_10107_),
    .B(_10312_),
    .Y(_10321_));
 sky130_fd_sc_hd__o211a_2 _14109_ (.A1(\decode.regfile.registers_26[24] ),
    .A2(_10315_),
    .B1(_10321_),
    .C1(_10317_),
    .X(_00172_));
 sky130_fd_sc_hd__nand2_2 _14110_ (.A(_10112_),
    .B(_10312_),
    .Y(_10322_));
 sky130_fd_sc_hd__o211a_2 _14111_ (.A1(\decode.regfile.registers_26[25] ),
    .A2(_10315_),
    .B1(_10322_),
    .C1(_10317_),
    .X(_00173_));
 sky130_fd_sc_hd__nand2_2 _14112_ (.A(_10117_),
    .B(_10312_),
    .Y(_10323_));
 sky130_fd_sc_hd__o211a_2 _14113_ (.A1(\decode.regfile.registers_26[26] ),
    .A2(_10315_),
    .B1(_10323_),
    .C1(_10317_),
    .X(_00174_));
 sky130_fd_sc_hd__nand2_2 _14114_ (.A(_10122_),
    .B(_10312_),
    .Y(_10324_));
 sky130_fd_sc_hd__o211a_2 _14115_ (.A1(\decode.regfile.registers_26[27] ),
    .A2(_10315_),
    .B1(_10324_),
    .C1(_10317_),
    .X(_00175_));
 sky130_fd_sc_hd__nand2_2 _14116_ (.A(_10128_),
    .B(_10286_),
    .Y(_10325_));
 sky130_fd_sc_hd__o211a_2 _14117_ (.A1(\decode.regfile.registers_26[28] ),
    .A2(_10315_),
    .B1(_10325_),
    .C1(_10317_),
    .X(_00176_));
 sky130_fd_sc_hd__nand2_2 _14118_ (.A(_10136_),
    .B(_10286_),
    .Y(_10326_));
 sky130_fd_sc_hd__o211a_2 _14119_ (.A1(\decode.regfile.registers_26[29] ),
    .A2(_10315_),
    .B1(_10326_),
    .C1(_10317_),
    .X(_00177_));
 sky130_fd_sc_hd__nand2_2 _14120_ (.A(_10142_),
    .B(_10286_),
    .Y(_10327_));
 sky130_fd_sc_hd__buf_1 _14121_ (.A(_10290_),
    .X(_10328_));
 sky130_fd_sc_hd__o211a_2 _14122_ (.A1(\decode.regfile.registers_26[30] ),
    .A2(_10288_),
    .B1(_10327_),
    .C1(_10328_),
    .X(_00178_));
 sky130_fd_sc_hd__nand2_2 _14123_ (.A(_10147_),
    .B(_10286_),
    .Y(_10329_));
 sky130_fd_sc_hd__o211a_2 _14124_ (.A1(\decode.regfile.registers_26[31] ),
    .A2(_10288_),
    .B1(_10329_),
    .C1(_10328_),
    .X(_00179_));
 sky130_fd_sc_hd__and4b_2 _14125_ (.A_N(_09930_),
    .B(_10194_),
    .C(_10149_),
    .D(_10150_),
    .X(_10330_));
 sky130_fd_sc_hd__buf_1 _14126_ (.A(_10330_),
    .X(_10331_));
 sky130_fd_sc_hd__buf_1 _14127_ (.A(_10331_),
    .X(_10332_));
 sky130_fd_sc_hd__buf_1 _14128_ (.A(_10331_),
    .X(_10333_));
 sky130_fd_sc_hd__nand2_2 _14129_ (.A(_09950_),
    .B(_10333_),
    .Y(_10334_));
 sky130_fd_sc_hd__o211a_2 _14130_ (.A1(\decode.regfile.registers_27[0] ),
    .A2(_10332_),
    .B1(_10334_),
    .C1(_10328_),
    .X(_00180_));
 sky130_fd_sc_hd__nand2_2 _14131_ (.A(_09964_),
    .B(_10333_),
    .Y(_10335_));
 sky130_fd_sc_hd__o211a_2 _14132_ (.A1(\decode.regfile.registers_27[1] ),
    .A2(_10332_),
    .B1(_10335_),
    .C1(_10328_),
    .X(_00181_));
 sky130_fd_sc_hd__nand2_2 _14133_ (.A(_09970_),
    .B(_10333_),
    .Y(_10336_));
 sky130_fd_sc_hd__o211a_2 _14134_ (.A1(\decode.regfile.registers_27[2] ),
    .A2(_10332_),
    .B1(_10336_),
    .C1(_10328_),
    .X(_00182_));
 sky130_fd_sc_hd__nand2_2 _14135_ (.A(_09975_),
    .B(_10333_),
    .Y(_10337_));
 sky130_fd_sc_hd__o211a_2 _14136_ (.A1(\decode.regfile.registers_27[3] ),
    .A2(_10332_),
    .B1(_10337_),
    .C1(_10328_),
    .X(_00183_));
 sky130_fd_sc_hd__nand2_2 _14137_ (.A(_09984_),
    .B(_10333_),
    .Y(_10338_));
 sky130_fd_sc_hd__o211a_2 _14138_ (.A1(\decode.regfile.registers_27[4] ),
    .A2(_10332_),
    .B1(_10338_),
    .C1(_10328_),
    .X(_00184_));
 sky130_fd_sc_hd__nand2_2 _14139_ (.A(_09993_),
    .B(_10333_),
    .Y(_10339_));
 sky130_fd_sc_hd__o211a_2 _14140_ (.A1(\decode.regfile.registers_27[5] ),
    .A2(_10332_),
    .B1(_10339_),
    .C1(_10328_),
    .X(_00185_));
 sky130_fd_sc_hd__nand2_2 _14141_ (.A(_09999_),
    .B(_10333_),
    .Y(_10340_));
 sky130_fd_sc_hd__o211a_2 _14142_ (.A1(\decode.regfile.registers_27[6] ),
    .A2(_10332_),
    .B1(_10340_),
    .C1(_10328_),
    .X(_00186_));
 sky130_fd_sc_hd__nand2_2 _14143_ (.A(_10008_),
    .B(_10333_),
    .Y(_10341_));
 sky130_fd_sc_hd__o211a_2 _14144_ (.A1(\decode.regfile.registers_27[7] ),
    .A2(_10332_),
    .B1(_10341_),
    .C1(_10328_),
    .X(_00187_));
 sky130_fd_sc_hd__buf_1 _14145_ (.A(_10331_),
    .X(_10342_));
 sky130_fd_sc_hd__nand2_2 _14146_ (.A(_10015_),
    .B(_10342_),
    .Y(_10343_));
 sky130_fd_sc_hd__buf_1 _14147_ (.A(_10290_),
    .X(_10344_));
 sky130_fd_sc_hd__o211a_2 _14148_ (.A1(\decode.regfile.registers_27[8] ),
    .A2(_10332_),
    .B1(_10343_),
    .C1(_10344_),
    .X(_00188_));
 sky130_fd_sc_hd__nand2_2 _14149_ (.A(_10025_),
    .B(_10342_),
    .Y(_10345_));
 sky130_fd_sc_hd__o211a_2 _14150_ (.A1(\decode.regfile.registers_27[9] ),
    .A2(_10332_),
    .B1(_10345_),
    .C1(_10344_),
    .X(_00189_));
 sky130_fd_sc_hd__buf_1 _14151_ (.A(_10331_),
    .X(_10346_));
 sky130_fd_sc_hd__nand2_2 _14152_ (.A(_10031_),
    .B(_10342_),
    .Y(_10347_));
 sky130_fd_sc_hd__o211a_2 _14153_ (.A1(\decode.regfile.registers_27[10] ),
    .A2(_10346_),
    .B1(_10347_),
    .C1(_10344_),
    .X(_00190_));
 sky130_fd_sc_hd__nand2_2 _14154_ (.A(_10036_),
    .B(_10342_),
    .Y(_10348_));
 sky130_fd_sc_hd__o211a_2 _14155_ (.A1(\decode.regfile.registers_27[11] ),
    .A2(_10346_),
    .B1(_10348_),
    .C1(_10344_),
    .X(_00191_));
 sky130_fd_sc_hd__nand2_2 _14156_ (.A(_10042_),
    .B(_10342_),
    .Y(_10349_));
 sky130_fd_sc_hd__o211a_2 _14157_ (.A1(\decode.regfile.registers_27[12] ),
    .A2(_10346_),
    .B1(_10349_),
    .C1(_10344_),
    .X(_00192_));
 sky130_fd_sc_hd__nand2_2 _14158_ (.A(_10048_),
    .B(_10342_),
    .Y(_10350_));
 sky130_fd_sc_hd__o211a_2 _14159_ (.A1(\decode.regfile.registers_27[13] ),
    .A2(_10346_),
    .B1(_10350_),
    .C1(_10344_),
    .X(_00193_));
 sky130_fd_sc_hd__nand2_2 _14160_ (.A(_10053_),
    .B(_10342_),
    .Y(_10351_));
 sky130_fd_sc_hd__o211a_2 _14161_ (.A1(\decode.regfile.registers_27[14] ),
    .A2(_10346_),
    .B1(_10351_),
    .C1(_10344_),
    .X(_00194_));
 sky130_fd_sc_hd__nand2_2 _14162_ (.A(_10058_),
    .B(_10342_),
    .Y(_10352_));
 sky130_fd_sc_hd__o211a_2 _14163_ (.A1(\decode.regfile.registers_27[15] ),
    .A2(_10346_),
    .B1(_10352_),
    .C1(_10344_),
    .X(_00195_));
 sky130_fd_sc_hd__nand2_2 _14164_ (.A(_10064_),
    .B(_10342_),
    .Y(_10353_));
 sky130_fd_sc_hd__o211a_2 _14165_ (.A1(\decode.regfile.registers_27[16] ),
    .A2(_10346_),
    .B1(_10353_),
    .C1(_10344_),
    .X(_00196_));
 sky130_fd_sc_hd__nand2_2 _14166_ (.A(_10069_),
    .B(_10342_),
    .Y(_10354_));
 sky130_fd_sc_hd__o211a_2 _14167_ (.A1(\decode.regfile.registers_27[17] ),
    .A2(_10346_),
    .B1(_10354_),
    .C1(_10344_),
    .X(_00197_));
 sky130_fd_sc_hd__buf_1 _14168_ (.A(_10331_),
    .X(_10355_));
 sky130_fd_sc_hd__nand2_2 _14169_ (.A(_10074_),
    .B(_10355_),
    .Y(_10356_));
 sky130_fd_sc_hd__buf_1 _14170_ (.A(_10290_),
    .X(_10357_));
 sky130_fd_sc_hd__o211a_2 _14171_ (.A1(\decode.regfile.registers_27[18] ),
    .A2(_10346_),
    .B1(_10356_),
    .C1(_10357_),
    .X(_00198_));
 sky130_fd_sc_hd__nand2_2 _14172_ (.A(_10081_),
    .B(_10355_),
    .Y(_10358_));
 sky130_fd_sc_hd__o211a_2 _14173_ (.A1(\decode.regfile.registers_27[19] ),
    .A2(_10346_),
    .B1(_10358_),
    .C1(_10357_),
    .X(_00199_));
 sky130_fd_sc_hd__buf_1 _14174_ (.A(_10331_),
    .X(_10359_));
 sky130_fd_sc_hd__nand2_2 _14175_ (.A(_10087_),
    .B(_10355_),
    .Y(_10360_));
 sky130_fd_sc_hd__o211a_2 _14176_ (.A1(\decode.regfile.registers_27[20] ),
    .A2(_10359_),
    .B1(_10360_),
    .C1(_10357_),
    .X(_00200_));
 sky130_fd_sc_hd__nand2_2 _14177_ (.A(_10092_),
    .B(_10355_),
    .Y(_10361_));
 sky130_fd_sc_hd__o211a_2 _14178_ (.A1(\decode.regfile.registers_27[21] ),
    .A2(_10359_),
    .B1(_10361_),
    .C1(_10357_),
    .X(_00201_));
 sky130_fd_sc_hd__nand2_2 _14179_ (.A(_10097_),
    .B(_10355_),
    .Y(_10362_));
 sky130_fd_sc_hd__o211a_2 _14180_ (.A1(\decode.regfile.registers_27[22] ),
    .A2(_10359_),
    .B1(_10362_),
    .C1(_10357_),
    .X(_00202_));
 sky130_fd_sc_hd__nand2_2 _14181_ (.A(_10102_),
    .B(_10355_),
    .Y(_10363_));
 sky130_fd_sc_hd__o211a_2 _14182_ (.A1(\decode.regfile.registers_27[23] ),
    .A2(_10359_),
    .B1(_10363_),
    .C1(_10357_),
    .X(_00203_));
 sky130_fd_sc_hd__nand2_2 _14183_ (.A(_10107_),
    .B(_10355_),
    .Y(_10364_));
 sky130_fd_sc_hd__o211a_2 _14184_ (.A1(\decode.regfile.registers_27[24] ),
    .A2(_10359_),
    .B1(_10364_),
    .C1(_10357_),
    .X(_00204_));
 sky130_fd_sc_hd__nand2_2 _14185_ (.A(_10112_),
    .B(_10355_),
    .Y(_10365_));
 sky130_fd_sc_hd__o211a_2 _14186_ (.A1(\decode.regfile.registers_27[25] ),
    .A2(_10359_),
    .B1(_10365_),
    .C1(_10357_),
    .X(_00205_));
 sky130_fd_sc_hd__nand2_2 _14187_ (.A(_10117_),
    .B(_10355_),
    .Y(_10366_));
 sky130_fd_sc_hd__o211a_2 _14188_ (.A1(\decode.regfile.registers_27[26] ),
    .A2(_10359_),
    .B1(_10366_),
    .C1(_10357_),
    .X(_00206_));
 sky130_fd_sc_hd__nand2_2 _14189_ (.A(_10122_),
    .B(_10355_),
    .Y(_10367_));
 sky130_fd_sc_hd__o211a_2 _14190_ (.A1(\decode.regfile.registers_27[27] ),
    .A2(_10359_),
    .B1(_10367_),
    .C1(_10357_),
    .X(_00207_));
 sky130_fd_sc_hd__nand2_2 _14191_ (.A(_10128_),
    .B(_10331_),
    .Y(_10368_));
 sky130_fd_sc_hd__buf_1 _14192_ (.A(_10290_),
    .X(_10369_));
 sky130_fd_sc_hd__o211a_2 _14193_ (.A1(\decode.regfile.registers_27[28] ),
    .A2(_10359_),
    .B1(_10368_),
    .C1(_10369_),
    .X(_00208_));
 sky130_fd_sc_hd__nand2_2 _14194_ (.A(_10136_),
    .B(_10331_),
    .Y(_10370_));
 sky130_fd_sc_hd__o211a_2 _14195_ (.A1(\decode.regfile.registers_27[29] ),
    .A2(_10359_),
    .B1(_10370_),
    .C1(_10369_),
    .X(_00209_));
 sky130_fd_sc_hd__nand2_2 _14196_ (.A(_10142_),
    .B(_10331_),
    .Y(_10371_));
 sky130_fd_sc_hd__o211a_2 _14197_ (.A1(\decode.regfile.registers_27[30] ),
    .A2(_10333_),
    .B1(_10371_),
    .C1(_10369_),
    .X(_00210_));
 sky130_fd_sc_hd__nand2_2 _14198_ (.A(_10147_),
    .B(_10331_),
    .Y(_10372_));
 sky130_fd_sc_hd__o211a_2 _14199_ (.A1(\decode.regfile.registers_27[31] ),
    .A2(_10333_),
    .B1(_10372_),
    .C1(_10369_),
    .X(_00211_));
 sky130_fd_sc_hd__buf_1 _14200_ (.A(_09929_),
    .X(_10373_));
 sky130_fd_sc_hd__and4_2 _14201_ (.A(_10373_),
    .B(_10195_),
    .C(_09933_),
    .D(_10196_),
    .X(_10374_));
 sky130_fd_sc_hd__buf_1 _14202_ (.A(_10374_),
    .X(_10375_));
 sky130_fd_sc_hd__buf_1 _14203_ (.A(_10375_),
    .X(_10376_));
 sky130_fd_sc_hd__buf_1 _14204_ (.A(_10375_),
    .X(_10377_));
 sky130_fd_sc_hd__nand2_2 _14205_ (.A(_09950_),
    .B(_10377_),
    .Y(_10378_));
 sky130_fd_sc_hd__o211a_2 _14206_ (.A1(\decode.regfile.registers_28[0] ),
    .A2(_10376_),
    .B1(_10378_),
    .C1(_10369_),
    .X(_00212_));
 sky130_fd_sc_hd__nand2_2 _14207_ (.A(_09964_),
    .B(_10377_),
    .Y(_10379_));
 sky130_fd_sc_hd__o211a_2 _14208_ (.A1(\decode.regfile.registers_28[1] ),
    .A2(_10376_),
    .B1(_10379_),
    .C1(_10369_),
    .X(_00213_));
 sky130_fd_sc_hd__nand2_2 _14209_ (.A(_09970_),
    .B(_10377_),
    .Y(_10380_));
 sky130_fd_sc_hd__o211a_2 _14210_ (.A1(\decode.regfile.registers_28[2] ),
    .A2(_10376_),
    .B1(_10380_),
    .C1(_10369_),
    .X(_00214_));
 sky130_fd_sc_hd__nand2_2 _14211_ (.A(_09975_),
    .B(_10377_),
    .Y(_10381_));
 sky130_fd_sc_hd__o211a_2 _14212_ (.A1(\decode.regfile.registers_28[3] ),
    .A2(_10376_),
    .B1(_10381_),
    .C1(_10369_),
    .X(_00215_));
 sky130_fd_sc_hd__nand2_2 _14213_ (.A(_09984_),
    .B(_10377_),
    .Y(_10382_));
 sky130_fd_sc_hd__o211a_2 _14214_ (.A1(\decode.regfile.registers_28[4] ),
    .A2(_10376_),
    .B1(_10382_),
    .C1(_10369_),
    .X(_00216_));
 sky130_fd_sc_hd__nand2_2 _14215_ (.A(_09993_),
    .B(_10377_),
    .Y(_10383_));
 sky130_fd_sc_hd__o211a_2 _14216_ (.A1(\decode.regfile.registers_28[5] ),
    .A2(_10376_),
    .B1(_10383_),
    .C1(_10369_),
    .X(_00217_));
 sky130_fd_sc_hd__nand2_2 _14217_ (.A(_09999_),
    .B(_10377_),
    .Y(_10384_));
 sky130_fd_sc_hd__buf_1 _14218_ (.A(_10290_),
    .X(_10385_));
 sky130_fd_sc_hd__o211a_2 _14219_ (.A1(\decode.regfile.registers_28[6] ),
    .A2(_10376_),
    .B1(_10384_),
    .C1(_10385_),
    .X(_00218_));
 sky130_fd_sc_hd__nand2_2 _14220_ (.A(_10008_),
    .B(_10377_),
    .Y(_10386_));
 sky130_fd_sc_hd__o211a_2 _14221_ (.A1(\decode.regfile.registers_28[7] ),
    .A2(_10376_),
    .B1(_10386_),
    .C1(_10385_),
    .X(_00219_));
 sky130_fd_sc_hd__buf_1 _14222_ (.A(_10375_),
    .X(_10387_));
 sky130_fd_sc_hd__nand2_2 _14223_ (.A(_10015_),
    .B(_10387_),
    .Y(_10388_));
 sky130_fd_sc_hd__o211a_2 _14224_ (.A1(\decode.regfile.registers_28[8] ),
    .A2(_10376_),
    .B1(_10388_),
    .C1(_10385_),
    .X(_00220_));
 sky130_fd_sc_hd__nand2_2 _14225_ (.A(_10025_),
    .B(_10387_),
    .Y(_10389_));
 sky130_fd_sc_hd__o211a_2 _14226_ (.A1(\decode.regfile.registers_28[9] ),
    .A2(_10376_),
    .B1(_10389_),
    .C1(_10385_),
    .X(_00221_));
 sky130_fd_sc_hd__buf_1 _14227_ (.A(_10375_),
    .X(_10390_));
 sky130_fd_sc_hd__nand2_2 _14228_ (.A(_10031_),
    .B(_10387_),
    .Y(_10391_));
 sky130_fd_sc_hd__o211a_2 _14229_ (.A1(\decode.regfile.registers_28[10] ),
    .A2(_10390_),
    .B1(_10391_),
    .C1(_10385_),
    .X(_00222_));
 sky130_fd_sc_hd__nand2_2 _14230_ (.A(_10036_),
    .B(_10387_),
    .Y(_10392_));
 sky130_fd_sc_hd__o211a_2 _14231_ (.A1(\decode.regfile.registers_28[11] ),
    .A2(_10390_),
    .B1(_10392_),
    .C1(_10385_),
    .X(_00223_));
 sky130_fd_sc_hd__nand2_2 _14232_ (.A(_10042_),
    .B(_10387_),
    .Y(_10393_));
 sky130_fd_sc_hd__o211a_2 _14233_ (.A1(\decode.regfile.registers_28[12] ),
    .A2(_10390_),
    .B1(_10393_),
    .C1(_10385_),
    .X(_00224_));
 sky130_fd_sc_hd__nand2_2 _14234_ (.A(_10048_),
    .B(_10387_),
    .Y(_10394_));
 sky130_fd_sc_hd__o211a_2 _14235_ (.A1(\decode.regfile.registers_28[13] ),
    .A2(_10390_),
    .B1(_10394_),
    .C1(_10385_),
    .X(_00225_));
 sky130_fd_sc_hd__nand2_2 _14236_ (.A(_10053_),
    .B(_10387_),
    .Y(_10395_));
 sky130_fd_sc_hd__o211a_2 _14237_ (.A1(\decode.regfile.registers_28[14] ),
    .A2(_10390_),
    .B1(_10395_),
    .C1(_10385_),
    .X(_00226_));
 sky130_fd_sc_hd__nand2_2 _14238_ (.A(_10058_),
    .B(_10387_),
    .Y(_10396_));
 sky130_fd_sc_hd__o211a_2 _14239_ (.A1(\decode.regfile.registers_28[15] ),
    .A2(_10390_),
    .B1(_10396_),
    .C1(_10385_),
    .X(_00227_));
 sky130_fd_sc_hd__nand2_2 _14240_ (.A(_10064_),
    .B(_10387_),
    .Y(_10397_));
 sky130_fd_sc_hd__buf_1 _14241_ (.A(_10290_),
    .X(_10398_));
 sky130_fd_sc_hd__o211a_2 _14242_ (.A1(\decode.regfile.registers_28[16] ),
    .A2(_10390_),
    .B1(_10397_),
    .C1(_10398_),
    .X(_00228_));
 sky130_fd_sc_hd__nand2_2 _14243_ (.A(_10069_),
    .B(_10387_),
    .Y(_10399_));
 sky130_fd_sc_hd__o211a_2 _14244_ (.A1(\decode.regfile.registers_28[17] ),
    .A2(_10390_),
    .B1(_10399_),
    .C1(_10398_),
    .X(_00229_));
 sky130_fd_sc_hd__buf_1 _14245_ (.A(_10375_),
    .X(_10400_));
 sky130_fd_sc_hd__nand2_2 _14246_ (.A(_10074_),
    .B(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__o211a_2 _14247_ (.A1(\decode.regfile.registers_28[18] ),
    .A2(_10390_),
    .B1(_10401_),
    .C1(_10398_),
    .X(_00230_));
 sky130_fd_sc_hd__nand2_2 _14248_ (.A(_10081_),
    .B(_10400_),
    .Y(_10402_));
 sky130_fd_sc_hd__o211a_2 _14249_ (.A1(\decode.regfile.registers_28[19] ),
    .A2(_10390_),
    .B1(_10402_),
    .C1(_10398_),
    .X(_00231_));
 sky130_fd_sc_hd__buf_1 _14250_ (.A(_10375_),
    .X(_10403_));
 sky130_fd_sc_hd__nand2_2 _14251_ (.A(_10087_),
    .B(_10400_),
    .Y(_10404_));
 sky130_fd_sc_hd__o211a_2 _14252_ (.A1(\decode.regfile.registers_28[20] ),
    .A2(_10403_),
    .B1(_10404_),
    .C1(_10398_),
    .X(_00232_));
 sky130_fd_sc_hd__nand2_2 _14253_ (.A(_10092_),
    .B(_10400_),
    .Y(_10405_));
 sky130_fd_sc_hd__o211a_2 _14254_ (.A1(\decode.regfile.registers_28[21] ),
    .A2(_10403_),
    .B1(_10405_),
    .C1(_10398_),
    .X(_00233_));
 sky130_fd_sc_hd__nand2_2 _14255_ (.A(_10097_),
    .B(_10400_),
    .Y(_10406_));
 sky130_fd_sc_hd__o211a_2 _14256_ (.A1(\decode.regfile.registers_28[22] ),
    .A2(_10403_),
    .B1(_10406_),
    .C1(_10398_),
    .X(_00234_));
 sky130_fd_sc_hd__nand2_2 _14257_ (.A(_10102_),
    .B(_10400_),
    .Y(_10407_));
 sky130_fd_sc_hd__o211a_2 _14258_ (.A1(\decode.regfile.registers_28[23] ),
    .A2(_10403_),
    .B1(_10407_),
    .C1(_10398_),
    .X(_00235_));
 sky130_fd_sc_hd__nand2_2 _14259_ (.A(_10107_),
    .B(_10400_),
    .Y(_10408_));
 sky130_fd_sc_hd__o211a_2 _14260_ (.A1(\decode.regfile.registers_28[24] ),
    .A2(_10403_),
    .B1(_10408_),
    .C1(_10398_),
    .X(_00236_));
 sky130_fd_sc_hd__nand2_2 _14261_ (.A(_10112_),
    .B(_10400_),
    .Y(_10409_));
 sky130_fd_sc_hd__o211a_2 _14262_ (.A1(\decode.regfile.registers_28[25] ),
    .A2(_10403_),
    .B1(_10409_),
    .C1(_10398_),
    .X(_00237_));
 sky130_fd_sc_hd__nand2_2 _14263_ (.A(_10117_),
    .B(_10400_),
    .Y(_10410_));
 sky130_fd_sc_hd__buf_1 _14264_ (.A(_10290_),
    .X(_10411_));
 sky130_fd_sc_hd__o211a_2 _14265_ (.A1(\decode.regfile.registers_28[26] ),
    .A2(_10403_),
    .B1(_10410_),
    .C1(_10411_),
    .X(_00238_));
 sky130_fd_sc_hd__nand2_2 _14266_ (.A(_10122_),
    .B(_10400_),
    .Y(_10412_));
 sky130_fd_sc_hd__o211a_2 _14267_ (.A1(\decode.regfile.registers_28[27] ),
    .A2(_10403_),
    .B1(_10412_),
    .C1(_10411_),
    .X(_00239_));
 sky130_fd_sc_hd__nand2_2 _14268_ (.A(_10128_),
    .B(_10375_),
    .Y(_10413_));
 sky130_fd_sc_hd__o211a_2 _14269_ (.A1(\decode.regfile.registers_28[28] ),
    .A2(_10403_),
    .B1(_10413_),
    .C1(_10411_),
    .X(_00240_));
 sky130_fd_sc_hd__nand2_2 _14270_ (.A(_10136_),
    .B(_10375_),
    .Y(_10414_));
 sky130_fd_sc_hd__o211a_2 _14271_ (.A1(\decode.regfile.registers_28[29] ),
    .A2(_10403_),
    .B1(_10414_),
    .C1(_10411_),
    .X(_00241_));
 sky130_fd_sc_hd__nand2_2 _14272_ (.A(_10142_),
    .B(_10375_),
    .Y(_10415_));
 sky130_fd_sc_hd__o211a_2 _14273_ (.A1(\decode.regfile.registers_28[30] ),
    .A2(_10377_),
    .B1(_10415_),
    .C1(_10411_),
    .X(_00242_));
 sky130_fd_sc_hd__nand2_2 _14274_ (.A(_10147_),
    .B(_10375_),
    .Y(_10416_));
 sky130_fd_sc_hd__o211a_2 _14275_ (.A1(\decode.regfile.registers_28[31] ),
    .A2(_10377_),
    .B1(_10416_),
    .C1(_10411_),
    .X(_00243_));
 sky130_fd_sc_hd__and4_2 _14276_ (.A(_09929_),
    .B(_10195_),
    .C(_09933_),
    .D(_10240_),
    .X(_10417_));
 sky130_fd_sc_hd__buf_1 _14277_ (.A(_10417_),
    .X(_10418_));
 sky130_fd_sc_hd__buf_1 _14278_ (.A(_10418_),
    .X(_10419_));
 sky130_fd_sc_hd__buf_1 _14279_ (.A(_10418_),
    .X(_10420_));
 sky130_fd_sc_hd__nand2_2 _14280_ (.A(_10420_),
    .B(_10245_),
    .Y(_10421_));
 sky130_fd_sc_hd__o211a_2 _14281_ (.A1(\decode.regfile.registers_29[0] ),
    .A2(_10419_),
    .B1(_10421_),
    .C1(_10411_),
    .X(_00244_));
 sky130_fd_sc_hd__nand2_2 _14282_ (.A(_09964_),
    .B(_10420_),
    .Y(_10422_));
 sky130_fd_sc_hd__o211a_2 _14283_ (.A1(\decode.regfile.registers_29[1] ),
    .A2(_10419_),
    .B1(_10422_),
    .C1(_10411_),
    .X(_00245_));
 sky130_fd_sc_hd__nand2_2 _14284_ (.A(_09970_),
    .B(_10420_),
    .Y(_10423_));
 sky130_fd_sc_hd__o211a_2 _14285_ (.A1(\decode.regfile.registers_29[2] ),
    .A2(_10419_),
    .B1(_10423_),
    .C1(_10411_),
    .X(_00246_));
 sky130_fd_sc_hd__nand2_2 _14286_ (.A(_09975_),
    .B(_10420_),
    .Y(_10424_));
 sky130_fd_sc_hd__o211a_2 _14287_ (.A1(\decode.regfile.registers_29[3] ),
    .A2(_10419_),
    .B1(_10424_),
    .C1(_10411_),
    .X(_00247_));
 sky130_fd_sc_hd__nand2_2 _14288_ (.A(_09984_),
    .B(_10420_),
    .Y(_10425_));
 sky130_fd_sc_hd__buf_1 _14289_ (.A(_10130_),
    .X(_10426_));
 sky130_fd_sc_hd__buf_1 _14290_ (.A(_10426_),
    .X(_10427_));
 sky130_fd_sc_hd__o211a_2 _14291_ (.A1(\decode.regfile.registers_29[4] ),
    .A2(_10419_),
    .B1(_10425_),
    .C1(_10427_),
    .X(_00248_));
 sky130_fd_sc_hd__nand2_2 _14292_ (.A(_09993_),
    .B(_10420_),
    .Y(_10428_));
 sky130_fd_sc_hd__o211a_2 _14293_ (.A1(\decode.regfile.registers_29[5] ),
    .A2(_10419_),
    .B1(_10428_),
    .C1(_10427_),
    .X(_00249_));
 sky130_fd_sc_hd__nand2_2 _14294_ (.A(_09999_),
    .B(_10420_),
    .Y(_10429_));
 sky130_fd_sc_hd__o211a_2 _14295_ (.A1(\decode.regfile.registers_29[6] ),
    .A2(_10419_),
    .B1(_10429_),
    .C1(_10427_),
    .X(_00250_));
 sky130_fd_sc_hd__nand2_2 _14296_ (.A(_10008_),
    .B(_10420_),
    .Y(_10430_));
 sky130_fd_sc_hd__o211a_2 _14297_ (.A1(\decode.regfile.registers_29[7] ),
    .A2(_10419_),
    .B1(_10430_),
    .C1(_10427_),
    .X(_00251_));
 sky130_fd_sc_hd__buf_1 _14298_ (.A(_10418_),
    .X(_10431_));
 sky130_fd_sc_hd__nand2_2 _14299_ (.A(_10015_),
    .B(_10431_),
    .Y(_10432_));
 sky130_fd_sc_hd__o211a_2 _14300_ (.A1(\decode.regfile.registers_29[8] ),
    .A2(_10419_),
    .B1(_10432_),
    .C1(_10427_),
    .X(_00252_));
 sky130_fd_sc_hd__nand2_2 _14301_ (.A(_10025_),
    .B(_10431_),
    .Y(_10433_));
 sky130_fd_sc_hd__o211a_2 _14302_ (.A1(\decode.regfile.registers_29[9] ),
    .A2(_10419_),
    .B1(_10433_),
    .C1(_10427_),
    .X(_00253_));
 sky130_fd_sc_hd__buf_1 _14303_ (.A(_10418_),
    .X(_10434_));
 sky130_fd_sc_hd__nand2_2 _14304_ (.A(_10031_),
    .B(_10431_),
    .Y(_10435_));
 sky130_fd_sc_hd__o211a_2 _14305_ (.A1(\decode.regfile.registers_29[10] ),
    .A2(_10434_),
    .B1(_10435_),
    .C1(_10427_),
    .X(_00254_));
 sky130_fd_sc_hd__nand2_2 _14306_ (.A(_10036_),
    .B(_10431_),
    .Y(_10436_));
 sky130_fd_sc_hd__o211a_2 _14307_ (.A1(\decode.regfile.registers_29[11] ),
    .A2(_10434_),
    .B1(_10436_),
    .C1(_10427_),
    .X(_00255_));
 sky130_fd_sc_hd__nand2_2 _14308_ (.A(_10042_),
    .B(_10431_),
    .Y(_10437_));
 sky130_fd_sc_hd__o211a_2 _14309_ (.A1(\decode.regfile.registers_29[12] ),
    .A2(_10434_),
    .B1(_10437_),
    .C1(_10427_),
    .X(_00256_));
 sky130_fd_sc_hd__nand2_2 _14310_ (.A(_10048_),
    .B(_10431_),
    .Y(_10438_));
 sky130_fd_sc_hd__o211a_2 _14311_ (.A1(\decode.regfile.registers_29[13] ),
    .A2(_10434_),
    .B1(_10438_),
    .C1(_10427_),
    .X(_00257_));
 sky130_fd_sc_hd__nand2_2 _14312_ (.A(_10053_),
    .B(_10431_),
    .Y(_10439_));
 sky130_fd_sc_hd__buf_1 _14313_ (.A(_10426_),
    .X(_10440_));
 sky130_fd_sc_hd__o211a_2 _14314_ (.A1(\decode.regfile.registers_29[14] ),
    .A2(_10434_),
    .B1(_10439_),
    .C1(_10440_),
    .X(_00258_));
 sky130_fd_sc_hd__nand2_2 _14315_ (.A(_10058_),
    .B(_10431_),
    .Y(_10441_));
 sky130_fd_sc_hd__o211a_2 _14316_ (.A1(\decode.regfile.registers_29[15] ),
    .A2(_10434_),
    .B1(_10441_),
    .C1(_10440_),
    .X(_00259_));
 sky130_fd_sc_hd__nand2_2 _14317_ (.A(_10064_),
    .B(_10431_),
    .Y(_10442_));
 sky130_fd_sc_hd__o211a_2 _14318_ (.A1(\decode.regfile.registers_29[16] ),
    .A2(_10434_),
    .B1(_10442_),
    .C1(_10440_),
    .X(_00260_));
 sky130_fd_sc_hd__nand2_2 _14319_ (.A(_10069_),
    .B(_10431_),
    .Y(_10443_));
 sky130_fd_sc_hd__o211a_2 _14320_ (.A1(\decode.regfile.registers_29[17] ),
    .A2(_10434_),
    .B1(_10443_),
    .C1(_10440_),
    .X(_00261_));
 sky130_fd_sc_hd__buf_1 _14321_ (.A(_10418_),
    .X(_10444_));
 sky130_fd_sc_hd__nand2_2 _14322_ (.A(_10074_),
    .B(_10444_),
    .Y(_10445_));
 sky130_fd_sc_hd__o211a_2 _14323_ (.A1(\decode.regfile.registers_29[18] ),
    .A2(_10434_),
    .B1(_10445_),
    .C1(_10440_),
    .X(_00262_));
 sky130_fd_sc_hd__nand2_2 _14324_ (.A(_10081_),
    .B(_10444_),
    .Y(_10446_));
 sky130_fd_sc_hd__o211a_2 _14325_ (.A1(\decode.regfile.registers_29[19] ),
    .A2(_10434_),
    .B1(_10446_),
    .C1(_10440_),
    .X(_00263_));
 sky130_fd_sc_hd__buf_1 _14326_ (.A(_10418_),
    .X(_10447_));
 sky130_fd_sc_hd__nand2_2 _14327_ (.A(_10087_),
    .B(_10444_),
    .Y(_10448_));
 sky130_fd_sc_hd__o211a_2 _14328_ (.A1(\decode.regfile.registers_29[20] ),
    .A2(_10447_),
    .B1(_10448_),
    .C1(_10440_),
    .X(_00264_));
 sky130_fd_sc_hd__nand2_2 _14329_ (.A(_10092_),
    .B(_10444_),
    .Y(_10449_));
 sky130_fd_sc_hd__o211a_2 _14330_ (.A1(\decode.regfile.registers_29[21] ),
    .A2(_10447_),
    .B1(_10449_),
    .C1(_10440_),
    .X(_00265_));
 sky130_fd_sc_hd__nand2_2 _14331_ (.A(_10097_),
    .B(_10444_),
    .Y(_10450_));
 sky130_fd_sc_hd__o211a_2 _14332_ (.A1(\decode.regfile.registers_29[22] ),
    .A2(_10447_),
    .B1(_10450_),
    .C1(_10440_),
    .X(_00266_));
 sky130_fd_sc_hd__nand2_2 _14333_ (.A(_10102_),
    .B(_10444_),
    .Y(_10451_));
 sky130_fd_sc_hd__o211a_2 _14334_ (.A1(\decode.regfile.registers_29[23] ),
    .A2(_10447_),
    .B1(_10451_),
    .C1(_10440_),
    .X(_00267_));
 sky130_fd_sc_hd__nand2_2 _14335_ (.A(_10107_),
    .B(_10444_),
    .Y(_10452_));
 sky130_fd_sc_hd__buf_1 _14336_ (.A(_10426_),
    .X(_10453_));
 sky130_fd_sc_hd__o211a_2 _14337_ (.A1(\decode.regfile.registers_29[24] ),
    .A2(_10447_),
    .B1(_10452_),
    .C1(_10453_),
    .X(_00268_));
 sky130_fd_sc_hd__nand2_2 _14338_ (.A(_10112_),
    .B(_10444_),
    .Y(_10454_));
 sky130_fd_sc_hd__o211a_2 _14339_ (.A1(\decode.regfile.registers_29[25] ),
    .A2(_10447_),
    .B1(_10454_),
    .C1(_10453_),
    .X(_00269_));
 sky130_fd_sc_hd__nand2_2 _14340_ (.A(_10117_),
    .B(_10444_),
    .Y(_10455_));
 sky130_fd_sc_hd__o211a_2 _14341_ (.A1(\decode.regfile.registers_29[26] ),
    .A2(_10447_),
    .B1(_10455_),
    .C1(_10453_),
    .X(_00270_));
 sky130_fd_sc_hd__nand2_2 _14342_ (.A(_10122_),
    .B(_10444_),
    .Y(_10456_));
 sky130_fd_sc_hd__o211a_2 _14343_ (.A1(\decode.regfile.registers_29[27] ),
    .A2(_10447_),
    .B1(_10456_),
    .C1(_10453_),
    .X(_00271_));
 sky130_fd_sc_hd__nand2_2 _14344_ (.A(_10128_),
    .B(_10418_),
    .Y(_10457_));
 sky130_fd_sc_hd__o211a_2 _14345_ (.A1(\decode.regfile.registers_29[28] ),
    .A2(_10447_),
    .B1(_10457_),
    .C1(_10453_),
    .X(_00272_));
 sky130_fd_sc_hd__nand2_2 _14346_ (.A(_10136_),
    .B(_10418_),
    .Y(_10458_));
 sky130_fd_sc_hd__o211a_2 _14347_ (.A1(\decode.regfile.registers_29[29] ),
    .A2(_10447_),
    .B1(_10458_),
    .C1(_10453_),
    .X(_00273_));
 sky130_fd_sc_hd__nand2_2 _14348_ (.A(_10142_),
    .B(_10418_),
    .Y(_10459_));
 sky130_fd_sc_hd__o211a_2 _14349_ (.A1(\decode.regfile.registers_29[30] ),
    .A2(_10420_),
    .B1(_10459_),
    .C1(_10453_),
    .X(_00274_));
 sky130_fd_sc_hd__nand2_2 _14350_ (.A(_10147_),
    .B(_10418_),
    .Y(_10460_));
 sky130_fd_sc_hd__o211a_2 _14351_ (.A1(\decode.regfile.registers_29[31] ),
    .A2(_10420_),
    .B1(_10460_),
    .C1(_10453_),
    .X(_00275_));
 sky130_fd_sc_hd__and4_2 _14352_ (.A(_10373_),
    .B(_10195_),
    .C(_09932_),
    .D(_10149_),
    .X(_10461_));
 sky130_fd_sc_hd__buf_1 _14353_ (.A(_10461_),
    .X(_10462_));
 sky130_fd_sc_hd__buf_1 _14354_ (.A(_10462_),
    .X(_10463_));
 sky130_fd_sc_hd__buf_1 _14355_ (.A(_10462_),
    .X(_10464_));
 sky130_fd_sc_hd__nand2_2 _14356_ (.A(_09950_),
    .B(_10464_),
    .Y(_10465_));
 sky130_fd_sc_hd__o211a_2 _14357_ (.A1(\decode.regfile.registers_30[0] ),
    .A2(_10463_),
    .B1(_10465_),
    .C1(_10453_),
    .X(_00276_));
 sky130_fd_sc_hd__nand2_2 _14358_ (.A(_09964_),
    .B(_10464_),
    .Y(_10466_));
 sky130_fd_sc_hd__o211a_2 _14359_ (.A1(\decode.regfile.registers_30[1] ),
    .A2(_10463_),
    .B1(_10466_),
    .C1(_10453_),
    .X(_00277_));
 sky130_fd_sc_hd__nand2_2 _14360_ (.A(_09970_),
    .B(_10464_),
    .Y(_10467_));
 sky130_fd_sc_hd__buf_1 _14361_ (.A(_10426_),
    .X(_10468_));
 sky130_fd_sc_hd__o211a_2 _14362_ (.A1(\decode.regfile.registers_30[2] ),
    .A2(_10463_),
    .B1(_10467_),
    .C1(_10468_),
    .X(_00278_));
 sky130_fd_sc_hd__nand2_2 _14363_ (.A(_09975_),
    .B(_10464_),
    .Y(_10469_));
 sky130_fd_sc_hd__o211a_2 _14364_ (.A1(\decode.regfile.registers_30[3] ),
    .A2(_10463_),
    .B1(_10469_),
    .C1(_10468_),
    .X(_00279_));
 sky130_fd_sc_hd__nand2_2 _14365_ (.A(_09984_),
    .B(_10464_),
    .Y(_10470_));
 sky130_fd_sc_hd__o211a_2 _14366_ (.A1(\decode.regfile.registers_30[4] ),
    .A2(_10463_),
    .B1(_10470_),
    .C1(_10468_),
    .X(_00280_));
 sky130_fd_sc_hd__nand2_2 _14367_ (.A(_09993_),
    .B(_10464_),
    .Y(_10471_));
 sky130_fd_sc_hd__o211a_2 _14368_ (.A1(\decode.regfile.registers_30[5] ),
    .A2(_10463_),
    .B1(_10471_),
    .C1(_10468_),
    .X(_00281_));
 sky130_fd_sc_hd__nand2_2 _14369_ (.A(_09999_),
    .B(_10464_),
    .Y(_10472_));
 sky130_fd_sc_hd__o211a_2 _14370_ (.A1(\decode.regfile.registers_30[6] ),
    .A2(_10463_),
    .B1(_10472_),
    .C1(_10468_),
    .X(_00282_));
 sky130_fd_sc_hd__nand2_2 _14371_ (.A(_10008_),
    .B(_10464_),
    .Y(_10473_));
 sky130_fd_sc_hd__o211a_2 _14372_ (.A1(\decode.regfile.registers_30[7] ),
    .A2(_10463_),
    .B1(_10473_),
    .C1(_10468_),
    .X(_00283_));
 sky130_fd_sc_hd__buf_1 _14373_ (.A(_10462_),
    .X(_10474_));
 sky130_fd_sc_hd__nand2_2 _14374_ (.A(_10015_),
    .B(_10474_),
    .Y(_10475_));
 sky130_fd_sc_hd__o211a_2 _14375_ (.A1(\decode.regfile.registers_30[8] ),
    .A2(_10463_),
    .B1(_10475_),
    .C1(_10468_),
    .X(_00284_));
 sky130_fd_sc_hd__nand2_2 _14376_ (.A(_10025_),
    .B(_10474_),
    .Y(_10476_));
 sky130_fd_sc_hd__o211a_2 _14377_ (.A1(\decode.regfile.registers_30[9] ),
    .A2(_10463_),
    .B1(_10476_),
    .C1(_10468_),
    .X(_00285_));
 sky130_fd_sc_hd__buf_1 _14378_ (.A(_10462_),
    .X(_10477_));
 sky130_fd_sc_hd__nand2_2 _14379_ (.A(_10031_),
    .B(_10474_),
    .Y(_10478_));
 sky130_fd_sc_hd__o211a_2 _14380_ (.A1(\decode.regfile.registers_30[10] ),
    .A2(_10477_),
    .B1(_10478_),
    .C1(_10468_),
    .X(_00286_));
 sky130_fd_sc_hd__nand2_2 _14381_ (.A(_10036_),
    .B(_10474_),
    .Y(_10479_));
 sky130_fd_sc_hd__o211a_2 _14382_ (.A1(\decode.regfile.registers_30[11] ),
    .A2(_10477_),
    .B1(_10479_),
    .C1(_10468_),
    .X(_00287_));
 sky130_fd_sc_hd__nand2_2 _14383_ (.A(_10042_),
    .B(_10474_),
    .Y(_10480_));
 sky130_fd_sc_hd__buf_1 _14384_ (.A(_10426_),
    .X(_10481_));
 sky130_fd_sc_hd__o211a_2 _14385_ (.A1(\decode.regfile.registers_30[12] ),
    .A2(_10477_),
    .B1(_10480_),
    .C1(_10481_),
    .X(_00288_));
 sky130_fd_sc_hd__nand2_2 _14386_ (.A(_10048_),
    .B(_10474_),
    .Y(_10482_));
 sky130_fd_sc_hd__o211a_2 _14387_ (.A1(\decode.regfile.registers_30[13] ),
    .A2(_10477_),
    .B1(_10482_),
    .C1(_10481_),
    .X(_00289_));
 sky130_fd_sc_hd__nand2_2 _14388_ (.A(_10053_),
    .B(_10474_),
    .Y(_10483_));
 sky130_fd_sc_hd__o211a_2 _14389_ (.A1(\decode.regfile.registers_30[14] ),
    .A2(_10477_),
    .B1(_10483_),
    .C1(_10481_),
    .X(_00290_));
 sky130_fd_sc_hd__nand2_2 _14390_ (.A(_10058_),
    .B(_10474_),
    .Y(_10484_));
 sky130_fd_sc_hd__o211a_2 _14391_ (.A1(\decode.regfile.registers_30[15] ),
    .A2(_10477_),
    .B1(_10484_),
    .C1(_10481_),
    .X(_00291_));
 sky130_fd_sc_hd__nand2_2 _14392_ (.A(_10064_),
    .B(_10474_),
    .Y(_10485_));
 sky130_fd_sc_hd__o211a_2 _14393_ (.A1(\decode.regfile.registers_30[16] ),
    .A2(_10477_),
    .B1(_10485_),
    .C1(_10481_),
    .X(_00292_));
 sky130_fd_sc_hd__nand2_2 _14394_ (.A(_10069_),
    .B(_10474_),
    .Y(_10486_));
 sky130_fd_sc_hd__o211a_2 _14395_ (.A1(\decode.regfile.registers_30[17] ),
    .A2(_10477_),
    .B1(_10486_),
    .C1(_10481_),
    .X(_00293_));
 sky130_fd_sc_hd__buf_1 _14396_ (.A(_10462_),
    .X(_10487_));
 sky130_fd_sc_hd__nand2_2 _14397_ (.A(_10074_),
    .B(_10487_),
    .Y(_10488_));
 sky130_fd_sc_hd__o211a_2 _14398_ (.A1(\decode.regfile.registers_30[18] ),
    .A2(_10477_),
    .B1(_10488_),
    .C1(_10481_),
    .X(_00294_));
 sky130_fd_sc_hd__nand2_2 _14399_ (.A(_10081_),
    .B(_10487_),
    .Y(_10489_));
 sky130_fd_sc_hd__o211a_2 _14400_ (.A1(\decode.regfile.registers_30[19] ),
    .A2(_10477_),
    .B1(_10489_),
    .C1(_10481_),
    .X(_00295_));
 sky130_fd_sc_hd__buf_1 _14401_ (.A(_10462_),
    .X(_10490_));
 sky130_fd_sc_hd__nand2_2 _14402_ (.A(_10087_),
    .B(_10487_),
    .Y(_10491_));
 sky130_fd_sc_hd__o211a_2 _14403_ (.A1(\decode.regfile.registers_30[20] ),
    .A2(_10490_),
    .B1(_10491_),
    .C1(_10481_),
    .X(_00296_));
 sky130_fd_sc_hd__nand2_2 _14404_ (.A(_10092_),
    .B(_10487_),
    .Y(_10492_));
 sky130_fd_sc_hd__o211a_2 _14405_ (.A1(\decode.regfile.registers_30[21] ),
    .A2(_10490_),
    .B1(_10492_),
    .C1(_10481_),
    .X(_00297_));
 sky130_fd_sc_hd__nand2_2 _14406_ (.A(_10097_),
    .B(_10487_),
    .Y(_10493_));
 sky130_fd_sc_hd__buf_1 _14407_ (.A(_10426_),
    .X(_10494_));
 sky130_fd_sc_hd__o211a_2 _14408_ (.A1(\decode.regfile.registers_30[22] ),
    .A2(_10490_),
    .B1(_10493_),
    .C1(_10494_),
    .X(_00298_));
 sky130_fd_sc_hd__nand2_2 _14409_ (.A(_10102_),
    .B(_10487_),
    .Y(_10495_));
 sky130_fd_sc_hd__o211a_2 _14410_ (.A1(\decode.regfile.registers_30[23] ),
    .A2(_10490_),
    .B1(_10495_),
    .C1(_10494_),
    .X(_00299_));
 sky130_fd_sc_hd__nand2_2 _14411_ (.A(_10107_),
    .B(_10487_),
    .Y(_10496_));
 sky130_fd_sc_hd__o211a_2 _14412_ (.A1(\decode.regfile.registers_30[24] ),
    .A2(_10490_),
    .B1(_10496_),
    .C1(_10494_),
    .X(_00300_));
 sky130_fd_sc_hd__nand2_2 _14413_ (.A(_10112_),
    .B(_10487_),
    .Y(_10497_));
 sky130_fd_sc_hd__o211a_2 _14414_ (.A1(\decode.regfile.registers_30[25] ),
    .A2(_10490_),
    .B1(_10497_),
    .C1(_10494_),
    .X(_00301_));
 sky130_fd_sc_hd__nand2_2 _14415_ (.A(_10117_),
    .B(_10487_),
    .Y(_10498_));
 sky130_fd_sc_hd__o211a_2 _14416_ (.A1(\decode.regfile.registers_30[26] ),
    .A2(_10490_),
    .B1(_10498_),
    .C1(_10494_),
    .X(_00302_));
 sky130_fd_sc_hd__nand2_2 _14417_ (.A(_10122_),
    .B(_10487_),
    .Y(_10499_));
 sky130_fd_sc_hd__o211a_2 _14418_ (.A1(\decode.regfile.registers_30[27] ),
    .A2(_10490_),
    .B1(_10499_),
    .C1(_10494_),
    .X(_00303_));
 sky130_fd_sc_hd__nand2_2 _14419_ (.A(_10128_),
    .B(_10462_),
    .Y(_10500_));
 sky130_fd_sc_hd__o211a_2 _14420_ (.A1(\decode.regfile.registers_30[28] ),
    .A2(_10490_),
    .B1(_10500_),
    .C1(_10494_),
    .X(_00304_));
 sky130_fd_sc_hd__nand2_2 _14421_ (.A(_10136_),
    .B(_10462_),
    .Y(_10501_));
 sky130_fd_sc_hd__o211a_2 _14422_ (.A1(\decode.regfile.registers_30[29] ),
    .A2(_10490_),
    .B1(_10501_),
    .C1(_10494_),
    .X(_00305_));
 sky130_fd_sc_hd__nand2_2 _14423_ (.A(_10142_),
    .B(_10462_),
    .Y(_10502_));
 sky130_fd_sc_hd__o211a_2 _14424_ (.A1(\decode.regfile.registers_30[30] ),
    .A2(_10464_),
    .B1(_10502_),
    .C1(_10494_),
    .X(_00306_));
 sky130_fd_sc_hd__nand2_2 _14425_ (.A(_10147_),
    .B(_10462_),
    .Y(_10503_));
 sky130_fd_sc_hd__o211a_2 _14426_ (.A1(\decode.regfile.registers_30[31] ),
    .A2(_10464_),
    .B1(_10503_),
    .C1(_10494_),
    .X(_00307_));
 sky130_fd_sc_hd__and4_2 _14427_ (.A(_10373_),
    .B(_10195_),
    .C(_09933_),
    .D(_10150_),
    .X(_10504_));
 sky130_fd_sc_hd__buf_1 _14428_ (.A(_10504_),
    .X(_10505_));
 sky130_fd_sc_hd__buf_1 _14429_ (.A(_10505_),
    .X(_10506_));
 sky130_fd_sc_hd__buf_1 _14430_ (.A(_10505_),
    .X(_10507_));
 sky130_fd_sc_hd__nand2_2 _14431_ (.A(_09950_),
    .B(_10507_),
    .Y(_10508_));
 sky130_fd_sc_hd__buf_1 _14432_ (.A(_10426_),
    .X(_10509_));
 sky130_fd_sc_hd__o211a_2 _14433_ (.A1(\decode.regfile.registers_31[0] ),
    .A2(_10506_),
    .B1(_10508_),
    .C1(_10509_),
    .X(_00308_));
 sky130_fd_sc_hd__nand2_2 _14434_ (.A(_09964_),
    .B(_10507_),
    .Y(_10510_));
 sky130_fd_sc_hd__o211a_2 _14435_ (.A1(\decode.regfile.registers_31[1] ),
    .A2(_10506_),
    .B1(_10510_),
    .C1(_10509_),
    .X(_00309_));
 sky130_fd_sc_hd__nand2_2 _14436_ (.A(_09970_),
    .B(_10507_),
    .Y(_10511_));
 sky130_fd_sc_hd__o211a_2 _14437_ (.A1(\decode.regfile.registers_31[2] ),
    .A2(_10506_),
    .B1(_10511_),
    .C1(_10509_),
    .X(_00310_));
 sky130_fd_sc_hd__nand2_2 _14438_ (.A(_09975_),
    .B(_10507_),
    .Y(_10512_));
 sky130_fd_sc_hd__o211a_2 _14439_ (.A1(\decode.regfile.registers_31[3] ),
    .A2(_10506_),
    .B1(_10512_),
    .C1(_10509_),
    .X(_00311_));
 sky130_fd_sc_hd__nand2_2 _14440_ (.A(_09984_),
    .B(_10507_),
    .Y(_10513_));
 sky130_fd_sc_hd__o211a_2 _14441_ (.A1(\decode.regfile.registers_31[4] ),
    .A2(_10506_),
    .B1(_10513_),
    .C1(_10509_),
    .X(_00312_));
 sky130_fd_sc_hd__nand2_2 _14442_ (.A(_09993_),
    .B(_10507_),
    .Y(_10514_));
 sky130_fd_sc_hd__o211a_2 _14443_ (.A1(\decode.regfile.registers_31[5] ),
    .A2(_10506_),
    .B1(_10514_),
    .C1(_10509_),
    .X(_00313_));
 sky130_fd_sc_hd__nand2_2 _14444_ (.A(_09999_),
    .B(_10507_),
    .Y(_10515_));
 sky130_fd_sc_hd__o211a_2 _14445_ (.A1(\decode.regfile.registers_31[6] ),
    .A2(_10506_),
    .B1(_10515_),
    .C1(_10509_),
    .X(_00314_));
 sky130_fd_sc_hd__nand2_2 _14446_ (.A(_10008_),
    .B(_10507_),
    .Y(_10516_));
 sky130_fd_sc_hd__o211a_2 _14447_ (.A1(\decode.regfile.registers_31[7] ),
    .A2(_10506_),
    .B1(_10516_),
    .C1(_10509_),
    .X(_00315_));
 sky130_fd_sc_hd__buf_1 _14448_ (.A(_10505_),
    .X(_10517_));
 sky130_fd_sc_hd__nand2_2 _14449_ (.A(_10015_),
    .B(_10517_),
    .Y(_10518_));
 sky130_fd_sc_hd__o211a_2 _14450_ (.A1(\decode.regfile.registers_31[8] ),
    .A2(_10506_),
    .B1(_10518_),
    .C1(_10509_),
    .X(_00316_));
 sky130_fd_sc_hd__nand2_2 _14451_ (.A(_10025_),
    .B(_10517_),
    .Y(_10519_));
 sky130_fd_sc_hd__o211a_2 _14452_ (.A1(\decode.regfile.registers_31[9] ),
    .A2(_10506_),
    .B1(_10519_),
    .C1(_10509_),
    .X(_00317_));
 sky130_fd_sc_hd__buf_1 _14453_ (.A(_10505_),
    .X(_10520_));
 sky130_fd_sc_hd__nand2_2 _14454_ (.A(_10031_),
    .B(_10517_),
    .Y(_10521_));
 sky130_fd_sc_hd__buf_1 _14455_ (.A(_10426_),
    .X(_10522_));
 sky130_fd_sc_hd__o211a_2 _14456_ (.A1(\decode.regfile.registers_31[10] ),
    .A2(_10520_),
    .B1(_10521_),
    .C1(_10522_),
    .X(_00318_));
 sky130_fd_sc_hd__nand2_2 _14457_ (.A(_10036_),
    .B(_10517_),
    .Y(_10523_));
 sky130_fd_sc_hd__o211a_2 _14458_ (.A1(\decode.regfile.registers_31[11] ),
    .A2(_10520_),
    .B1(_10523_),
    .C1(_10522_),
    .X(_00319_));
 sky130_fd_sc_hd__nand2_2 _14459_ (.A(_10042_),
    .B(_10517_),
    .Y(_10524_));
 sky130_fd_sc_hd__o211a_2 _14460_ (.A1(\decode.regfile.registers_31[12] ),
    .A2(_10520_),
    .B1(_10524_),
    .C1(_10522_),
    .X(_00320_));
 sky130_fd_sc_hd__nand2_2 _14461_ (.A(_10048_),
    .B(_10517_),
    .Y(_10525_));
 sky130_fd_sc_hd__o211a_2 _14462_ (.A1(\decode.regfile.registers_31[13] ),
    .A2(_10520_),
    .B1(_10525_),
    .C1(_10522_),
    .X(_00321_));
 sky130_fd_sc_hd__nand2_2 _14463_ (.A(_10053_),
    .B(_10517_),
    .Y(_10526_));
 sky130_fd_sc_hd__o211a_2 _14464_ (.A1(\decode.regfile.registers_31[14] ),
    .A2(_10520_),
    .B1(_10526_),
    .C1(_10522_),
    .X(_00322_));
 sky130_fd_sc_hd__nand2_2 _14465_ (.A(_10058_),
    .B(_10517_),
    .Y(_10527_));
 sky130_fd_sc_hd__o211a_2 _14466_ (.A1(\decode.regfile.registers_31[15] ),
    .A2(_10520_),
    .B1(_10527_),
    .C1(_10522_),
    .X(_00323_));
 sky130_fd_sc_hd__nand2_2 _14467_ (.A(_10064_),
    .B(_10517_),
    .Y(_10528_));
 sky130_fd_sc_hd__o211a_2 _14468_ (.A1(\decode.regfile.registers_31[16] ),
    .A2(_10520_),
    .B1(_10528_),
    .C1(_10522_),
    .X(_00324_));
 sky130_fd_sc_hd__nand2_2 _14469_ (.A(_10069_),
    .B(_10517_),
    .Y(_10529_));
 sky130_fd_sc_hd__o211a_2 _14470_ (.A1(\decode.regfile.registers_31[17] ),
    .A2(_10520_),
    .B1(_10529_),
    .C1(_10522_),
    .X(_00325_));
 sky130_fd_sc_hd__buf_1 _14471_ (.A(_10505_),
    .X(_10530_));
 sky130_fd_sc_hd__nand2_2 _14472_ (.A(_10074_),
    .B(_10530_),
    .Y(_10531_));
 sky130_fd_sc_hd__o211a_2 _14473_ (.A1(\decode.regfile.registers_31[18] ),
    .A2(_10520_),
    .B1(_10531_),
    .C1(_10522_),
    .X(_00326_));
 sky130_fd_sc_hd__nand2_2 _14474_ (.A(_10081_),
    .B(_10530_),
    .Y(_10532_));
 sky130_fd_sc_hd__o211a_2 _14475_ (.A1(\decode.regfile.registers_31[19] ),
    .A2(_10520_),
    .B1(_10532_),
    .C1(_10522_),
    .X(_00327_));
 sky130_fd_sc_hd__buf_1 _14476_ (.A(_10505_),
    .X(_10533_));
 sky130_fd_sc_hd__nand2_2 _14477_ (.A(_10087_),
    .B(_10530_),
    .Y(_10534_));
 sky130_fd_sc_hd__buf_1 _14478_ (.A(_10426_),
    .X(_10535_));
 sky130_fd_sc_hd__o211a_2 _14479_ (.A1(\decode.regfile.registers_31[20] ),
    .A2(_10533_),
    .B1(_10534_),
    .C1(_10535_),
    .X(_00328_));
 sky130_fd_sc_hd__nand2_2 _14480_ (.A(_10092_),
    .B(_10530_),
    .Y(_10536_));
 sky130_fd_sc_hd__o211a_2 _14481_ (.A1(\decode.regfile.registers_31[21] ),
    .A2(_10533_),
    .B1(_10536_),
    .C1(_10535_),
    .X(_00329_));
 sky130_fd_sc_hd__nand2_2 _14482_ (.A(_10097_),
    .B(_10530_),
    .Y(_10537_));
 sky130_fd_sc_hd__o211a_2 _14483_ (.A1(\decode.regfile.registers_31[22] ),
    .A2(_10533_),
    .B1(_10537_),
    .C1(_10535_),
    .X(_00330_));
 sky130_fd_sc_hd__nand2_2 _14484_ (.A(_10102_),
    .B(_10530_),
    .Y(_10538_));
 sky130_fd_sc_hd__o211a_2 _14485_ (.A1(\decode.regfile.registers_31[23] ),
    .A2(_10533_),
    .B1(_10538_),
    .C1(_10535_),
    .X(_00331_));
 sky130_fd_sc_hd__nand2_2 _14486_ (.A(_10107_),
    .B(_10530_),
    .Y(_10539_));
 sky130_fd_sc_hd__o211a_2 _14487_ (.A1(\decode.regfile.registers_31[24] ),
    .A2(_10533_),
    .B1(_10539_),
    .C1(_10535_),
    .X(_00332_));
 sky130_fd_sc_hd__nand2_2 _14488_ (.A(_10112_),
    .B(_10530_),
    .Y(_10540_));
 sky130_fd_sc_hd__o211a_2 _14489_ (.A1(\decode.regfile.registers_31[25] ),
    .A2(_10533_),
    .B1(_10540_),
    .C1(_10535_),
    .X(_00333_));
 sky130_fd_sc_hd__nand2_2 _14490_ (.A(_10117_),
    .B(_10530_),
    .Y(_10541_));
 sky130_fd_sc_hd__o211a_2 _14491_ (.A1(\decode.regfile.registers_31[26] ),
    .A2(_10533_),
    .B1(_10541_),
    .C1(_10535_),
    .X(_00334_));
 sky130_fd_sc_hd__nand2_2 _14492_ (.A(_10122_),
    .B(_10530_),
    .Y(_10542_));
 sky130_fd_sc_hd__o211a_2 _14493_ (.A1(\decode.regfile.registers_31[27] ),
    .A2(_10533_),
    .B1(_10542_),
    .C1(_10535_),
    .X(_00335_));
 sky130_fd_sc_hd__nand2_2 _14494_ (.A(_10128_),
    .B(_10505_),
    .Y(_10543_));
 sky130_fd_sc_hd__o211a_2 _14495_ (.A1(\decode.regfile.registers_31[28] ),
    .A2(_10533_),
    .B1(_10543_),
    .C1(_10535_),
    .X(_00336_));
 sky130_fd_sc_hd__nand2_2 _14496_ (.A(_10136_),
    .B(_10505_),
    .Y(_10544_));
 sky130_fd_sc_hd__o211a_2 _14497_ (.A1(\decode.regfile.registers_31[29] ),
    .A2(_10533_),
    .B1(_10544_),
    .C1(_10535_),
    .X(_00337_));
 sky130_fd_sc_hd__nand2_2 _14498_ (.A(_10142_),
    .B(_10505_),
    .Y(_10545_));
 sky130_fd_sc_hd__buf_1 _14499_ (.A(_10426_),
    .X(_10546_));
 sky130_fd_sc_hd__o211a_2 _14500_ (.A1(\decode.regfile.registers_31[30] ),
    .A2(_10507_),
    .B1(_10545_),
    .C1(_10546_),
    .X(_00338_));
 sky130_fd_sc_hd__nand2_2 _14501_ (.A(_10147_),
    .B(_10505_),
    .Y(_10547_));
 sky130_fd_sc_hd__o211a_2 _14502_ (.A1(\decode.regfile.registers_31[31] ),
    .A2(_10507_),
    .B1(_10547_),
    .C1(_10546_),
    .X(_00339_));
 sky130_fd_sc_hd__mux4_2 _14503_ (.A0(\fetch.btb.btbTable[0][1] ),
    .A1(\fetch.btb.btbTable[1][1] ),
    .A2(\fetch.btb.btbTable[2][1] ),
    .A3(\fetch.btb.btbTable[3][1] ),
    .S0(_09891_),
    .S1(_09888_),
    .X(_10548_));
 sky130_fd_sc_hd__mux4_2 _14504_ (.A0(\fetch.btb.btbTable[4][1] ),
    .A1(\fetch.btb.btbTable[5][1] ),
    .A2(\fetch.btb.btbTable[6][1] ),
    .A3(\fetch.btb.btbTable[7][1] ),
    .S0(_09891_),
    .S1(_09888_),
    .X(_10549_));
 sky130_fd_sc_hd__a22o_2 _14505_ (.A1(_10548_),
    .A2(_09917_),
    .B1(_09916_),
    .B2(_10549_),
    .X(_10550_));
 sky130_fd_sc_hd__mux4_2 _14506_ (.A0(\fetch.btb.btbTable[12][1] ),
    .A1(\fetch.btb.btbTable[13][1] ),
    .A2(\fetch.btb.btbTable[14][1] ),
    .A3(\fetch.btb.btbTable[15][1] ),
    .S0(_09891_),
    .S1(_09888_),
    .X(_10551_));
 sky130_fd_sc_hd__mux4_2 _14507_ (.A0(\fetch.btb.btbTable[8][1] ),
    .A1(\fetch.btb.btbTable[9][1] ),
    .A2(\fetch.btb.btbTable[10][1] ),
    .A3(\fetch.btb.btbTable[11][1] ),
    .S0(_09891_),
    .S1(_09888_),
    .X(_10552_));
 sky130_fd_sc_hd__and3b_2 _14508_ (.A_N(_09879_),
    .B(_10552_),
    .C(_09882_),
    .X(_10553_));
 sky130_fd_sc_hd__a31o_2 _14509_ (.A1(_09879_),
    .A2(_09882_),
    .A3(_10551_),
    .B1(_10553_),
    .X(_10554_));
 sky130_fd_sc_hd__mux4_2 _14510_ (.A0(\fetch.btb.btbTable[0][0] ),
    .A1(\fetch.btb.btbTable[1][0] ),
    .A2(\fetch.btb.btbTable[2][0] ),
    .A3(\fetch.btb.btbTable[3][0] ),
    .S0(_09891_),
    .S1(_09888_),
    .X(_10555_));
 sky130_fd_sc_hd__buf_1 _14511_ (.A(_09891_),
    .X(_10556_));
 sky130_fd_sc_hd__buf_1 _14512_ (.A(_09888_),
    .X(_10557_));
 sky130_fd_sc_hd__mux4_2 _14513_ (.A0(\fetch.btb.btbTable[4][0] ),
    .A1(\fetch.btb.btbTable[5][0] ),
    .A2(\fetch.btb.btbTable[6][0] ),
    .A3(\fetch.btb.btbTable[7][0] ),
    .S0(_10556_),
    .S1(_10557_),
    .X(_10558_));
 sky130_fd_sc_hd__a22o_2 _14514_ (.A1(_10555_),
    .A2(_09917_),
    .B1(_09916_),
    .B2(_10558_),
    .X(_10559_));
 sky130_fd_sc_hd__mux4_2 _14515_ (.A0(\fetch.btb.btbTable[12][0] ),
    .A1(\fetch.btb.btbTable[13][0] ),
    .A2(\fetch.btb.btbTable[14][0] ),
    .A3(\fetch.btb.btbTable[15][0] ),
    .S0(_10556_),
    .S1(_10557_),
    .X(_10560_));
 sky130_fd_sc_hd__mux4_2 _14516_ (.A0(\fetch.btb.btbTable[8][0] ),
    .A1(\fetch.btb.btbTable[9][0] ),
    .A2(\fetch.btb.btbTable[10][0] ),
    .A3(\fetch.btb.btbTable[11][0] ),
    .S0(_09891_),
    .S1(_09888_),
    .X(_10561_));
 sky130_fd_sc_hd__and3b_2 _14517_ (.A_N(_09879_),
    .B(_10561_),
    .C(_09882_),
    .X(_10562_));
 sky130_fd_sc_hd__a31o_2 _14518_ (.A1(_09879_),
    .A2(_09882_),
    .A3(_10560_),
    .B1(_10562_),
    .X(_10563_));
 sky130_fd_sc_hd__o22ai_2 _14519_ (.A1(_10550_),
    .A2(_10554_),
    .B1(_10559_),
    .B2(_10563_),
    .Y(_10564_));
 sky130_fd_sc_hd__nand2_2 _14520_ (.A(_09900_),
    .B(\fetch.btb.io_branch ),
    .Y(_10565_));
 sky130_fd_sc_hd__nor4_2 _14521_ (.A(_10550_),
    .B(_10554_),
    .C(_10559_),
    .D(_10563_),
    .Y(_10566_));
 sky130_fd_sc_hd__nor2_2 _14522_ (.A(_10565_),
    .B(_10566_),
    .Y(_10567_));
 sky130_fd_sc_hd__a31o_2 _14523_ (.A1(\fetch.bht.bhtTable_tag_MPORT_en ),
    .A2(\fetch.btb.io_branch ),
    .A3(_10564_),
    .B1(_10567_),
    .X(_10568_));
 sky130_fd_sc_hd__nand2_2 _14524_ (.A(_10568_),
    .B(_09890_),
    .Y(_10569_));
 sky130_fd_sc_hd__or3b_2 _14525_ (.A(_10569_),
    .B(_09881_),
    .C_N(_09884_),
    .X(_10570_));
 sky130_fd_sc_hd__xnor2_2 _14526_ (.A(\fetch.btb.btbTable[9][0] ),
    .B(_10570_),
    .Y(_00340_));
 sky130_fd_sc_hd__nand3b_2 _14527_ (.A_N(_10566_),
    .B(_10565_),
    .C(_10564_),
    .Y(_10571_));
 sky130_fd_sc_hd__o21ai_2 _14528_ (.A1(_10565_),
    .A2(_10564_),
    .B1(_10571_),
    .Y(_10572_));
 sky130_fd_sc_hd__buf_1 _14529_ (.A(_10572_),
    .X(_10573_));
 sky130_fd_sc_hd__mux2_2 _14530_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[9][1] ),
    .S(_10570_),
    .X(_10574_));
 sky130_fd_sc_hd__buf_1 _14531_ (.A(_10574_),
    .X(_00341_));
 sky130_fd_sc_hd__buf_1 _14532_ (.A(reset),
    .X(_10575_));
 sky130_fd_sc_hd__buf_1 _14533_ (.A(_10575_),
    .X(_10576_));
 sky130_fd_sc_hd__buf_1 _14534_ (.A(_10576_),
    .X(_10577_));
 sky130_fd_sc_hd__or4bb_2 _14535_ (.A(\decode.control.io_opcode[3] ),
    .B(\decode.control.io_opcode[2] ),
    .C_N(\decode.control.io_opcode[1] ),
    .D_N(\decode.control.io_opcode[0] ),
    .X(_10578_));
 sky130_fd_sc_hd__buf_1 _14536_ (.A(\decode.control.io_opcode[6] ),
    .X(_10579_));
 sky130_fd_sc_hd__and4bb_2 _14537_ (.A_N(\decode.control.io_opcode[3] ),
    .B_N(\decode.control.io_opcode[2] ),
    .C(\decode.control.io_opcode[1] ),
    .D(\decode.control.io_opcode[0] ),
    .X(_10580_));
 sky130_fd_sc_hd__and4_2 _14538_ (.A(\decode.control.io_opcode[6] ),
    .B(\decode.control.io_opcode[5] ),
    .C(\decode.control.io_opcode[4] ),
    .D(_10580_),
    .X(_10581_));
 sky130_fd_sc_hd__o21ai_2 _14539_ (.A1(\decode.control.io_funct3[1] ),
    .A2(\decode.control.io_funct3[0] ),
    .B1(_10581_),
    .Y(_10582_));
 sky130_fd_sc_hd__and3b_2 _14540_ (.A_N(\decode.control.io_opcode[4] ),
    .B(\decode.control.io_opcode[5] ),
    .C(\decode.control.io_opcode[6] ),
    .X(_10583_));
 sky130_fd_sc_hd__and3_2 _14541_ (.A(\decode.control.io_opcode[2] ),
    .B(\decode.control.io_opcode[1] ),
    .C(\decode.control.io_opcode[0] ),
    .X(_10584_));
 sky130_fd_sc_hd__nand2_2 _14542_ (.A(_10583_),
    .B(_10584_),
    .Y(_10585_));
 sky130_fd_sc_hd__o2bb2a_2 _14543_ (.A1_N(_10580_),
    .A2_N(_10583_),
    .B1(\decode.control.io_opcode[3] ),
    .B2(_10585_),
    .X(_10586_));
 sky130_fd_sc_hd__o221a_2 _14544_ (.A1(_10578_),
    .A2(_10579_),
    .B1(\decode.control.io_funct3[2] ),
    .B2(_10582_),
    .C1(_10586_),
    .X(_10587_));
 sky130_fd_sc_hd__buf_1 _14545_ (.A(\decode.immGen._imm_T_24[17] ),
    .X(_10588_));
 sky130_fd_sc_hd__buf_1 _14546_ (.A(_10588_),
    .X(_10589_));
 sky130_fd_sc_hd__xor2_2 _14547_ (.A(_10589_),
    .B(\decode.id_ex_ex_rd_reg[2] ),
    .X(_10590_));
 sky130_fd_sc_hd__inv_2 _14548_ (.A(\decode.immGen._imm_T_24[19] ),
    .Y(_10591_));
 sky130_fd_sc_hd__buf_1 _14549_ (.A(_10591_),
    .X(_10592_));
 sky130_fd_sc_hd__buf_1 _14550_ (.A(_10592_),
    .X(_10593_));
 sky130_fd_sc_hd__buf_1 _14551_ (.A(_10593_),
    .X(_10594_));
 sky130_fd_sc_hd__buf_1 _14552_ (.A(_10594_),
    .X(_10595_));
 sky130_fd_sc_hd__inv_2 _14553_ (.A(\decode.id_ex_ex_rd_reg[3] ),
    .Y(_10596_));
 sky130_fd_sc_hd__buf_1 _14554_ (.A(\decode.immGen._imm_T_24[18] ),
    .X(_10597_));
 sky130_fd_sc_hd__buf_1 _14555_ (.A(_10597_),
    .X(_10598_));
 sky130_fd_sc_hd__buf_1 _14556_ (.A(_10598_),
    .X(_10599_));
 sky130_fd_sc_hd__a2bb2o_2 _14557_ (.A1_N(\decode.id_ex_ex_rd_reg[4] ),
    .A2_N(_10595_),
    .B1(_10596_),
    .B2(_10599_),
    .X(_10600_));
 sky130_fd_sc_hd__inv_2 _14558_ (.A(\decode.immGen._imm_T_24[16] ),
    .Y(_10601_));
 sky130_fd_sc_hd__buf_1 _14559_ (.A(_10601_),
    .X(_10602_));
 sky130_fd_sc_hd__buf_1 _14560_ (.A(_10602_),
    .X(_10603_));
 sky130_fd_sc_hd__buf_1 _14561_ (.A(_10603_),
    .X(_10604_));
 sky130_fd_sc_hd__inv_2 _14562_ (.A(\decode.immGen._imm_T_24[18] ),
    .Y(_10605_));
 sky130_fd_sc_hd__buf_1 _14563_ (.A(_10605_),
    .X(_10606_));
 sky130_fd_sc_hd__buf_1 _14564_ (.A(\decode.immGen._imm_T_24[16] ),
    .X(_10607_));
 sky130_fd_sc_hd__buf_1 _14565_ (.A(_10607_),
    .X(_10608_));
 sky130_fd_sc_hd__buf_1 _14566_ (.A(_10608_),
    .X(_10609_));
 sky130_fd_sc_hd__buf_1 _14567_ (.A(_10609_),
    .X(_10610_));
 sky130_fd_sc_hd__buf_1 _14568_ (.A(_10610_),
    .X(_10611_));
 sky130_fd_sc_hd__buf_1 _14569_ (.A(_10611_),
    .X(_10612_));
 sky130_fd_sc_hd__inv_2 _14570_ (.A(\decode.id_ex_ex_rd_reg[1] ),
    .Y(_10613_));
 sky130_fd_sc_hd__buf_1 _14571_ (.A(\decode.immGen._imm_T_24[15] ),
    .X(_10614_));
 sky130_fd_sc_hd__buf_1 _14572_ (.A(_10614_),
    .X(_10615_));
 sky130_fd_sc_hd__buf_1 _14573_ (.A(_10615_),
    .X(_10616_));
 sky130_fd_sc_hd__buf_1 _14574_ (.A(_10616_),
    .X(_10617_));
 sky130_fd_sc_hd__buf_1 _14575_ (.A(_10617_),
    .X(_10618_));
 sky130_fd_sc_hd__buf_1 _14576_ (.A(_10618_),
    .X(_10619_));
 sky130_fd_sc_hd__xor2_2 _14577_ (.A(_10619_),
    .B(\decode.id_ex_ex_rd_reg[0] ),
    .X(_10620_));
 sky130_fd_sc_hd__a221o_2 _14578_ (.A1(_10612_),
    .A2(_10613_),
    .B1(\decode.id_ex_ex_rd_reg[4] ),
    .B2(_10595_),
    .C1(_10620_),
    .X(_10621_));
 sky130_fd_sc_hd__a221o_2 _14579_ (.A1(_10604_),
    .A2(\decode.id_ex_ex_rd_reg[1] ),
    .B1(\decode.id_ex_ex_rd_reg[3] ),
    .B2(_10606_),
    .C1(_10621_),
    .X(_10622_));
 sky130_fd_sc_hd__inv_2 _14580_ (.A(\decode.immGen._imm_T_24[1] ),
    .Y(_10623_));
 sky130_fd_sc_hd__buf_1 _14581_ (.A(_10623_),
    .X(_10624_));
 sky130_fd_sc_hd__buf_1 _14582_ (.A(_10624_),
    .X(_10625_));
 sky130_fd_sc_hd__nand2_2 _14583_ (.A(_10625_),
    .B(_10613_),
    .Y(_10626_));
 sky130_fd_sc_hd__buf_1 _14584_ (.A(\decode.immGen._imm_T_24[1] ),
    .X(_10627_));
 sky130_fd_sc_hd__buf_1 _14585_ (.A(_10627_),
    .X(_10628_));
 sky130_fd_sc_hd__buf_1 _14586_ (.A(_10628_),
    .X(_10629_));
 sky130_fd_sc_hd__buf_1 _14587_ (.A(_10629_),
    .X(_10630_));
 sky130_fd_sc_hd__buf_1 _14588_ (.A(_10630_),
    .X(_10631_));
 sky130_fd_sc_hd__buf_1 _14589_ (.A(_10631_),
    .X(_10632_));
 sky130_fd_sc_hd__buf_1 _14590_ (.A(_10632_),
    .X(_10633_));
 sky130_fd_sc_hd__nand2_2 _14591_ (.A(_10633_),
    .B(\decode.id_ex_ex_rd_reg[1] ),
    .Y(_10634_));
 sky130_fd_sc_hd__buf_1 _14592_ (.A(\decode.immGen._imm_T_24[11] ),
    .X(_10635_));
 sky130_fd_sc_hd__buf_1 _14593_ (.A(_10635_),
    .X(_10636_));
 sky130_fd_sc_hd__buf_1 _14594_ (.A(_10636_),
    .X(_10637_));
 sky130_fd_sc_hd__buf_1 _14595_ (.A(_10637_),
    .X(_10638_));
 sky130_fd_sc_hd__buf_1 _14596_ (.A(_10638_),
    .X(_10639_));
 sky130_fd_sc_hd__buf_1 _14597_ (.A(_10639_),
    .X(_10640_));
 sky130_fd_sc_hd__or2_2 _14598_ (.A(_10640_),
    .B(\decode.id_ex_ex_rd_reg[0] ),
    .X(_10641_));
 sky130_fd_sc_hd__buf_1 _14599_ (.A(_10640_),
    .X(_10642_));
 sky130_fd_sc_hd__nand2_2 _14600_ (.A(_10642_),
    .B(\decode.id_ex_ex_rd_reg[0] ),
    .Y(_10643_));
 sky130_fd_sc_hd__a22o_2 _14601_ (.A1(_10626_),
    .A2(_10634_),
    .B1(_10641_),
    .B2(_10643_),
    .X(_10644_));
 sky130_fd_sc_hd__buf_1 _14602_ (.A(\decode.immGen._imm_T_24[4] ),
    .X(_10645_));
 sky130_fd_sc_hd__buf_1 _14603_ (.A(_10645_),
    .X(_10646_));
 sky130_fd_sc_hd__buf_1 _14604_ (.A(_10646_),
    .X(_10647_));
 sky130_fd_sc_hd__buf_1 _14605_ (.A(_10647_),
    .X(_10648_));
 sky130_fd_sc_hd__buf_1 _14606_ (.A(_10648_),
    .X(_10649_));
 sky130_fd_sc_hd__buf_1 _14607_ (.A(_10649_),
    .X(_10650_));
 sky130_fd_sc_hd__buf_1 _14608_ (.A(_10650_),
    .X(_10651_));
 sky130_fd_sc_hd__buf_1 _14609_ (.A(_10651_),
    .X(_10652_));
 sky130_fd_sc_hd__xor2_2 _14610_ (.A(_10652_),
    .B(\decode.id_ex_ex_rd_reg[4] ),
    .X(_10653_));
 sky130_fd_sc_hd__buf_1 _14611_ (.A(\decode.immGen._imm_T_24[2] ),
    .X(_10654_));
 sky130_fd_sc_hd__buf_1 _14612_ (.A(_10654_),
    .X(_10655_));
 sky130_fd_sc_hd__and2_2 _14613_ (.A(_10655_),
    .B(\decode.id_ex_ex_rd_reg[2] ),
    .X(_10656_));
 sky130_fd_sc_hd__buf_1 _14614_ (.A(_10655_),
    .X(_10657_));
 sky130_fd_sc_hd__nor2_2 _14615_ (.A(_10657_),
    .B(\decode.id_ex_ex_rd_reg[2] ),
    .Y(_10658_));
 sky130_fd_sc_hd__buf_1 _14616_ (.A(\decode.immGen._imm_T_24[3] ),
    .X(_10659_));
 sky130_fd_sc_hd__buf_1 _14617_ (.A(_10659_),
    .X(_10660_));
 sky130_fd_sc_hd__or2_2 _14618_ (.A(_10660_),
    .B(\decode.id_ex_ex_rd_reg[3] ),
    .X(_10661_));
 sky130_fd_sc_hd__buf_1 _14619_ (.A(_10660_),
    .X(_10662_));
 sky130_fd_sc_hd__nand2_2 _14620_ (.A(_10662_),
    .B(\decode.id_ex_ex_rd_reg[3] ),
    .Y(_10663_));
 sky130_fd_sc_hd__a2bb2o_2 _14621_ (.A1_N(_10656_),
    .A2_N(_10658_),
    .B1(_10661_),
    .B2(_10663_),
    .X(_10664_));
 sky130_fd_sc_hd__nor2_2 _14622_ (.A(\decode.control.io_opcode[6] ),
    .B(_10578_),
    .Y(_10665_));
 sky130_fd_sc_hd__and3b_2 _14623_ (.A_N(\decode.control.io_opcode[4] ),
    .B(_10580_),
    .C(\decode.control.io_opcode[5] ),
    .X(_10666_));
 sky130_fd_sc_hd__buf_1 _14624_ (.A(_10666_),
    .X(_10667_));
 sky130_fd_sc_hd__a31o_2 _14625_ (.A1(\decode.control.io_opcode[5] ),
    .A2(\decode.control.io_opcode[4] ),
    .A3(_10665_),
    .B1(_10667_),
    .X(_10668_));
 sky130_fd_sc_hd__or4b_2 _14626_ (.A(_10644_),
    .B(_10653_),
    .C(_10664_),
    .D_N(_10668_),
    .X(_10669_));
 sky130_fd_sc_hd__o41a_2 _14627_ (.A1(_10587_),
    .A2(_10590_),
    .A3(_10600_),
    .A4(_10622_),
    .B1(_10669_),
    .X(_10670_));
 sky130_fd_sc_hd__and2b_2 _14628_ (.A_N(_10670_),
    .B(\decode.id_ex_memread_reg ),
    .X(_10671_));
 sky130_fd_sc_hd__buf_1 _14629_ (.A(_10671_),
    .X(_10672_));
 sky130_fd_sc_hd__buf_1 _14630_ (.A(_10672_),
    .X(_10673_));
 sky130_fd_sc_hd__inv_2 _14631_ (.A(\execute.io_target_pc[1] ),
    .Y(_10674_));
 sky130_fd_sc_hd__inv_2 _14632_ (.A(\decode.id_ex_pc_reg[16] ),
    .Y(_10675_));
 sky130_fd_sc_hd__a22oi_2 _14633_ (.A1(_10674_),
    .A2(\decode.id_ex_pc_reg[1] ),
    .B1(_10675_),
    .B2(\execute.io_target_pc[16] ),
    .Y(_10676_));
 sky130_fd_sc_hd__inv_2 _14634_ (.A(\decode.id_ex_pc_reg[22] ),
    .Y(_10677_));
 sky130_fd_sc_hd__buf_1 _14635_ (.A(\decode.id_ex_pc_reg[6] ),
    .X(_10678_));
 sky130_fd_sc_hd__or2b_2 _14636_ (.A(\execute.io_target_pc[6] ),
    .B_N(_10678_),
    .X(_10679_));
 sky130_fd_sc_hd__inv_2 _14637_ (.A(\decode.id_ex_pc_reg[8] ),
    .Y(_10680_));
 sky130_fd_sc_hd__buf_1 _14638_ (.A(\decode.id_ex_pc_reg[15] ),
    .X(_10681_));
 sky130_fd_sc_hd__inv_2 _14639_ (.A(_10681_),
    .Y(_10682_));
 sky130_fd_sc_hd__a22oi_2 _14640_ (.A1(_10680_),
    .A2(\execute.io_target_pc[8] ),
    .B1(_10682_),
    .B2(\execute.io_target_pc[15] ),
    .Y(_10683_));
 sky130_fd_sc_hd__inv_2 _14641_ (.A(\decode.id_ex_pc_reg[30] ),
    .Y(_10684_));
 sky130_fd_sc_hd__o2bb2a_2 _14642_ (.A1_N(_10684_),
    .A2_N(\execute.io_target_pc[30] ),
    .B1(_10680_),
    .B2(\execute.io_target_pc[8] ),
    .X(_10685_));
 sky130_fd_sc_hd__o2111a_2 _14643_ (.A1(\execute.io_target_pc[22] ),
    .A2(_10677_),
    .B1(_10679_),
    .C1(_10683_),
    .D1(_10685_),
    .X(_10686_));
 sky130_fd_sc_hd__inv_2 _14644_ (.A(\execute.io_target_pc[27] ),
    .Y(_10687_));
 sky130_fd_sc_hd__inv_2 _14645_ (.A(\execute.io_target_pc[11] ),
    .Y(_10688_));
 sky130_fd_sc_hd__buf_1 _14646_ (.A(\decode.id_ex_pc_reg[11] ),
    .X(_10689_));
 sky130_fd_sc_hd__inv_2 _14647_ (.A(\decode.id_ex_pc_reg[4] ),
    .Y(_10690_));
 sky130_fd_sc_hd__o2bb2a_2 _14648_ (.A1_N(_10688_),
    .A2_N(_10689_),
    .B1(\execute.io_target_pc[4] ),
    .B2(_10690_),
    .X(_10691_));
 sky130_fd_sc_hd__inv_2 _14649_ (.A(\decode.id_ex_pc_reg[19] ),
    .Y(_10692_));
 sky130_fd_sc_hd__inv_2 _14650_ (.A(\decode.id_ex_pc_reg[24] ),
    .Y(_10693_));
 sky130_fd_sc_hd__buf_1 _14651_ (.A(\decode.id_ex_pc_reg[12] ),
    .X(_10694_));
 sky130_fd_sc_hd__and2_2 _14652_ (.A(_10694_),
    .B(\execute.io_target_pc[12] ),
    .X(_10695_));
 sky130_fd_sc_hd__nor2_2 _14653_ (.A(_10694_),
    .B(\execute.io_target_pc[12] ),
    .Y(_10696_));
 sky130_fd_sc_hd__buf_1 _14654_ (.A(\decode.id_ex_pc_reg[29] ),
    .X(_10697_));
 sky130_fd_sc_hd__inv_2 _14655_ (.A(\execute.io_target_pc[29] ),
    .Y(_10698_));
 sky130_fd_sc_hd__a2bb2o_2 _14656_ (.A1_N(_10695_),
    .A2_N(_10696_),
    .B1(_10697_),
    .B2(_10698_),
    .X(_10699_));
 sky130_fd_sc_hd__a221oi_2 _14657_ (.A1(_10692_),
    .A2(\execute.io_target_pc[19] ),
    .B1(_10693_),
    .B2(\execute.io_target_pc[24] ),
    .C1(_10699_),
    .Y(_10700_));
 sky130_fd_sc_hd__o211a_2 _14658_ (.A1(\decode.id_ex_pc_reg[27] ),
    .A2(_10687_),
    .B1(_10691_),
    .C1(_10700_),
    .X(_10701_));
 sky130_fd_sc_hd__inv_2 _14659_ (.A(\decode.id_ex_pc_reg[14] ),
    .Y(_10702_));
 sky130_fd_sc_hd__inv_2 _14660_ (.A(\execute.io_target_pc[0] ),
    .Y(_10703_));
 sky130_fd_sc_hd__buf_1 _14661_ (.A(\decode.id_ex_pc_reg[5] ),
    .X(_10704_));
 sky130_fd_sc_hd__inv_2 _14662_ (.A(_10704_),
    .Y(_10705_));
 sky130_fd_sc_hd__buf_1 _14663_ (.A(\decode.id_ex_pc_reg[9] ),
    .X(_10706_));
 sky130_fd_sc_hd__inv_2 _14664_ (.A(_10706_),
    .Y(_10707_));
 sky130_fd_sc_hd__a22oi_2 _14665_ (.A1(_10705_),
    .A2(\execute.io_target_pc[5] ),
    .B1(_10707_),
    .B2(\execute.io_target_pc[9] ),
    .Y(_10708_));
 sky130_fd_sc_hd__inv_2 _14666_ (.A(\execute.io_target_pc[13] ),
    .Y(_10709_));
 sky130_fd_sc_hd__buf_1 _14667_ (.A(\decode.id_ex_pc_reg[13] ),
    .X(_10710_));
 sky130_fd_sc_hd__inv_2 _14668_ (.A(\decode.id_ex_pc_reg[2] ),
    .Y(_10711_));
 sky130_fd_sc_hd__o2bb2a_2 _14669_ (.A1_N(_10709_),
    .A2_N(_10710_),
    .B1(\execute.io_target_pc[2] ),
    .B2(_10711_),
    .X(_10712_));
 sky130_fd_sc_hd__inv_2 _14670_ (.A(\decode.id_ex_pc_reg[18] ),
    .Y(_10713_));
 sky130_fd_sc_hd__o2bb2a_2 _14671_ (.A1_N(_10687_),
    .A2_N(\decode.id_ex_pc_reg[27] ),
    .B1(\execute.io_target_pc[18] ),
    .B2(_10713_),
    .X(_10714_));
 sky130_fd_sc_hd__o2111ai_2 _14672_ (.A1(\decode.id_ex_pc_reg[0] ),
    .A2(_10703_),
    .B1(_10708_),
    .C1(_10712_),
    .D1(_10714_),
    .Y(_10715_));
 sky130_fd_sc_hd__inv_2 _14673_ (.A(\decode.id_ex_pc_reg[20] ),
    .Y(_10716_));
 sky130_fd_sc_hd__inv_2 _14674_ (.A(\execute.io_target_pc[21] ),
    .Y(_10717_));
 sky130_fd_sc_hd__a22o_2 _14675_ (.A1(_10690_),
    .A2(\execute.io_target_pc[4] ),
    .B1(\decode.id_ex_pc_reg[21] ),
    .B2(_10717_),
    .X(_10718_));
 sky130_fd_sc_hd__a221o_2 _14676_ (.A1(_10703_),
    .A2(\decode.id_ex_pc_reg[0] ),
    .B1(_10716_),
    .B2(\execute.io_target_pc[20] ),
    .C1(_10718_),
    .X(_10719_));
 sky130_fd_sc_hd__inv_2 _14677_ (.A(\decode.id_ex_pc_reg[26] ),
    .Y(_10720_));
 sky130_fd_sc_hd__inv_2 _14678_ (.A(\decode.id_ex_pc_reg[10] ),
    .Y(_10721_));
 sky130_fd_sc_hd__a22oi_2 _14679_ (.A1(_10721_),
    .A2(\execute.io_target_pc[10] ),
    .B1(_10720_),
    .B2(\execute.io_target_pc[26] ),
    .Y(_10722_));
 sky130_fd_sc_hd__or2_2 _14680_ (.A(\execute.io_target_pc[30] ),
    .B(_10684_),
    .X(_10723_));
 sky130_fd_sc_hd__o211a_2 _14681_ (.A1(_10720_),
    .A2(\execute.io_target_pc[26] ),
    .B1(_10722_),
    .C1(_10723_),
    .X(_10724_));
 sky130_fd_sc_hd__inv_2 _14682_ (.A(\decode.id_ex_pc_reg[25] ),
    .Y(_10725_));
 sky130_fd_sc_hd__o2bb2a_2 _14683_ (.A1_N(_10725_),
    .A2_N(\execute.io_target_pc[25] ),
    .B1(_10721_),
    .B2(\execute.io_target_pc[10] ),
    .X(_10726_));
 sky130_fd_sc_hd__o221a_2 _14684_ (.A1(_10707_),
    .A2(\execute.io_target_pc[9] ),
    .B1(_10725_),
    .B2(\execute.io_target_pc[25] ),
    .C1(_10726_),
    .X(_10727_));
 sky130_fd_sc_hd__or2b_2 _14685_ (.A(_10678_),
    .B_N(\execute.io_target_pc[6] ),
    .X(_10728_));
 sky130_fd_sc_hd__o221a_2 _14686_ (.A1(\execute.io_target_pc[15] ),
    .A2(_10682_),
    .B1(\execute.io_target_pc[14] ),
    .B2(_10702_),
    .C1(_10728_),
    .X(_10729_));
 sky130_fd_sc_hd__buf_1 _14687_ (.A(\decode.id_ex_pc_reg[7] ),
    .X(_10730_));
 sky130_fd_sc_hd__inv_2 _14688_ (.A(_10730_),
    .Y(_10731_));
 sky130_fd_sc_hd__inv_2 _14689_ (.A(\decode.id_ex_pc_reg[23] ),
    .Y(_10732_));
 sky130_fd_sc_hd__inv_2 _14690_ (.A(\decode.id_ex_pc_reg[31] ),
    .Y(_10733_));
 sky130_fd_sc_hd__a22oi_2 _14691_ (.A1(_10732_),
    .A2(\execute.io_target_pc[23] ),
    .B1(_10733_),
    .B2(\execute.io_target_pc[31] ),
    .Y(_10734_));
 sky130_fd_sc_hd__o221a_2 _14692_ (.A1(_10731_),
    .A2(\execute.io_target_pc[7] ),
    .B1(\decode.id_ex_pc_reg[21] ),
    .B2(_10717_),
    .C1(_10734_),
    .X(_10735_));
 sky130_fd_sc_hd__inv_2 _14693_ (.A(\decode.id_ex_pc_reg[17] ),
    .Y(_10736_));
 sky130_fd_sc_hd__o2bb2a_2 _14694_ (.A1_N(\execute.io_target_pc[17] ),
    .A2_N(_10736_),
    .B1(_10688_),
    .B2(_10689_),
    .X(_10737_));
 sky130_fd_sc_hd__o221a_2 _14695_ (.A1(_10674_),
    .A2(\decode.id_ex_pc_reg[1] ),
    .B1(_10710_),
    .B2(_10709_),
    .C1(_10737_),
    .X(_10738_));
 sky130_fd_sc_hd__o2111a_2 _14696_ (.A1(_10675_),
    .A2(\execute.io_target_pc[16] ),
    .B1(_10729_),
    .C1(_10735_),
    .D1(_10738_),
    .X(_10739_));
 sky130_fd_sc_hd__nand4b_2 _14697_ (.A_N(_10719_),
    .B(_10724_),
    .C(_10727_),
    .D(_10739_),
    .Y(_10740_));
 sky130_fd_sc_hd__nand2_2 _14698_ (.A(_10731_),
    .B(\execute.io_target_pc[7] ),
    .Y(_10741_));
 sky130_fd_sc_hd__o22a_2 _14699_ (.A1(\execute.io_target_pc[20] ),
    .A2(_10716_),
    .B1(\execute.io_target_pc[17] ),
    .B2(_10736_),
    .X(_10742_));
 sky130_fd_sc_hd__inv_2 _14700_ (.A(\decode.id_ex_pc_reg[28] ),
    .Y(_10743_));
 sky130_fd_sc_hd__o22a_2 _14701_ (.A1(\decode.id_ex_pc_reg[29] ),
    .A2(_10698_),
    .B1(_10732_),
    .B2(\execute.io_target_pc[23] ),
    .X(_10744_));
 sky130_fd_sc_hd__o221a_2 _14702_ (.A1(_10705_),
    .A2(\execute.io_target_pc[5] ),
    .B1(_10692_),
    .B2(\execute.io_target_pc[19] ),
    .C1(_10744_),
    .X(_10745_));
 sky130_fd_sc_hd__a22o_2 _14703_ (.A1(_10711_),
    .A2(\execute.io_target_pc[2] ),
    .B1(_10743_),
    .B2(\execute.io_target_pc[28] ),
    .X(_10746_));
 sky130_fd_sc_hd__buf_1 _14704_ (.A(\decode.id_ex_pc_reg[3] ),
    .X(_10747_));
 sky130_fd_sc_hd__inv_2 _14705_ (.A(_10747_),
    .Y(_10748_));
 sky130_fd_sc_hd__o22a_2 _14706_ (.A1(\execute.io_target_pc[24] ),
    .A2(_10693_),
    .B1(\execute.io_target_pc[3] ),
    .B2(_10748_),
    .X(_10749_));
 sky130_fd_sc_hd__a22oi_2 _14707_ (.A1(_10748_),
    .A2(\execute.io_target_pc[3] ),
    .B1(_10677_),
    .B2(\execute.io_target_pc[22] ),
    .Y(_10750_));
 sky130_fd_sc_hd__nand2_2 _14708_ (.A(_10713_),
    .B(\execute.io_target_pc[18] ),
    .Y(_10751_));
 sky130_fd_sc_hd__and4b_2 _14709_ (.A_N(_10746_),
    .B(_10749_),
    .C(_10750_),
    .D(_10751_),
    .X(_10752_));
 sky130_fd_sc_hd__o211a_2 _14710_ (.A1(_10743_),
    .A2(\execute.io_target_pc[28] ),
    .B1(_10745_),
    .C1(_10752_),
    .X(_10753_));
 sky130_fd_sc_hd__o2111ai_2 _14711_ (.A1(_10733_),
    .A2(\execute.io_target_pc[31] ),
    .B1(_10741_),
    .C1(_10742_),
    .D1(_10753_),
    .Y(_10754_));
 sky130_fd_sc_hd__a2111oi_2 _14712_ (.A1(_10702_),
    .A2(\execute.io_target_pc[14] ),
    .B1(_10715_),
    .C1(_10740_),
    .D1(_10754_),
    .Y(_10755_));
 sky130_fd_sc_hd__a41oi_2 _14713_ (.A1(_10676_),
    .A2(_10686_),
    .A3(_10701_),
    .A4(_10755_),
    .B1(_09900_),
    .Y(_10756_));
 sky130_fd_sc_hd__buf_1 _14714_ (.A(_10756_),
    .X(_10757_));
 sky130_fd_sc_hd__or3_2 _14715_ (.A(\csr.io_trapped ),
    .B(\csr.io_mret ),
    .C(_10757_),
    .X(_10758_));
 sky130_fd_sc_hd__buf_1 _14716_ (.A(\csr.io_mem_pc[27] ),
    .X(_10759_));
 sky130_fd_sc_hd__buf_1 _14717_ (.A(\csr.io_mem_pc[26] ),
    .X(_10760_));
 sky130_fd_sc_hd__and3_2 _14718_ (.A(\csr.io_mem_pc[5] ),
    .B(\csr.io_mem_pc[6] ),
    .C(_09928_),
    .X(_10761_));
 sky130_fd_sc_hd__and4_2 _14719_ (.A(\csr.io_mem_pc[7] ),
    .B(\csr.io_mem_pc[8] ),
    .C(\csr.io_mem_pc[9] ),
    .D(_10761_),
    .X(_10762_));
 sky130_fd_sc_hd__and4_2 _14720_ (.A(\csr.io_mem_pc[10] ),
    .B(\csr.io_mem_pc[11] ),
    .C(\csr.io_mem_pc[12] ),
    .D(_10762_),
    .X(_10763_));
 sky130_fd_sc_hd__and4_2 _14721_ (.A(\csr.io_mem_pc[13] ),
    .B(\csr.io_mem_pc[14] ),
    .C(\csr.io_mem_pc[15] ),
    .D(_10763_),
    .X(_10764_));
 sky130_fd_sc_hd__and4_2 _14722_ (.A(\csr.io_mem_pc[16] ),
    .B(\csr.io_mem_pc[17] ),
    .C(\csr.io_mem_pc[18] ),
    .D(_10764_),
    .X(_10765_));
 sky130_fd_sc_hd__and4_2 _14723_ (.A(\csr.io_mem_pc[19] ),
    .B(\csr.io_mem_pc[20] ),
    .C(\csr.io_mem_pc[21] ),
    .D(_10765_),
    .X(_10766_));
 sky130_fd_sc_hd__buf_1 _14724_ (.A(_10766_),
    .X(_10767_));
 sky130_fd_sc_hd__and3_2 _14725_ (.A(\csr.io_mem_pc[22] ),
    .B(\csr.io_mem_pc[23] ),
    .C(_10767_),
    .X(_10768_));
 sky130_fd_sc_hd__and4_2 _14726_ (.A(\csr.io_mem_pc[24] ),
    .B(\csr.io_mem_pc[25] ),
    .C(_10760_),
    .D(_10768_),
    .X(_10769_));
 sky130_fd_sc_hd__and4_2 _14727_ (.A(_10759_),
    .B(\csr.io_mem_pc[28] ),
    .C(\csr.io_mem_pc[29] ),
    .D(_10769_),
    .X(_10770_));
 sky130_fd_sc_hd__buf_1 _14728_ (.A(\csr.io_mem_pc[28] ),
    .X(_10771_));
 sky130_fd_sc_hd__buf_1 _14729_ (.A(\csr.io_mem_pc[24] ),
    .X(_10772_));
 sky130_fd_sc_hd__buf_1 _14730_ (.A(\csr.io_mem_pc[25] ),
    .X(_10773_));
 sky130_fd_sc_hd__and3_2 _14731_ (.A(\csr.io_mem_pc[26] ),
    .B(\csr.io_mem_pc[27] ),
    .C(_10768_),
    .X(_10774_));
 sky130_fd_sc_hd__and3_2 _14732_ (.A(_10772_),
    .B(_10773_),
    .C(_10774_),
    .X(_10775_));
 sky130_fd_sc_hd__a21oi_2 _14733_ (.A1(_10771_),
    .A2(_10775_),
    .B1(\csr.io_mem_pc[29] ),
    .Y(_10776_));
 sky130_fd_sc_hd__buf_1 _14734_ (.A(\csr.io_mem_pc[30] ),
    .X(_10777_));
 sky130_fd_sc_hd__nand2_2 _14735_ (.A(_10684_),
    .B(_10777_),
    .Y(_10778_));
 sky130_fd_sc_hd__or2_2 _14736_ (.A(_10777_),
    .B(_10684_),
    .X(_10779_));
 sky130_fd_sc_hd__o211a_2 _14737_ (.A1(_10697_),
    .A2(_10776_),
    .B1(_10778_),
    .C1(_10779_),
    .X(_10780_));
 sky130_fd_sc_hd__and3_2 _14738_ (.A(\csr.io_mem_pc[27] ),
    .B(\csr.io_mem_pc[28] ),
    .C(_10769_),
    .X(_10781_));
 sky130_fd_sc_hd__a21oi_2 _14739_ (.A1(_10759_),
    .A2(_10769_),
    .B1(\csr.io_mem_pc[28] ),
    .Y(_10782_));
 sky130_fd_sc_hd__o21a_2 _14740_ (.A1(_10781_),
    .A2(_10782_),
    .B1(\decode.id_ex_pc_reg[28] ),
    .X(_10783_));
 sky130_fd_sc_hd__a211oi_2 _14741_ (.A1(_10771_),
    .A2(_10775_),
    .B1(_10782_),
    .C1(\decode.id_ex_pc_reg[28] ),
    .Y(_10784_));
 sky130_fd_sc_hd__a211oi_2 _14742_ (.A1(_10697_),
    .A2(_10776_),
    .B1(_10783_),
    .C1(_10784_),
    .Y(_10785_));
 sky130_fd_sc_hd__buf_1 _14743_ (.A(\decode.id_ex_pc_reg[23] ),
    .X(_10786_));
 sky130_fd_sc_hd__buf_1 _14744_ (.A(\csr.io_mem_pc[22] ),
    .X(_10787_));
 sky130_fd_sc_hd__a21oi_2 _14745_ (.A1(_10787_),
    .A2(_10767_),
    .B1(\csr.io_mem_pc[23] ),
    .Y(_10788_));
 sky130_fd_sc_hd__or2_2 _14746_ (.A(_10768_),
    .B(_10788_),
    .X(_10789_));
 sky130_fd_sc_hd__buf_1 _14747_ (.A(\decode.id_ex_pc_reg[25] ),
    .X(_10790_));
 sky130_fd_sc_hd__a21oi_2 _14748_ (.A1(\csr.io_mem_pc[24] ),
    .A2(_10768_),
    .B1(\csr.io_mem_pc[25] ),
    .Y(_10791_));
 sky130_fd_sc_hd__and3_2 _14749_ (.A(\csr.io_mem_pc[24] ),
    .B(\csr.io_mem_pc[25] ),
    .C(_10768_),
    .X(_10792_));
 sky130_fd_sc_hd__or3_2 _14750_ (.A(_10790_),
    .B(_10791_),
    .C(_10792_),
    .X(_10793_));
 sky130_fd_sc_hd__o21ai_2 _14751_ (.A1(_10791_),
    .A2(_10792_),
    .B1(_10790_),
    .Y(_10794_));
 sky130_fd_sc_hd__buf_1 _14752_ (.A(\csr.io_mem_pc[20] ),
    .X(_10795_));
 sky130_fd_sc_hd__and3_2 _14753_ (.A(\csr.io_mem_pc[19] ),
    .B(_10795_),
    .C(_10765_),
    .X(_10796_));
 sky130_fd_sc_hd__nor2_2 _14754_ (.A(\csr.io_mem_pc[21] ),
    .B(_10796_),
    .Y(_10797_));
 sky130_fd_sc_hd__buf_1 _14755_ (.A(\decode.id_ex_pc_reg[21] ),
    .X(_10798_));
 sky130_fd_sc_hd__o21a_2 _14756_ (.A1(_10767_),
    .A2(_10797_),
    .B1(_10798_),
    .X(_10799_));
 sky130_fd_sc_hd__buf_1 _14757_ (.A(\csr.io_mem_pc[19] ),
    .X(_10800_));
 sky130_fd_sc_hd__xnor2_2 _14758_ (.A(_10800_),
    .B(_10765_),
    .Y(_10801_));
 sky130_fd_sc_hd__nand2_2 _14759_ (.A(_10801_),
    .B(\decode.id_ex_pc_reg[19] ),
    .Y(_10802_));
 sky130_fd_sc_hd__buf_1 _14760_ (.A(\csr.io_mem_pc[17] ),
    .X(_10803_));
 sky130_fd_sc_hd__nand2_2 _14761_ (.A(\csr.io_mem_pc[16] ),
    .B(_10764_),
    .Y(_10804_));
 sky130_fd_sc_hd__xor2_2 _14762_ (.A(_10803_),
    .B(_10804_),
    .X(_10805_));
 sky130_fd_sc_hd__buf_1 _14763_ (.A(\decode.id_ex_pc_reg[17] ),
    .X(_10806_));
 sky130_fd_sc_hd__buf_1 _14764_ (.A(\csr.io_mem_pc[15] ),
    .X(_10807_));
 sky130_fd_sc_hd__and3_2 _14765_ (.A(\csr.io_mem_pc[13] ),
    .B(\csr.io_mem_pc[14] ),
    .C(_10763_),
    .X(_10808_));
 sky130_fd_sc_hd__nor2_2 _14766_ (.A(_10807_),
    .B(_10808_),
    .Y(_10809_));
 sky130_fd_sc_hd__xnor2_2 _14767_ (.A(\csr.io_mem_pc[13] ),
    .B(_10763_),
    .Y(_10810_));
 sky130_fd_sc_hd__nand2_2 _14768_ (.A(_10810_),
    .B(\decode.id_ex_pc_reg[13] ),
    .Y(_10811_));
 sky130_fd_sc_hd__buf_1 _14769_ (.A(\csr.io_mem_pc[11] ),
    .X(_10812_));
 sky130_fd_sc_hd__nand2_2 _14770_ (.A(\csr.io_mem_pc[10] ),
    .B(_10762_),
    .Y(_10813_));
 sky130_fd_sc_hd__xor2_2 _14771_ (.A(_10812_),
    .B(_10813_),
    .X(_10814_));
 sky130_fd_sc_hd__and3_2 _14772_ (.A(\csr.io_mem_pc[4] ),
    .B(\csr.io_mem_pc[5] ),
    .C(_09894_),
    .X(_10815_));
 sky130_fd_sc_hd__and3_2 _14773_ (.A(\csr.io_mem_pc[6] ),
    .B(\csr.io_mem_pc[7] ),
    .C(_10815_),
    .X(_10816_));
 sky130_fd_sc_hd__buf_1 _14774_ (.A(\csr.io_mem_pc[9] ),
    .X(_10817_));
 sky130_fd_sc_hd__a21oi_2 _14775_ (.A1(\csr.io_mem_pc[8] ),
    .A2(_10816_),
    .B1(_10817_),
    .Y(_10818_));
 sky130_fd_sc_hd__nand2_2 _14776_ (.A(_10814_),
    .B(\decode.id_ex_pc_reg[11] ),
    .Y(_10819_));
 sky130_fd_sc_hd__buf_1 _14777_ (.A(\csr.io_mem_pc[6] ),
    .X(_10820_));
 sky130_fd_sc_hd__buf_1 _14778_ (.A(\csr.io_mem_pc[7] ),
    .X(_10821_));
 sky130_fd_sc_hd__a21oi_2 _14779_ (.A1(_10820_),
    .A2(_10815_),
    .B1(_10821_),
    .Y(_10822_));
 sky130_fd_sc_hd__o21ai_2 _14780_ (.A1(_10762_),
    .A2(_10818_),
    .B1(\decode.id_ex_pc_reg[9] ),
    .Y(_10823_));
 sky130_fd_sc_hd__nor3_2 _14781_ (.A(_10747_),
    .B(_09887_),
    .C(_09890_),
    .Y(_10824_));
 sky130_fd_sc_hd__nor3_2 _14782_ (.A(_10748_),
    .B(_09892_),
    .C(_09894_),
    .Y(_10825_));
 sky130_fd_sc_hd__xnor2_2 _14783_ (.A(\decode.id_ex_pc_reg[31] ),
    .B(\csr.io_mem_pc[31] ),
    .Y(_10826_));
 sky130_fd_sc_hd__a21o_2 _14784_ (.A1(_10684_),
    .A2(\csr.io_mem_pc[30] ),
    .B1(_10826_),
    .X(_10827_));
 sky130_fd_sc_hd__a21oi_2 _14785_ (.A1(\csr.io_mem_pc[2] ),
    .A2(\csr.io_mem_pc[3] ),
    .B1(\csr.io_mem_pc[4] ),
    .Y(_10828_));
 sky130_fd_sc_hd__or2_2 _14786_ (.A(_09928_),
    .B(_10828_),
    .X(_10829_));
 sky130_fd_sc_hd__and2_2 _14787_ (.A(\decode.id_ex_pc_reg[0] ),
    .B(\csr.io_mem_pc[0] ),
    .X(_10830_));
 sky130_fd_sc_hd__nor2_2 _14788_ (.A(\decode.id_ex_pc_reg[0] ),
    .B(\csr.io_mem_pc[0] ),
    .Y(_10831_));
 sky130_fd_sc_hd__nor2_2 _14789_ (.A(\decode.id_ex_pc_reg[1] ),
    .B(\csr.io_mem_pc[1] ),
    .Y(_10832_));
 sky130_fd_sc_hd__and2_2 _14790_ (.A(\decode.id_ex_pc_reg[1] ),
    .B(\csr.io_mem_pc[1] ),
    .X(_10833_));
 sky130_fd_sc_hd__buf_1 _14791_ (.A(\decode.id_ex_pc_reg[2] ),
    .X(_10834_));
 sky130_fd_sc_hd__nand2_2 _14792_ (.A(_09891_),
    .B(_10834_),
    .Y(_10835_));
 sky130_fd_sc_hd__or2_2 _14793_ (.A(\csr.io_mem_pc[2] ),
    .B(_10834_),
    .X(_10836_));
 sky130_fd_sc_hd__o211a_2 _14794_ (.A1(_10832_),
    .A2(_10833_),
    .B1(_10835_),
    .C1(_10836_),
    .X(_10837_));
 sky130_fd_sc_hd__o221ai_2 _14795_ (.A1(_10830_),
    .A2(_10831_),
    .B1(\decode.id_ex_pc_reg[4] ),
    .B2(_10829_),
    .C1(_10837_),
    .Y(_10838_));
 sky130_fd_sc_hd__a21oi_2 _14796_ (.A1(\decode.id_ex_pc_reg[4] ),
    .A2(_10829_),
    .B1(_10838_),
    .Y(_10839_));
 sky130_fd_sc_hd__o21ai_2 _14797_ (.A1(_10816_),
    .A2(_10822_),
    .B1(_10730_),
    .Y(_10840_));
 sky130_fd_sc_hd__o2111a_2 _14798_ (.A1(_10824_),
    .A2(_10825_),
    .B1(_10827_),
    .C1(_10839_),
    .D1(_10840_),
    .X(_10841_));
 sky130_fd_sc_hd__o311a_2 _14799_ (.A1(_10730_),
    .A2(_10816_),
    .A3(_10822_),
    .B1(_10823_),
    .C1(_10841_),
    .X(_10842_));
 sky130_fd_sc_hd__o311a_2 _14800_ (.A1(_10706_),
    .A2(_10762_),
    .A3(_10818_),
    .B1(_10819_),
    .C1(_10842_),
    .X(_10843_));
 sky130_fd_sc_hd__o221a_2 _14801_ (.A1(\decode.id_ex_pc_reg[13] ),
    .A2(_10810_),
    .B1(_10814_),
    .B2(_10689_),
    .C1(_10843_),
    .X(_10844_));
 sky130_fd_sc_hd__o311a_2 _14802_ (.A1(\decode.id_ex_pc_reg[15] ),
    .A2(_10764_),
    .A3(_10809_),
    .B1(_10811_),
    .C1(_10844_),
    .X(_10845_));
 sky130_fd_sc_hd__o21ai_2 _14803_ (.A1(_10764_),
    .A2(_10809_),
    .B1(_10681_),
    .Y(_10846_));
 sky130_fd_sc_hd__nand2_2 _14804_ (.A(_10805_),
    .B(_10806_),
    .Y(_10847_));
 sky130_fd_sc_hd__and3_2 _14805_ (.A(_10845_),
    .B(_10846_),
    .C(_10847_),
    .X(_10848_));
 sky130_fd_sc_hd__o221a_2 _14806_ (.A1(\decode.id_ex_pc_reg[19] ),
    .A2(_10801_),
    .B1(_10805_),
    .B2(_10806_),
    .C1(_10848_),
    .X(_10849_));
 sky130_fd_sc_hd__o311ai_2 _14807_ (.A1(\decode.id_ex_pc_reg[21] ),
    .A2(_10767_),
    .A3(_10797_),
    .B1(_10802_),
    .C1(_10849_),
    .Y(_10850_));
 sky130_fd_sc_hd__a211oi_2 _14808_ (.A1(_10786_),
    .A2(_10789_),
    .B1(_10799_),
    .C1(_10850_),
    .Y(_10851_));
 sky130_fd_sc_hd__o2111a_2 _14809_ (.A1(_10786_),
    .A2(_10789_),
    .B1(_10793_),
    .C1(_10794_),
    .D1(_10851_),
    .X(_10852_));
 sky130_fd_sc_hd__nor2_2 _14810_ (.A(\csr.io_mem_pc[27] ),
    .B(_10769_),
    .Y(_10853_));
 sky130_fd_sc_hd__buf_1 _14811_ (.A(\decode.id_ex_pc_reg[27] ),
    .X(_10854_));
 sky130_fd_sc_hd__o21ai_2 _14812_ (.A1(_10775_),
    .A2(_10853_),
    .B1(_10854_),
    .Y(_10855_));
 sky130_fd_sc_hd__a311o_2 _14813_ (.A1(_10772_),
    .A2(_10773_),
    .A3(_10774_),
    .B1(_10853_),
    .C1(\decode.id_ex_pc_reg[27] ),
    .X(_10856_));
 sky130_fd_sc_hd__and3_2 _14814_ (.A(_10852_),
    .B(_10855_),
    .C(_10856_),
    .X(_10857_));
 sky130_fd_sc_hd__nor2_2 _14815_ (.A(_10760_),
    .B(_10792_),
    .Y(_10858_));
 sky130_fd_sc_hd__a21o_2 _14816_ (.A1(_10779_),
    .A2(_10826_),
    .B1(_10697_),
    .X(_10859_));
 sky130_fd_sc_hd__nand2_2 _14817_ (.A(_10770_),
    .B(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__xnor2_2 _14818_ (.A(\csr.io_mem_pc[24] ),
    .B(_10768_),
    .Y(_10861_));
 sky130_fd_sc_hd__o21ai_2 _14819_ (.A1(_10769_),
    .A2(_10858_),
    .B1(\decode.id_ex_pc_reg[26] ),
    .Y(_10862_));
 sky130_fd_sc_hd__xnor2_2 _14820_ (.A(_10787_),
    .B(_10767_),
    .Y(_10863_));
 sky130_fd_sc_hd__buf_1 _14821_ (.A(\decode.id_ex_pc_reg[22] ),
    .X(_10864_));
 sky130_fd_sc_hd__a21oi_2 _14822_ (.A1(_10800_),
    .A2(_10765_),
    .B1(_10795_),
    .Y(_10865_));
 sky130_fd_sc_hd__or2_2 _14823_ (.A(_10796_),
    .B(_10865_),
    .X(_10866_));
 sky130_fd_sc_hd__buf_1 _14824_ (.A(\decode.id_ex_pc_reg[20] ),
    .X(_10867_));
 sky130_fd_sc_hd__buf_1 _14825_ (.A(\csr.io_mem_pc[16] ),
    .X(_10868_));
 sky130_fd_sc_hd__a31oi_2 _14826_ (.A1(_10868_),
    .A2(_10803_),
    .A3(_10764_),
    .B1(\csr.io_mem_pc[18] ),
    .Y(_10869_));
 sky130_fd_sc_hd__or2_2 _14827_ (.A(_10765_),
    .B(_10869_),
    .X(_10870_));
 sky130_fd_sc_hd__buf_1 _14828_ (.A(\csr.io_mem_pc[13] ),
    .X(_10871_));
 sky130_fd_sc_hd__buf_1 _14829_ (.A(\csr.io_mem_pc[14] ),
    .X(_10872_));
 sky130_fd_sc_hd__a41o_2 _14830_ (.A1(_10871_),
    .A2(_10872_),
    .A3(_10807_),
    .A4(_10763_),
    .B1(_10868_),
    .X(_10873_));
 sky130_fd_sc_hd__a21o_2 _14831_ (.A1(_10804_),
    .A2(_10873_),
    .B1(_10675_),
    .X(_10874_));
 sky130_fd_sc_hd__nand2_2 _14832_ (.A(_10804_),
    .B(_10873_),
    .Y(_10875_));
 sky130_fd_sc_hd__a21oi_2 _14833_ (.A1(_10871_),
    .A2(_10763_),
    .B1(_10872_),
    .Y(_10876_));
 sky130_fd_sc_hd__or2_2 _14834_ (.A(_10808_),
    .B(_10876_),
    .X(_10877_));
 sky130_fd_sc_hd__buf_1 _14835_ (.A(\csr.io_mem_pc[10] ),
    .X(_10878_));
 sky130_fd_sc_hd__a31oi_2 _14836_ (.A1(_10878_),
    .A2(_10812_),
    .A3(_10762_),
    .B1(\csr.io_mem_pc[12] ),
    .Y(_10879_));
 sky130_fd_sc_hd__or2_2 _14837_ (.A(_10763_),
    .B(_10879_),
    .X(_10880_));
 sky130_fd_sc_hd__buf_1 _14838_ (.A(\csr.io_mem_pc[8] ),
    .X(_10881_));
 sky130_fd_sc_hd__a31o_2 _14839_ (.A1(_10881_),
    .A2(_10817_),
    .A3(_10816_),
    .B1(_10878_),
    .X(_10882_));
 sky130_fd_sc_hd__a21o_2 _14840_ (.A1(_10813_),
    .A2(_10882_),
    .B1(_10721_),
    .X(_10883_));
 sky130_fd_sc_hd__nand2_2 _14841_ (.A(_10881_),
    .B(_10816_),
    .Y(_10884_));
 sky130_fd_sc_hd__a31o_2 _14842_ (.A1(_10820_),
    .A2(_10821_),
    .A3(_10815_),
    .B1(\csr.io_mem_pc[8] ),
    .X(_10885_));
 sky130_fd_sc_hd__and3_2 _14843_ (.A(_10721_),
    .B(_10813_),
    .C(_10882_),
    .X(_10886_));
 sky130_fd_sc_hd__a31o_2 _14844_ (.A1(\csr.io_mem_pc[4] ),
    .A2(_09891_),
    .A3(_09888_),
    .B1(\csr.io_mem_pc[5] ),
    .X(_10887_));
 sky130_fd_sc_hd__or3b_2 _14845_ (.A(_10705_),
    .B(_10815_),
    .C_N(_10887_),
    .X(_10888_));
 sky130_fd_sc_hd__nand2_2 _14846_ (.A(\csr.io_mem_pc[5] ),
    .B(_09928_),
    .Y(_10889_));
 sky130_fd_sc_hd__a21o_2 _14847_ (.A1(_10889_),
    .A2(_10887_),
    .B1(_10704_),
    .X(_10890_));
 sky130_fd_sc_hd__a21oi_2 _14848_ (.A1(\csr.io_mem_pc[5] ),
    .A2(_09928_),
    .B1(_10820_),
    .Y(_10891_));
 sky130_fd_sc_hd__nor3_2 _14849_ (.A(_10678_),
    .B(_10761_),
    .C(_10891_),
    .Y(_10892_));
 sky130_fd_sc_hd__o21a_2 _14850_ (.A1(_10761_),
    .A2(_10891_),
    .B1(_10678_),
    .X(_10893_));
 sky130_fd_sc_hd__a211oi_2 _14851_ (.A1(_10888_),
    .A2(_10890_),
    .B1(_10892_),
    .C1(_10893_),
    .Y(_10894_));
 sky130_fd_sc_hd__a21o_2 _14852_ (.A1(_10884_),
    .A2(_10885_),
    .B1(_10680_),
    .X(_10895_));
 sky130_fd_sc_hd__nand2_2 _14853_ (.A(_10894_),
    .B(_10895_),
    .Y(_10896_));
 sky130_fd_sc_hd__a311oi_2 _14854_ (.A1(_10680_),
    .A2(_10884_),
    .A3(_10885_),
    .B1(_10886_),
    .C1(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__o211ai_2 _14855_ (.A1(\decode.id_ex_pc_reg[12] ),
    .A2(_10880_),
    .B1(_10883_),
    .C1(_10897_),
    .Y(_10898_));
 sky130_fd_sc_hd__a221oi_2 _14856_ (.A1(\decode.id_ex_pc_reg[14] ),
    .A2(_10877_),
    .B1(_10880_),
    .B2(_10694_),
    .C1(_10898_),
    .Y(_10899_));
 sky130_fd_sc_hd__o221a_2 _14857_ (.A1(\decode.id_ex_pc_reg[16] ),
    .A2(_10875_),
    .B1(_10877_),
    .B2(\decode.id_ex_pc_reg[14] ),
    .C1(_10899_),
    .X(_10900_));
 sky130_fd_sc_hd__o211ai_2 _14858_ (.A1(\decode.id_ex_pc_reg[18] ),
    .A2(_10870_),
    .B1(_10874_),
    .C1(_10900_),
    .Y(_10901_));
 sky130_fd_sc_hd__a221oi_2 _14859_ (.A1(\decode.id_ex_pc_reg[20] ),
    .A2(_10866_),
    .B1(_10870_),
    .B2(\decode.id_ex_pc_reg[18] ),
    .C1(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__o221ai_2 _14860_ (.A1(\decode.id_ex_pc_reg[22] ),
    .A2(_10863_),
    .B1(_10866_),
    .B2(_10867_),
    .C1(_10902_),
    .Y(_10903_));
 sky130_fd_sc_hd__a221oi_2 _14861_ (.A1(\decode.id_ex_pc_reg[24] ),
    .A2(_10861_),
    .B1(_10863_),
    .B2(_10864_),
    .C1(_10903_),
    .Y(_10904_));
 sky130_fd_sc_hd__o211a_2 _14862_ (.A1(\decode.id_ex_pc_reg[24] ),
    .A2(_10861_),
    .B1(_10862_),
    .C1(_10904_),
    .X(_10905_));
 sky130_fd_sc_hd__o311a_2 _14863_ (.A1(\decode.id_ex_pc_reg[26] ),
    .A2(_10769_),
    .A3(_10858_),
    .B1(_10860_),
    .C1(_10905_),
    .X(_10906_));
 sky130_fd_sc_hd__o2111a_2 _14864_ (.A1(_10770_),
    .A2(_10780_),
    .B1(_10785_),
    .C1(_10857_),
    .D1(_10906_),
    .X(_10907_));
 sky130_fd_sc_hd__nor2_2 _14865_ (.A(\fetch.bht.bhtTable_tag_MPORT_en ),
    .B(_10907_),
    .Y(_10908_));
 sky130_fd_sc_hd__or2_2 _14866_ (.A(_10758_),
    .B(_10908_),
    .X(_10909_));
 sky130_fd_sc_hd__buf_1 _14867_ (.A(_10909_),
    .X(_10910_));
 sky130_fd_sc_hd__buf_1 _14868_ (.A(_10910_),
    .X(_10911_));
 sky130_fd_sc_hd__nor4_2 _14869_ (.A(_10577_),
    .B(_10587_),
    .C(_10673_),
    .D(_10911_),
    .Y(_00342_));
 sky130_fd_sc_hd__buf_1 _14870_ (.A(_10575_),
    .X(_10912_));
 sky130_fd_sc_hd__buf_1 _14871_ (.A(_10909_),
    .X(_10913_));
 sky130_fd_sc_hd__or2b_2 _14872_ (.A(_10670_),
    .B_N(\decode.id_ex_memread_reg ),
    .X(_10914_));
 sky130_fd_sc_hd__buf_1 _14873_ (.A(_10914_),
    .X(_10915_));
 sky130_fd_sc_hd__buf_1 _14874_ (.A(_10915_),
    .X(_10916_));
 sky130_fd_sc_hd__and4bb_2 _14875_ (.A_N(_10912_),
    .B_N(_10913_),
    .C(_10916_),
    .D(\decode.immGen._imm_T_10[0] ),
    .X(_10917_));
 sky130_fd_sc_hd__buf_1 _14876_ (.A(_10917_),
    .X(_00343_));
 sky130_fd_sc_hd__and4bb_2 _14877_ (.A_N(_10912_),
    .B_N(_10913_),
    .C(_10916_),
    .D(\decode.immGen._imm_T_10[1] ),
    .X(_10918_));
 sky130_fd_sc_hd__buf_1 _14878_ (.A(_10918_),
    .X(_00344_));
 sky130_fd_sc_hd__and4bb_2 _14879_ (.A_N(_10912_),
    .B_N(_10913_),
    .C(_10916_),
    .D(\decode.immGen._imm_T_10[2] ),
    .X(_10919_));
 sky130_fd_sc_hd__buf_1 _14880_ (.A(_10919_),
    .X(_00345_));
 sky130_fd_sc_hd__and4bb_2 _14881_ (.A_N(_10912_),
    .B_N(_10913_),
    .C(_10916_),
    .D(\decode.immGen._imm_T_10[3] ),
    .X(_10920_));
 sky130_fd_sc_hd__buf_1 _14882_ (.A(_10920_),
    .X(_00346_));
 sky130_fd_sc_hd__buf_1 _14883_ (.A(_10915_),
    .X(_10921_));
 sky130_fd_sc_hd__and4bb_2 _14884_ (.A_N(_10912_),
    .B_N(_10913_),
    .C(_10921_),
    .D(\decode.immGen._imm_T_10[4] ),
    .X(_10922_));
 sky130_fd_sc_hd__buf_1 _14885_ (.A(_10922_),
    .X(_00347_));
 sky130_fd_sc_hd__buf_1 _14886_ (.A(_10618_),
    .X(_10923_));
 sky130_fd_sc_hd__buf_1 _14887_ (.A(_10923_),
    .X(_10924_));
 sky130_fd_sc_hd__buf_1 _14888_ (.A(_10924_),
    .X(_10925_));
 sky130_fd_sc_hd__buf_1 _14889_ (.A(_10925_),
    .X(_10926_));
 sky130_fd_sc_hd__buf_1 _14890_ (.A(_10926_),
    .X(_10927_));
 sky130_fd_sc_hd__buf_1 _14891_ (.A(_10927_),
    .X(_10928_));
 sky130_fd_sc_hd__buf_1 _14892_ (.A(_10928_),
    .X(_10929_));
 sky130_fd_sc_hd__buf_1 _14893_ (.A(_10929_),
    .X(_10930_));
 sky130_fd_sc_hd__buf_1 _14894_ (.A(_10930_),
    .X(_10931_));
 sky130_fd_sc_hd__and4bb_2 _14895_ (.A_N(_10912_),
    .B_N(_10913_),
    .C(_10921_),
    .D(_10931_),
    .X(_10932_));
 sky130_fd_sc_hd__buf_1 _14896_ (.A(_10932_),
    .X(_00348_));
 sky130_fd_sc_hd__buf_1 _14897_ (.A(_10604_),
    .X(_10933_));
 sky130_fd_sc_hd__nor4_2 _14898_ (.A(_10933_),
    .B(_10577_),
    .C(_10673_),
    .D(_10911_),
    .Y(_00349_));
 sky130_fd_sc_hd__inv_2 _14899_ (.A(\decode.immGen._imm_T_24[17] ),
    .Y(_10934_));
 sky130_fd_sc_hd__buf_1 _14900_ (.A(_10934_),
    .X(_10935_));
 sky130_fd_sc_hd__buf_1 _14901_ (.A(_10935_),
    .X(_10936_));
 sky130_fd_sc_hd__buf_1 _14902_ (.A(_10936_),
    .X(_10937_));
 sky130_fd_sc_hd__nor4_2 _14903_ (.A(_10937_),
    .B(_10577_),
    .C(_10673_),
    .D(_10911_),
    .Y(_00350_));
 sky130_fd_sc_hd__nor4_2 _14904_ (.A(_10606_),
    .B(_10577_),
    .C(_10673_),
    .D(_10911_),
    .Y(_00351_));
 sky130_fd_sc_hd__buf_1 _14905_ (.A(_10595_),
    .X(_10938_));
 sky130_fd_sc_hd__buf_1 _14906_ (.A(_10938_),
    .X(_10939_));
 sky130_fd_sc_hd__buf_1 _14907_ (.A(_10939_),
    .X(_10940_));
 sky130_fd_sc_hd__nor4_2 _14908_ (.A(_10940_),
    .B(_10577_),
    .C(_10673_),
    .D(_10911_),
    .Y(_00352_));
 sky130_fd_sc_hd__buf_1 _14909_ (.A(\decode.control.io_funct3[0] ),
    .X(_10941_));
 sky130_fd_sc_hd__and4bb_2 _14910_ (.A_N(_10912_),
    .B_N(_10913_),
    .C(_10921_),
    .D(_10941_),
    .X(_10942_));
 sky130_fd_sc_hd__buf_1 _14911_ (.A(_10942_),
    .X(_00353_));
 sky130_fd_sc_hd__buf_1 _14912_ (.A(\decode.control.io_funct3[1] ),
    .X(_10943_));
 sky130_fd_sc_hd__buf_1 _14913_ (.A(_10943_),
    .X(_10944_));
 sky130_fd_sc_hd__and4bb_2 _14914_ (.A_N(_10912_),
    .B_N(_10913_),
    .C(_10921_),
    .D(_10944_),
    .X(_10945_));
 sky130_fd_sc_hd__buf_1 _14915_ (.A(_10945_),
    .X(_00354_));
 sky130_fd_sc_hd__buf_1 _14916_ (.A(\decode.control.io_funct3[2] ),
    .X(_10946_));
 sky130_fd_sc_hd__and4bb_2 _14917_ (.A_N(_10912_),
    .B_N(_10913_),
    .C(_10921_),
    .D(_10946_),
    .X(_10947_));
 sky130_fd_sc_hd__buf_1 _14918_ (.A(_10947_),
    .X(_00355_));
 sky130_fd_sc_hd__buf_1 _14919_ (.A(_10667_),
    .X(_10948_));
 sky130_fd_sc_hd__and4b_2 _14920_ (.A_N(\decode.control.io_opcode[4] ),
    .B(_10580_),
    .C(_10579_),
    .D(\decode.control.io_opcode[5] ),
    .X(_10949_));
 sky130_fd_sc_hd__nor2_2 _14921_ (.A(\decode.control.io_opcode[3] ),
    .B(_10585_),
    .Y(_10950_));
 sky130_fd_sc_hd__or2_2 _14922_ (.A(_10579_),
    .B(_10578_),
    .X(_10951_));
 sky130_fd_sc_hd__nor2_2 _14923_ (.A(\decode.control.io_opcode[5] ),
    .B(_10951_),
    .Y(_10952_));
 sky130_fd_sc_hd__or3_2 _14924_ (.A(_10949_),
    .B(_10950_),
    .C(_10952_),
    .X(_10953_));
 sky130_fd_sc_hd__buf_1 _14925_ (.A(_10953_),
    .X(_10954_));
 sky130_fd_sc_hd__buf_1 _14926_ (.A(_10642_),
    .X(_10955_));
 sky130_fd_sc_hd__buf_1 _14927_ (.A(_10955_),
    .X(_10956_));
 sky130_fd_sc_hd__buf_1 _14928_ (.A(_10956_),
    .X(_10957_));
 sky130_fd_sc_hd__buf_1 _14929_ (.A(_10957_),
    .X(_10958_));
 sky130_fd_sc_hd__buf_1 _14930_ (.A(_10958_),
    .X(_10959_));
 sky130_fd_sc_hd__buf_1 _14931_ (.A(_10959_),
    .X(_10960_));
 sky130_fd_sc_hd__buf_1 _14932_ (.A(_10960_),
    .X(_10961_));
 sky130_fd_sc_hd__buf_1 _14933_ (.A(_10961_),
    .X(_10962_));
 sky130_fd_sc_hd__and3b_2 _14934_ (.A_N(_10948_),
    .B(_10954_),
    .C(_10962_),
    .X(_10963_));
 sky130_fd_sc_hd__buf_1 _14935_ (.A(\decode.control.io_opcode[4] ),
    .X(_10964_));
 sky130_fd_sc_hd__buf_1 _14936_ (.A(\decode.control.io_opcode[5] ),
    .X(_10965_));
 sky130_fd_sc_hd__and4b_2 _14937_ (.A_N(_10964_),
    .B(_10665_),
    .C(\decode.immGen._imm_T_10[0] ),
    .D(_10965_),
    .X(_10966_));
 sky130_fd_sc_hd__and4_2 _14938_ (.A(\decode.control.io_opcode[2] ),
    .B(\decode.control.io_opcode[1] ),
    .C(\decode.control.io_opcode[0] ),
    .D(_10583_),
    .X(_10967_));
 sky130_fd_sc_hd__and4bb_2 _14939_ (.A_N(_10579_),
    .B_N(\decode.control.io_opcode[3] ),
    .C(\decode.control.io_opcode[4] ),
    .D(_10584_),
    .X(_10968_));
 sky130_fd_sc_hd__buf_1 _14940_ (.A(_10968_),
    .X(_10969_));
 sky130_fd_sc_hd__buf_1 _14941_ (.A(\csr.io_mret ),
    .X(_10970_));
 sky130_fd_sc_hd__or2_2 _14942_ (.A(\csr.io_trapped ),
    .B(_10970_),
    .X(_10971_));
 sky130_fd_sc_hd__or4_2 _14943_ (.A(_10971_),
    .B(_10757_),
    .C(_10672_),
    .D(_10908_),
    .X(_10972_));
 sky130_fd_sc_hd__nor2_2 _14944_ (.A(reset),
    .B(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__o41a_2 _14945_ (.A1(_10667_),
    .A2(_10967_),
    .A3(_10952_),
    .A4(_10969_),
    .B1(_10973_),
    .X(_10974_));
 sky130_fd_sc_hd__o21a_2 _14946_ (.A1(_10963_),
    .A2(_10966_),
    .B1(_10974_),
    .X(_00356_));
 sky130_fd_sc_hd__a41o_2 _14947_ (.A1(\decode.control.io_opcode[2] ),
    .A2(\decode.control.io_opcode[1] ),
    .A3(\decode.control.io_opcode[0] ),
    .A4(_10583_),
    .B1(_10952_),
    .X(_10975_));
 sky130_fd_sc_hd__buf_1 _14948_ (.A(_10633_),
    .X(_10976_));
 sky130_fd_sc_hd__buf_1 _14949_ (.A(_10976_),
    .X(_10977_));
 sky130_fd_sc_hd__buf_1 _14950_ (.A(_10977_),
    .X(_10978_));
 sky130_fd_sc_hd__buf_1 _14951_ (.A(_10978_),
    .X(_10979_));
 sky130_fd_sc_hd__buf_1 _14952_ (.A(_10979_),
    .X(_10980_));
 sky130_fd_sc_hd__buf_1 _14953_ (.A(_10980_),
    .X(_10981_));
 sky130_fd_sc_hd__a22o_2 _14954_ (.A1(\decode.immGen._imm_T_10[1] ),
    .A2(_10948_),
    .B1(_10975_),
    .B2(_10981_),
    .X(_10982_));
 sky130_fd_sc_hd__and2_2 _14955_ (.A(_10974_),
    .B(_10982_),
    .X(_10983_));
 sky130_fd_sc_hd__buf_1 _14956_ (.A(_10983_),
    .X(_00357_));
 sky130_fd_sc_hd__a22o_2 _14957_ (.A1(\decode.immGen._imm_T_10[2] ),
    .A2(_10667_),
    .B1(_10975_),
    .B2(_10657_),
    .X(_10984_));
 sky130_fd_sc_hd__and2_2 _14958_ (.A(_10974_),
    .B(_10984_),
    .X(_10985_));
 sky130_fd_sc_hd__buf_1 _14959_ (.A(_10985_),
    .X(_00358_));
 sky130_fd_sc_hd__a22o_2 _14960_ (.A1(\decode.immGen._imm_T_10[3] ),
    .A2(_10667_),
    .B1(_10975_),
    .B2(_10662_),
    .X(_10986_));
 sky130_fd_sc_hd__and2_2 _14961_ (.A(_10974_),
    .B(_10986_),
    .X(_10987_));
 sky130_fd_sc_hd__buf_1 _14962_ (.A(_10987_),
    .X(_00359_));
 sky130_fd_sc_hd__buf_1 _14963_ (.A(_10651_),
    .X(_10988_));
 sky130_fd_sc_hd__buf_1 _14964_ (.A(_10988_),
    .X(_10989_));
 sky130_fd_sc_hd__buf_1 _14965_ (.A(_10989_),
    .X(_10990_));
 sky130_fd_sc_hd__buf_1 _14966_ (.A(_10990_),
    .X(_10991_));
 sky130_fd_sc_hd__buf_1 _14967_ (.A(_10991_),
    .X(_10992_));
 sky130_fd_sc_hd__buf_1 _14968_ (.A(_10992_),
    .X(_10993_));
 sky130_fd_sc_hd__buf_1 _14969_ (.A(_10993_),
    .X(_10994_));
 sky130_fd_sc_hd__a22o_2 _14970_ (.A1(\decode.immGen._imm_T_10[4] ),
    .A2(_10667_),
    .B1(_10975_),
    .B2(_10994_),
    .X(_10995_));
 sky130_fd_sc_hd__and2_2 _14971_ (.A(_10974_),
    .B(_10995_),
    .X(_10996_));
 sky130_fd_sc_hd__buf_1 _14972_ (.A(_10996_),
    .X(_00360_));
 sky130_fd_sc_hd__buf_1 _14973_ (.A(_10967_),
    .X(_10997_));
 sky130_fd_sc_hd__buf_1 _14974_ (.A(_10973_),
    .X(_10998_));
 sky130_fd_sc_hd__buf_1 _14975_ (.A(_10998_),
    .X(_10999_));
 sky130_fd_sc_hd__o311a_2 _14976_ (.A1(_10948_),
    .A2(_10954_),
    .A3(_10997_),
    .B1(\decode.control.io_funct7[0] ),
    .C1(_10999_),
    .X(_00361_));
 sky130_fd_sc_hd__o311a_2 _14977_ (.A1(_10948_),
    .A2(_10954_),
    .A3(_10997_),
    .B1(\decode.control.io_funct7[1] ),
    .C1(_10999_),
    .X(_00362_));
 sky130_fd_sc_hd__o311a_2 _14978_ (.A1(_10948_),
    .A2(_10954_),
    .A3(_10997_),
    .B1(\decode.control.io_funct7[2] ),
    .C1(_10999_),
    .X(_00363_));
 sky130_fd_sc_hd__o311a_2 _14979_ (.A1(_10948_),
    .A2(_10954_),
    .A3(_10997_),
    .B1(\decode.control.io_funct7[3] ),
    .C1(_10999_),
    .X(_00364_));
 sky130_fd_sc_hd__o311a_2 _14980_ (.A1(_10948_),
    .A2(_10954_),
    .A3(_10997_),
    .B1(\decode.control.io_funct7[4] ),
    .C1(_10999_),
    .X(_00365_));
 sky130_fd_sc_hd__o311a_2 _14981_ (.A1(_10948_),
    .A2(_10954_),
    .A3(_10997_),
    .B1(\decode.control.io_funct7[5] ),
    .C1(_10999_),
    .X(_00366_));
 sky130_fd_sc_hd__nor2_2 _14982_ (.A(_10964_),
    .B(_10951_),
    .Y(_11000_));
 sky130_fd_sc_hd__o31a_2 _14983_ (.A1(_10950_),
    .A2(_10952_),
    .A3(_11000_),
    .B1(\decode.control.io_funct7[6] ),
    .X(_11001_));
 sky130_fd_sc_hd__nor4_2 _14984_ (.A(_10667_),
    .B(_10950_),
    .C(_10952_),
    .D(_10969_),
    .Y(_11002_));
 sky130_fd_sc_hd__a32o_2 _14985_ (.A1(_10962_),
    .A2(_10997_),
    .A3(_11002_),
    .B1(\decode.immGen._imm_T_10[0] ),
    .B2(_10949_),
    .X(_11003_));
 sky130_fd_sc_hd__o21a_2 _14986_ (.A1(_11001_),
    .A2(_11003_),
    .B1(_10974_),
    .X(_00367_));
 sky130_fd_sc_hd__buf_1 _14987_ (.A(_10998_),
    .X(_11004_));
 sky130_fd_sc_hd__a31o_2 _14988_ (.A1(\decode.control.io_opcode[3] ),
    .A2(_10583_),
    .A3(_10584_),
    .B1(_10968_),
    .X(_11005_));
 sky130_fd_sc_hd__buf_1 _14989_ (.A(_11005_),
    .X(_11006_));
 sky130_fd_sc_hd__o311a_2 _14990_ (.A1(_10948_),
    .A2(_10950_),
    .A3(_10952_),
    .B1(_10998_),
    .C1(\decode.control.io_funct7[6] ),
    .X(_11007_));
 sky130_fd_sc_hd__a31o_2 _14991_ (.A1(_10941_),
    .A2(_11004_),
    .A3(_11006_),
    .B1(_11007_),
    .X(_00368_));
 sky130_fd_sc_hd__a31o_2 _14992_ (.A1(_10944_),
    .A2(_11004_),
    .A3(_11006_),
    .B1(_11007_),
    .X(_00369_));
 sky130_fd_sc_hd__a31o_2 _14993_ (.A1(_10946_),
    .A2(_11004_),
    .A3(_11006_),
    .B1(_11007_),
    .X(_00370_));
 sky130_fd_sc_hd__a31o_2 _14994_ (.A1(_10931_),
    .A2(_11004_),
    .A3(_11006_),
    .B1(_11007_),
    .X(_00371_));
 sky130_fd_sc_hd__buf_1 _14995_ (.A(_10612_),
    .X(_11008_));
 sky130_fd_sc_hd__buf_1 _14996_ (.A(_11008_),
    .X(_11009_));
 sky130_fd_sc_hd__buf_1 _14997_ (.A(_11009_),
    .X(_11010_));
 sky130_fd_sc_hd__buf_1 _14998_ (.A(_11010_),
    .X(_11011_));
 sky130_fd_sc_hd__a31o_2 _14999_ (.A1(_11011_),
    .A2(_11004_),
    .A3(_11006_),
    .B1(_11007_),
    .X(_00372_));
 sky130_fd_sc_hd__buf_1 _15000_ (.A(_10589_),
    .X(_11012_));
 sky130_fd_sc_hd__a31o_2 _15001_ (.A1(_11012_),
    .A2(_11004_),
    .A3(_11006_),
    .B1(_11007_),
    .X(_00373_));
 sky130_fd_sc_hd__buf_1 _15002_ (.A(_10599_),
    .X(_11013_));
 sky130_fd_sc_hd__buf_1 _15003_ (.A(_11013_),
    .X(_11014_));
 sky130_fd_sc_hd__buf_1 _15004_ (.A(_11014_),
    .X(_11015_));
 sky130_fd_sc_hd__a31o_2 _15005_ (.A1(_11015_),
    .A2(_11004_),
    .A3(_11006_),
    .B1(_11007_),
    .X(_00374_));
 sky130_fd_sc_hd__buf_1 _15006_ (.A(\decode.immGen._imm_T_24[19] ),
    .X(_11016_));
 sky130_fd_sc_hd__buf_1 _15007_ (.A(_11016_),
    .X(_11017_));
 sky130_fd_sc_hd__buf_1 _15008_ (.A(_11017_),
    .X(_11018_));
 sky130_fd_sc_hd__buf_1 _15009_ (.A(_11018_),
    .X(_11019_));
 sky130_fd_sc_hd__buf_1 _15010_ (.A(_11019_),
    .X(_11020_));
 sky130_fd_sc_hd__buf_1 _15011_ (.A(_11020_),
    .X(_11021_));
 sky130_fd_sc_hd__buf_1 _15012_ (.A(_11021_),
    .X(_11022_));
 sky130_fd_sc_hd__buf_1 _15013_ (.A(_11022_),
    .X(_11023_));
 sky130_fd_sc_hd__buf_1 _15014_ (.A(_11023_),
    .X(_11024_));
 sky130_fd_sc_hd__buf_1 _15015_ (.A(_11024_),
    .X(_11025_));
 sky130_fd_sc_hd__buf_1 _15016_ (.A(_11025_),
    .X(_11026_));
 sky130_fd_sc_hd__buf_1 _15017_ (.A(_11026_),
    .X(_11027_));
 sky130_fd_sc_hd__a31o_2 _15018_ (.A1(_11027_),
    .A2(_11004_),
    .A3(_11006_),
    .B1(_11007_),
    .X(_00375_));
 sky130_fd_sc_hd__buf_1 _15019_ (.A(_10998_),
    .X(_11028_));
 sky130_fd_sc_hd__buf_1 _15020_ (.A(_10969_),
    .X(_11029_));
 sky130_fd_sc_hd__o311a_2 _15021_ (.A1(_10667_),
    .A2(_10954_),
    .A3(_10997_),
    .B1(\decode.control.io_funct7[6] ),
    .C1(_10973_),
    .X(_11030_));
 sky130_fd_sc_hd__buf_1 _15022_ (.A(_11030_),
    .X(_11031_));
 sky130_fd_sc_hd__a31o_2 _15023_ (.A1(_10962_),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00376_));
 sky130_fd_sc_hd__buf_1 _15024_ (.A(_10981_),
    .X(_11032_));
 sky130_fd_sc_hd__a31o_2 _15025_ (.A1(_11032_),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00377_));
 sky130_fd_sc_hd__a31o_2 _15026_ (.A1(_10657_),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00378_));
 sky130_fd_sc_hd__a31o_2 _15027_ (.A1(_10662_),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00379_));
 sky130_fd_sc_hd__buf_1 _15028_ (.A(_10994_),
    .X(_11033_));
 sky130_fd_sc_hd__a31o_2 _15029_ (.A1(_11033_),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00380_));
 sky130_fd_sc_hd__a31o_2 _15030_ (.A1(\decode.control.io_funct7[0] ),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00381_));
 sky130_fd_sc_hd__a31o_2 _15031_ (.A1(\decode.control.io_funct7[1] ),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00382_));
 sky130_fd_sc_hd__a31o_2 _15032_ (.A1(\decode.control.io_funct7[2] ),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00383_));
 sky130_fd_sc_hd__a31o_2 _15033_ (.A1(\decode.control.io_funct7[3] ),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00384_));
 sky130_fd_sc_hd__a31o_2 _15034_ (.A1(\decode.control.io_funct7[4] ),
    .A2(_11028_),
    .A3(_11029_),
    .B1(_11031_),
    .X(_00385_));
 sky130_fd_sc_hd__a31o_2 _15035_ (.A1(\decode.control.io_funct7[5] ),
    .A2(_10998_),
    .A3(_10969_),
    .B1(_11030_),
    .X(_00386_));
 sky130_fd_sc_hd__a21oi_2 _15036_ (.A1(_10965_),
    .A2(_10964_),
    .B1(_10951_),
    .Y(_11034_));
 sky130_fd_sc_hd__o311a_2 _15037_ (.A1(_10950_),
    .A2(_11034_),
    .A3(_10969_),
    .B1(\decode.control.io_funct7[6] ),
    .C1(_11004_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_2 _15038_ (.A(_10659_),
    .B(_10654_),
    .X(_11035_));
 sky130_fd_sc_hd__buf_1 _15039_ (.A(_11035_),
    .X(_11036_));
 sky130_fd_sc_hd__buf_1 _15040_ (.A(_11036_),
    .X(_11037_));
 sky130_fd_sc_hd__buf_1 _15041_ (.A(_11037_),
    .X(_11038_));
 sky130_fd_sc_hd__buf_1 _15042_ (.A(_11038_),
    .X(_11039_));
 sky130_fd_sc_hd__and3_2 _15043_ (.A(_10994_),
    .B(_10981_),
    .C(_11039_),
    .X(_11040_));
 sky130_fd_sc_hd__inv_2 _15044_ (.A(\decode.immGen._imm_T_24[11] ),
    .Y(_11041_));
 sky130_fd_sc_hd__buf_1 _15045_ (.A(_11041_),
    .X(_11042_));
 sky130_fd_sc_hd__buf_1 _15046_ (.A(_11042_),
    .X(_11043_));
 sky130_fd_sc_hd__buf_1 _15047_ (.A(_11043_),
    .X(_11044_));
 sky130_fd_sc_hd__buf_1 _15048_ (.A(_11044_),
    .X(_11045_));
 sky130_fd_sc_hd__buf_1 _15049_ (.A(_11045_),
    .X(_11046_));
 sky130_fd_sc_hd__buf_1 _15050_ (.A(_11046_),
    .X(_11047_));
 sky130_fd_sc_hd__buf_1 _15051_ (.A(_11047_),
    .X(_11048_));
 sky130_fd_sc_hd__buf_1 _15052_ (.A(_11048_),
    .X(_11049_));
 sky130_fd_sc_hd__buf_1 _15053_ (.A(_11049_),
    .X(_11050_));
 sky130_fd_sc_hd__nand2_2 _15054_ (.A(_10660_),
    .B(_10655_),
    .Y(_11051_));
 sky130_fd_sc_hd__buf_1 _15055_ (.A(_11051_),
    .X(_11052_));
 sky130_fd_sc_hd__buf_1 _15056_ (.A(_11052_),
    .X(_11053_));
 sky130_fd_sc_hd__buf_1 _15057_ (.A(_11053_),
    .X(_11054_));
 sky130_fd_sc_hd__inv_2 _15058_ (.A(\decode.immGen._imm_T_24[4] ),
    .Y(_11055_));
 sky130_fd_sc_hd__buf_1 _15059_ (.A(_11055_),
    .X(_11056_));
 sky130_fd_sc_hd__buf_1 _15060_ (.A(_11056_),
    .X(_11057_));
 sky130_fd_sc_hd__buf_1 _15061_ (.A(_11057_),
    .X(_11058_));
 sky130_fd_sc_hd__buf_1 _15062_ (.A(_11058_),
    .X(_11059_));
 sky130_fd_sc_hd__buf_1 _15063_ (.A(_11059_),
    .X(_11060_));
 sky130_fd_sc_hd__buf_1 _15064_ (.A(_11060_),
    .X(_11061_));
 sky130_fd_sc_hd__buf_1 _15065_ (.A(_11061_),
    .X(_11062_));
 sky130_fd_sc_hd__or4_2 _15066_ (.A(_10979_),
    .B(_11050_),
    .C(_11054_),
    .D(_11062_),
    .X(_11063_));
 sky130_fd_sc_hd__buf_1 _15067_ (.A(_11063_),
    .X(_11064_));
 sky130_fd_sc_hd__buf_1 _15068_ (.A(_10625_),
    .X(_11065_));
 sky130_fd_sc_hd__buf_1 _15069_ (.A(_11065_),
    .X(_11066_));
 sky130_fd_sc_hd__buf_1 _15070_ (.A(_11066_),
    .X(_11067_));
 sky130_fd_sc_hd__o2111a_2 _15071_ (.A1(_10961_),
    .A2(\decode.regfile.registers_28[0] ),
    .B1(_11067_),
    .C1(_11038_),
    .D1(_10994_),
    .X(_11068_));
 sky130_fd_sc_hd__nor2b_2 _15072_ (.A(_10654_),
    .B_N(_10659_),
    .Y(_11069_));
 sky130_fd_sc_hd__buf_1 _15073_ (.A(_11069_),
    .X(_11070_));
 sky130_fd_sc_hd__buf_1 _15074_ (.A(_11070_),
    .X(_11071_));
 sky130_fd_sc_hd__buf_1 _15075_ (.A(_11071_),
    .X(_11072_));
 sky130_fd_sc_hd__and3_2 _15076_ (.A(_10989_),
    .B(_11072_),
    .C(_11065_),
    .X(_11073_));
 sky130_fd_sc_hd__buf_1 _15077_ (.A(_11073_),
    .X(_11074_));
 sky130_fd_sc_hd__buf_1 _15078_ (.A(_11074_),
    .X(_11075_));
 sky130_fd_sc_hd__buf_1 _15079_ (.A(_11049_),
    .X(_11076_));
 sky130_fd_sc_hd__and3_2 _15080_ (.A(_11074_),
    .B(_11076_),
    .C(\decode.regfile.registers_24[0] ),
    .X(_11077_));
 sky130_fd_sc_hd__a31o_2 _15081_ (.A1(_10960_),
    .A2(\decode.regfile.registers_25[0] ),
    .A3(_11075_),
    .B1(_11077_),
    .X(_11078_));
 sky130_fd_sc_hd__buf_1 _15082_ (.A(_10990_),
    .X(_11079_));
 sky130_fd_sc_hd__buf_1 _15083_ (.A(_11072_),
    .X(_11080_));
 sky130_fd_sc_hd__and3_2 _15084_ (.A(_11079_),
    .B(_10979_),
    .C(_11080_),
    .X(_11081_));
 sky130_fd_sc_hd__nand2b_2 _15085_ (.A_N(\decode.immGen._imm_T_24[3] ),
    .B(_10654_),
    .Y(_11082_));
 sky130_fd_sc_hd__buf_1 _15086_ (.A(_11082_),
    .X(_11083_));
 sky130_fd_sc_hd__buf_1 _15087_ (.A(_11083_),
    .X(_11084_));
 sky130_fd_sc_hd__buf_1 _15088_ (.A(_11084_),
    .X(_11085_));
 sky130_fd_sc_hd__or4_2 _15089_ (.A(_11060_),
    .B(_11065_),
    .C(_11049_),
    .D(_11085_),
    .X(_11086_));
 sky130_fd_sc_hd__buf_1 _15090_ (.A(_11086_),
    .X(_11087_));
 sky130_fd_sc_hd__buf_1 _15091_ (.A(_11087_),
    .X(_11088_));
 sky130_fd_sc_hd__or4b_2 _15092_ (.A(_10657_),
    .B(_10977_),
    .C(_11060_),
    .D_N(_10662_),
    .X(_11089_));
 sky130_fd_sc_hd__buf_1 _15093_ (.A(_11089_),
    .X(_11090_));
 sky130_fd_sc_hd__nor2b_2 _15094_ (.A(\decode.immGen._imm_T_24[3] ),
    .B_N(\decode.immGen._imm_T_24[2] ),
    .Y(_11091_));
 sky130_fd_sc_hd__buf_1 _15095_ (.A(_11091_),
    .X(_11092_));
 sky130_fd_sc_hd__buf_1 _15096_ (.A(_11092_),
    .X(_11093_));
 sky130_fd_sc_hd__buf_1 _15097_ (.A(_10652_),
    .X(_11094_));
 sky130_fd_sc_hd__and4_2 _15098_ (.A(_11048_),
    .B(_11093_),
    .C(_11094_),
    .D(_10976_),
    .X(_11095_));
 sky130_fd_sc_hd__buf_1 _15099_ (.A(_11095_),
    .X(_11096_));
 sky130_fd_sc_hd__or3_2 _15100_ (.A(_10628_),
    .B(_11042_),
    .C(_11082_),
    .X(_11097_));
 sky130_fd_sc_hd__buf_1 _15101_ (.A(_11097_),
    .X(_11098_));
 sky130_fd_sc_hd__buf_1 _15102_ (.A(_11098_),
    .X(_11099_));
 sky130_fd_sc_hd__buf_1 _15103_ (.A(_11099_),
    .X(_11100_));
 sky130_fd_sc_hd__and4_2 _15104_ (.A(_10625_),
    .B(_11092_),
    .C(_11048_),
    .D(_10652_),
    .X(_11101_));
 sky130_fd_sc_hd__buf_1 _15105_ (.A(_11101_),
    .X(_11102_));
 sky130_fd_sc_hd__buf_1 _15106_ (.A(_11102_),
    .X(_11103_));
 sky130_fd_sc_hd__nand2_2 _15107_ (.A(_10650_),
    .B(_10632_),
    .Y(_11104_));
 sky130_fd_sc_hd__or4_2 _15108_ (.A(_10660_),
    .B(_10655_),
    .C(_10640_),
    .D(_11104_),
    .X(_11105_));
 sky130_fd_sc_hd__buf_1 _15109_ (.A(_11105_),
    .X(_11106_));
 sky130_fd_sc_hd__nor2_2 _15110_ (.A(\decode.immGen._imm_T_24[3] ),
    .B(\decode.immGen._imm_T_24[2] ),
    .Y(_11107_));
 sky130_fd_sc_hd__buf_1 _15111_ (.A(_11107_),
    .X(_11108_));
 sky130_fd_sc_hd__buf_1 _15112_ (.A(_11108_),
    .X(_11109_));
 sky130_fd_sc_hd__buf_1 _15113_ (.A(_11109_),
    .X(_11110_));
 sky130_fd_sc_hd__buf_1 _15114_ (.A(_11110_),
    .X(_11111_));
 sky130_fd_sc_hd__buf_1 _15115_ (.A(_11111_),
    .X(_11112_));
 sky130_fd_sc_hd__buf_1 _15116_ (.A(_11112_),
    .X(_11113_));
 sky130_fd_sc_hd__buf_1 _15117_ (.A(_11113_),
    .X(_11114_));
 sky130_fd_sc_hd__nor2b_2 _15118_ (.A(\decode.immGen._imm_T_24[1] ),
    .B_N(\decode.immGen._imm_T_24[11] ),
    .Y(_11115_));
 sky130_fd_sc_hd__buf_1 _15119_ (.A(_11115_),
    .X(_11116_));
 sky130_fd_sc_hd__buf_1 _15120_ (.A(_11116_),
    .X(_11117_));
 sky130_fd_sc_hd__buf_1 _15121_ (.A(_11117_),
    .X(_11118_));
 sky130_fd_sc_hd__buf_1 _15122_ (.A(_11118_),
    .X(_11119_));
 sky130_fd_sc_hd__or2_2 _15123_ (.A(_10659_),
    .B(\decode.immGen._imm_T_24[2] ),
    .X(_11120_));
 sky130_fd_sc_hd__buf_1 _15124_ (.A(_11120_),
    .X(_11121_));
 sky130_fd_sc_hd__or4_2 _15125_ (.A(_11058_),
    .B(_10631_),
    .C(_10638_),
    .D(_11121_),
    .X(_11122_));
 sky130_fd_sc_hd__buf_1 _15126_ (.A(_11122_),
    .X(_11123_));
 sky130_fd_sc_hd__buf_1 _15127_ (.A(_11123_),
    .X(_11124_));
 sky130_fd_sc_hd__buf_1 _15128_ (.A(_11121_),
    .X(_11125_));
 sky130_fd_sc_hd__or4_2 _15129_ (.A(_11058_),
    .B(_10632_),
    .C(_11047_),
    .D(_11125_),
    .X(_11126_));
 sky130_fd_sc_hd__buf_1 _15130_ (.A(_11126_),
    .X(_11127_));
 sky130_fd_sc_hd__buf_1 _15131_ (.A(_11127_),
    .X(_11128_));
 sky130_fd_sc_hd__buf_1 _15132_ (.A(_10645_),
    .X(_11129_));
 sky130_fd_sc_hd__or4b_2 _15133_ (.A(_11129_),
    .B(_10654_),
    .C(_10623_),
    .D_N(_10659_),
    .X(_11130_));
 sky130_fd_sc_hd__buf_1 _15134_ (.A(_11130_),
    .X(_11131_));
 sky130_fd_sc_hd__buf_1 _15135_ (.A(_11131_),
    .X(_11132_));
 sky130_fd_sc_hd__and3_2 _15136_ (.A(_11069_),
    .B(_10624_),
    .C(_11058_),
    .X(_11133_));
 sky130_fd_sc_hd__buf_1 _15137_ (.A(_11133_),
    .X(_11134_));
 sky130_fd_sc_hd__or3_2 _15138_ (.A(_10645_),
    .B(_10623_),
    .C(_11082_),
    .X(_11135_));
 sky130_fd_sc_hd__buf_1 _15139_ (.A(_11135_),
    .X(_11136_));
 sky130_fd_sc_hd__buf_1 _15140_ (.A(_11055_),
    .X(_11137_));
 sky130_fd_sc_hd__and3_2 _15141_ (.A(_11091_),
    .B(_10623_),
    .C(_11137_),
    .X(_11138_));
 sky130_fd_sc_hd__buf_1 _15142_ (.A(_11138_),
    .X(_11139_));
 sky130_fd_sc_hd__and3_2 _15143_ (.A(_11055_),
    .B(_10627_),
    .C(\decode.immGen._imm_T_24[11] ),
    .X(_11140_));
 sky130_fd_sc_hd__buf_1 _15144_ (.A(_11140_),
    .X(_11141_));
 sky130_fd_sc_hd__buf_1 _15145_ (.A(_11141_),
    .X(_11142_));
 sky130_fd_sc_hd__nor2_2 _15146_ (.A(\decode.immGen._imm_T_24[4] ),
    .B(\decode.immGen._imm_T_24[1] ),
    .Y(_11143_));
 sky130_fd_sc_hd__and3_2 _15147_ (.A(_11091_),
    .B(_11041_),
    .C(_11143_),
    .X(_11144_));
 sky130_fd_sc_hd__buf_1 _15148_ (.A(_11144_),
    .X(_11145_));
 sky130_fd_sc_hd__buf_1 _15149_ (.A(_11145_),
    .X(_11146_));
 sky130_fd_sc_hd__nand3_2 _15150_ (.A(\decode.immGen._imm_T_24[1] ),
    .B(_11107_),
    .C(_11041_),
    .Y(_11147_));
 sky130_fd_sc_hd__buf_1 _15151_ (.A(_11147_),
    .X(_11148_));
 sky130_fd_sc_hd__buf_1 _15152_ (.A(_11148_),
    .X(_11149_));
 sky130_fd_sc_hd__nand3b_2 _15153_ (.A_N(_10645_),
    .B(\decode.immGen._imm_T_24[1] ),
    .C(\decode.immGen._imm_T_24[11] ),
    .Y(_11150_));
 sky130_fd_sc_hd__or3_2 _15154_ (.A(_10659_),
    .B(_10654_),
    .C(_11150_),
    .X(_11151_));
 sky130_fd_sc_hd__buf_1 _15155_ (.A(_11151_),
    .X(_11152_));
 sky130_fd_sc_hd__nand4_2 _15156_ (.A(_11107_),
    .B(_10623_),
    .C(_11055_),
    .D(\decode.immGen._imm_T_24[11] ),
    .Y(_11153_));
 sky130_fd_sc_hd__buf_1 _15157_ (.A(_11153_),
    .X(_11154_));
 sky130_fd_sc_hd__and4_2 _15158_ (.A(\decode.immGen._imm_T_24[1] ),
    .B(_11107_),
    .C(_11041_),
    .D(_11055_),
    .X(_11155_));
 sky130_fd_sc_hd__buf_1 _15159_ (.A(_11155_),
    .X(_11156_));
 sky130_fd_sc_hd__buf_1 _15160_ (.A(_11108_),
    .X(_11157_));
 sky130_fd_sc_hd__and4_2 _15161_ (.A(\decode.regfile.registers_1[0] ),
    .B(_11116_),
    .C(_11137_),
    .D(_11157_),
    .X(_11158_));
 sky130_fd_sc_hd__a211o_2 _15162_ (.A1(_11154_),
    .A2(\decode.regfile.registers_0[0] ),
    .B1(_11156_),
    .C1(_11158_),
    .X(_11159_));
 sky130_fd_sc_hd__o311a_2 _15163_ (.A1(\decode.regfile.registers_2[0] ),
    .A2(_10647_),
    .A3(_11149_),
    .B1(_11152_),
    .C1(_11159_),
    .X(_11160_));
 sky130_fd_sc_hd__a311o_2 _15164_ (.A1(\decode.regfile.registers_3[0] ),
    .A2(_11111_),
    .A3(_11142_),
    .B1(_11146_),
    .C1(_11160_),
    .X(_11161_));
 sky130_fd_sc_hd__a2111o_2 _15165_ (.A1(_11044_),
    .A2(\decode.regfile.registers_4[0] ),
    .B1(_10648_),
    .C1(_10630_),
    .D1(_11084_),
    .X(_11162_));
 sky130_fd_sc_hd__a32o_2 _15166_ (.A1(\decode.regfile.registers_5[0] ),
    .A2(_10638_),
    .A3(_11139_),
    .B1(_11161_),
    .B2(_11162_),
    .X(_11163_));
 sky130_fd_sc_hd__and3_2 _15167_ (.A(_11069_),
    .B(_11041_),
    .C(_11143_),
    .X(_11164_));
 sky130_fd_sc_hd__buf_1 _15168_ (.A(_11164_),
    .X(_11165_));
 sky130_fd_sc_hd__buf_1 _15169_ (.A(_11165_),
    .X(_11166_));
 sky130_fd_sc_hd__buf_1 _15170_ (.A(_11142_),
    .X(_11167_));
 sky130_fd_sc_hd__and4_2 _15171_ (.A(_10627_),
    .B(_11091_),
    .C(_11041_),
    .D(_11137_),
    .X(_11168_));
 sky130_fd_sc_hd__buf_1 _15172_ (.A(_11168_),
    .X(_11169_));
 sky130_fd_sc_hd__buf_1 _15173_ (.A(_11169_),
    .X(_11170_));
 sky130_fd_sc_hd__a32o_2 _15174_ (.A1(\decode.regfile.registers_7[0] ),
    .A2(_11092_),
    .A3(_11167_),
    .B1(_11170_),
    .B2(\decode.regfile.registers_6[0] ),
    .X(_11171_));
 sky130_fd_sc_hd__a211o_2 _15175_ (.A1(_11136_),
    .A2(_11163_),
    .B1(_11166_),
    .C1(_11171_),
    .X(_11172_));
 sky130_fd_sc_hd__or4b_2 _15176_ (.A(_10645_),
    .B(_10654_),
    .C(_10627_),
    .D_N(_10659_),
    .X(_11173_));
 sky130_fd_sc_hd__buf_1 _15177_ (.A(_11173_),
    .X(_11174_));
 sky130_fd_sc_hd__buf_1 _15178_ (.A(_11174_),
    .X(_11175_));
 sky130_fd_sc_hd__a21o_2 _15179_ (.A1(\decode.regfile.registers_8[0] ),
    .A2(_11046_),
    .B1(_11175_),
    .X(_11176_));
 sky130_fd_sc_hd__a32o_2 _15180_ (.A1(\decode.regfile.registers_9[0] ),
    .A2(_10639_),
    .A3(_11134_),
    .B1(_11172_),
    .B2(_11176_),
    .X(_11177_));
 sky130_fd_sc_hd__buf_1 _15181_ (.A(_10635_),
    .X(_11178_));
 sky130_fd_sc_hd__and4_2 _15182_ (.A(_10629_),
    .B(_11178_),
    .C(_11069_),
    .D(_11058_),
    .X(_11179_));
 sky130_fd_sc_hd__buf_1 _15183_ (.A(_11179_),
    .X(_11180_));
 sky130_fd_sc_hd__buf_1 _15184_ (.A(_11180_),
    .X(_11181_));
 sky130_fd_sc_hd__and4_2 _15185_ (.A(_10628_),
    .B(_11069_),
    .C(_11042_),
    .D(_11057_),
    .X(_11182_));
 sky130_fd_sc_hd__buf_1 _15186_ (.A(_11182_),
    .X(_11183_));
 sky130_fd_sc_hd__buf_1 _15187_ (.A(_11183_),
    .X(_11184_));
 sky130_fd_sc_hd__and3_2 _15188_ (.A(_10660_),
    .B(_10655_),
    .C(_11143_),
    .X(_11185_));
 sky130_fd_sc_hd__buf_1 _15189_ (.A(_11185_),
    .X(_11186_));
 sky130_fd_sc_hd__buf_1 _15190_ (.A(_11186_),
    .X(_11187_));
 sky130_fd_sc_hd__a221o_2 _15191_ (.A1(\decode.regfile.registers_11[0] ),
    .A2(_11181_),
    .B1(_11184_),
    .B2(\decode.regfile.registers_10[0] ),
    .C1(_11187_),
    .X(_11188_));
 sky130_fd_sc_hd__a21o_2 _15192_ (.A1(_11132_),
    .A2(_11177_),
    .B1(_11188_),
    .X(_11189_));
 sky130_fd_sc_hd__buf_1 _15193_ (.A(_11129_),
    .X(_11190_));
 sky130_fd_sc_hd__buf_1 _15194_ (.A(_11190_),
    .X(_11191_));
 sky130_fd_sc_hd__buf_1 _15195_ (.A(_11178_),
    .X(_11192_));
 sky130_fd_sc_hd__or4_2 _15196_ (.A(_11191_),
    .B(_10630_),
    .C(_11192_),
    .D(_11051_),
    .X(_11193_));
 sky130_fd_sc_hd__buf_1 _15197_ (.A(_11193_),
    .X(_11194_));
 sky130_fd_sc_hd__or4_2 _15198_ (.A(_10648_),
    .B(_10630_),
    .C(_11044_),
    .D(_11051_),
    .X(_11195_));
 sky130_fd_sc_hd__buf_1 _15199_ (.A(_11195_),
    .X(_11196_));
 sky130_fd_sc_hd__or3_2 _15200_ (.A(_11191_),
    .B(_10624_),
    .C(_11051_),
    .X(_11197_));
 sky130_fd_sc_hd__buf_1 _15201_ (.A(_11197_),
    .X(_11198_));
 sky130_fd_sc_hd__buf_1 _15202_ (.A(_11198_),
    .X(_11199_));
 sky130_fd_sc_hd__o221a_2 _15203_ (.A1(_11194_),
    .A2(\decode.regfile.registers_12[0] ),
    .B1(\decode.regfile.registers_13[0] ),
    .B2(_11196_),
    .C1(_11199_),
    .X(_11200_));
 sky130_fd_sc_hd__and4_2 _15204_ (.A(_10624_),
    .B(_11111_),
    .C(_11045_),
    .D(_10648_),
    .X(_11201_));
 sky130_fd_sc_hd__buf_1 _15205_ (.A(_11201_),
    .X(_11202_));
 sky130_fd_sc_hd__buf_1 _15206_ (.A(_11202_),
    .X(_11203_));
 sky130_fd_sc_hd__buf_1 _15207_ (.A(_11167_),
    .X(_11204_));
 sky130_fd_sc_hd__buf_1 _15208_ (.A(_11204_),
    .X(_11205_));
 sky130_fd_sc_hd__and4_2 _15209_ (.A(_10631_),
    .B(_11035_),
    .C(_11044_),
    .D(_11058_),
    .X(_11206_));
 sky130_fd_sc_hd__buf_1 _15210_ (.A(_11206_),
    .X(_11207_));
 sky130_fd_sc_hd__buf_1 _15211_ (.A(_11207_),
    .X(_11208_));
 sky130_fd_sc_hd__a32o_2 _15212_ (.A1(\decode.regfile.registers_15[0] ),
    .A2(_11036_),
    .A3(_11205_),
    .B1(_11208_),
    .B2(\decode.regfile.registers_14[0] ),
    .X(_11209_));
 sky130_fd_sc_hd__a211o_2 _15213_ (.A1(_11189_),
    .A2(_11200_),
    .B1(_11203_),
    .C1(_11209_),
    .X(_11210_));
 sky130_fd_sc_hd__o211a_2 _15214_ (.A1(_11124_),
    .A2(\decode.regfile.registers_16[0] ),
    .B1(_11128_),
    .C1(_11210_),
    .X(_11211_));
 sky130_fd_sc_hd__a41o_2 _15215_ (.A1(\decode.regfile.registers_17[0] ),
    .A2(_11094_),
    .A3(_11114_),
    .A4(_11119_),
    .B1(_11211_),
    .X(_11212_));
 sky130_fd_sc_hd__o2111a_2 _15216_ (.A1(\decode.regfile.registers_18[0] ),
    .A2(_10955_),
    .B1(_11114_),
    .C1(_10989_),
    .D1(_10977_),
    .X(_11213_));
 sky130_fd_sc_hd__a21o_2 _15217_ (.A1(_11106_),
    .A2(_11212_),
    .B1(_11213_),
    .X(_11214_));
 sky130_fd_sc_hd__buf_1 _15218_ (.A(_11125_),
    .X(_11215_));
 sky130_fd_sc_hd__buf_1 _15219_ (.A(_11104_),
    .X(_11216_));
 sky130_fd_sc_hd__buf_1 _15220_ (.A(_11216_),
    .X(_11217_));
 sky130_fd_sc_hd__or4_2 _15221_ (.A(_11058_),
    .B(_10633_),
    .C(_10642_),
    .D(_11085_),
    .X(_11218_));
 sky130_fd_sc_hd__buf_1 _15222_ (.A(_11218_),
    .X(_11219_));
 sky130_fd_sc_hd__o41a_2 _15223_ (.A1(\decode.regfile.registers_19[0] ),
    .A2(_11049_),
    .A3(_11215_),
    .A4(_11217_),
    .B1(_11219_),
    .X(_11220_));
 sky130_fd_sc_hd__and3_2 _15224_ (.A(_10988_),
    .B(_11118_),
    .C(_11093_),
    .X(_11221_));
 sky130_fd_sc_hd__buf_1 _15225_ (.A(_11221_),
    .X(_11222_));
 sky130_fd_sc_hd__buf_1 _15226_ (.A(_11222_),
    .X(_11223_));
 sky130_fd_sc_hd__a221o_2 _15227_ (.A1(\decode.regfile.registers_20[0] ),
    .A2(_11103_),
    .B1(_11214_),
    .B2(_11220_),
    .C1(_11223_),
    .X(_11224_));
 sky130_fd_sc_hd__buf_1 _15228_ (.A(_10642_),
    .X(_11225_));
 sky130_fd_sc_hd__or4_2 _15229_ (.A(_11059_),
    .B(_11065_),
    .C(_11225_),
    .D(_11085_),
    .X(_11226_));
 sky130_fd_sc_hd__buf_1 _15230_ (.A(_11226_),
    .X(_11227_));
 sky130_fd_sc_hd__buf_1 _15231_ (.A(_11227_),
    .X(_11228_));
 sky130_fd_sc_hd__buf_1 _15232_ (.A(_11228_),
    .X(_11229_));
 sky130_fd_sc_hd__o311a_2 _15233_ (.A1(\decode.regfile.registers_21[0] ),
    .A2(_11061_),
    .A3(_11100_),
    .B1(_11224_),
    .C1(_11229_),
    .X(_11230_));
 sky130_fd_sc_hd__and4_2 _15234_ (.A(_10989_),
    .B(_10976_),
    .C(_10955_),
    .D(_11093_),
    .X(_11231_));
 sky130_fd_sc_hd__buf_1 _15235_ (.A(_11231_),
    .X(_11232_));
 sky130_fd_sc_hd__a211o_2 _15236_ (.A1(\decode.regfile.registers_22[0] ),
    .A2(_11096_),
    .B1(_11230_),
    .C1(_11232_),
    .X(_11233_));
 sky130_fd_sc_hd__o211a_2 _15237_ (.A1(_11088_),
    .A2(\decode.regfile.registers_23[0] ),
    .B1(_11090_),
    .C1(_11233_),
    .X(_11234_));
 sky130_fd_sc_hd__or4b_2 _15238_ (.A(_10657_),
    .B(_10957_),
    .C(_11217_),
    .D_N(_10662_),
    .X(_11235_));
 sky130_fd_sc_hd__buf_1 _15239_ (.A(_11235_),
    .X(_11236_));
 sky130_fd_sc_hd__or4b_2 _15240_ (.A(_10657_),
    .B(_11049_),
    .C(_11217_),
    .D_N(_10662_),
    .X(_11237_));
 sky130_fd_sc_hd__or4_2 _15241_ (.A(_10979_),
    .B(_10958_),
    .C(_11054_),
    .D(_11062_),
    .X(_11238_));
 sky130_fd_sc_hd__o221a_2 _15242_ (.A1(\decode.regfile.registers_26[0] ),
    .A2(_11236_),
    .B1(_11237_),
    .B2(\decode.regfile.registers_27[0] ),
    .C1(_11238_),
    .X(_11239_));
 sky130_fd_sc_hd__o31a_2 _15243_ (.A1(_11078_),
    .A2(_11081_),
    .A3(_11234_),
    .B1(_11239_),
    .X(_11240_));
 sky130_fd_sc_hd__o22a_2 _15244_ (.A1(_11064_),
    .A2(\decode.regfile.registers_29[0] ),
    .B1(_11068_),
    .B2(_11240_),
    .X(_11241_));
 sky130_fd_sc_hd__or4_2 _15245_ (.A(_11062_),
    .B(_11066_),
    .C(_11076_),
    .D(_11054_),
    .X(_11242_));
 sky130_fd_sc_hd__buf_1 _15246_ (.A(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__buf_1 _15247_ (.A(_11065_),
    .X(_11244_));
 sky130_fd_sc_hd__or4_2 _15248_ (.A(_10958_),
    .B(_11054_),
    .C(_11062_),
    .D(_11244_),
    .X(_11245_));
 sky130_fd_sc_hd__buf_1 _15249_ (.A(_11245_),
    .X(_11246_));
 sky130_fd_sc_hd__o22a_2 _15250_ (.A1(\decode.regfile.registers_31[0] ),
    .A2(_11243_),
    .B1(_11246_),
    .B2(\decode.regfile.registers_30[0] ),
    .X(_11247_));
 sky130_fd_sc_hd__o41a_2 _15251_ (.A1(_10994_),
    .A2(_10981_),
    .A3(_10960_),
    .A4(_11215_),
    .B1(_10973_),
    .X(_11248_));
 sky130_fd_sc_hd__buf_1 _15252_ (.A(_11248_),
    .X(_11249_));
 sky130_fd_sc_hd__o211a_2 _15253_ (.A1(_11040_),
    .A2(_11241_),
    .B1(_11247_),
    .C1(_11249_),
    .X(_00388_));
 sky130_fd_sc_hd__buf_1 _15254_ (.A(_11050_),
    .X(_11250_));
 sky130_fd_sc_hd__buf_1 _15255_ (.A(_11250_),
    .X(_11251_));
 sky130_fd_sc_hd__or3_2 _15256_ (.A(_11062_),
    .B(_11066_),
    .C(_11054_),
    .X(_11252_));
 sky130_fd_sc_hd__buf_1 _15257_ (.A(_11252_),
    .X(_11253_));
 sky130_fd_sc_hd__nor2_2 _15258_ (.A(_10962_),
    .B(\decode.regfile.registers_30[1] ),
    .Y(_11254_));
 sky130_fd_sc_hd__buf_1 _15259_ (.A(_11063_),
    .X(_11255_));
 sky130_fd_sc_hd__o2111a_2 _15260_ (.A1(_10960_),
    .A2(\decode.regfile.registers_28[1] ),
    .B1(_11067_),
    .C1(_11038_),
    .D1(_10994_),
    .X(_11256_));
 sky130_fd_sc_hd__or4b_2 _15261_ (.A(_10657_),
    .B(_11065_),
    .C(_11061_),
    .D_N(_10662_),
    .X(_11257_));
 sky130_fd_sc_hd__buf_1 _15262_ (.A(_11257_),
    .X(_11258_));
 sky130_fd_sc_hd__buf_1 _15263_ (.A(_11258_),
    .X(_11259_));
 sky130_fd_sc_hd__buf_1 _15264_ (.A(_11235_),
    .X(_11260_));
 sky130_fd_sc_hd__buf_1 _15265_ (.A(_11072_),
    .X(_11261_));
 sky130_fd_sc_hd__buf_1 _15266_ (.A(_11086_),
    .X(_11262_));
 sky130_fd_sc_hd__buf_1 _15267_ (.A(_10956_),
    .X(_11263_));
 sky130_fd_sc_hd__buf_1 _15268_ (.A(_10977_),
    .X(_11264_));
 sky130_fd_sc_hd__buf_1 _15269_ (.A(_10989_),
    .X(_11265_));
 sky130_fd_sc_hd__o2111a_2 _15270_ (.A1(_11263_),
    .A2(\decode.regfile.registers_22[1] ),
    .B1(_11093_),
    .C1(_11264_),
    .D1(_11265_),
    .X(_11266_));
 sky130_fd_sc_hd__buf_1 _15271_ (.A(_11060_),
    .X(_11267_));
 sky130_fd_sc_hd__and4_2 _15272_ (.A(_11047_),
    .B(_11111_),
    .C(_10651_),
    .D(_10633_),
    .X(_11268_));
 sky130_fd_sc_hd__buf_1 _15273_ (.A(_11268_),
    .X(_11269_));
 sky130_fd_sc_hd__and4_2 _15274_ (.A(_10651_),
    .B(_10633_),
    .C(_10640_),
    .D(_11111_),
    .X(_11270_));
 sky130_fd_sc_hd__buf_1 _15275_ (.A(_11270_),
    .X(_11271_));
 sky130_fd_sc_hd__and3_2 _15276_ (.A(_10660_),
    .B(_10655_),
    .C(_11167_),
    .X(_11272_));
 sky130_fd_sc_hd__buf_1 _15277_ (.A(_11272_),
    .X(_11273_));
 sky130_fd_sc_hd__buf_1 _15278_ (.A(_11273_),
    .X(_11274_));
 sky130_fd_sc_hd__and3_2 _15279_ (.A(_10637_),
    .B(_11143_),
    .C(_11035_),
    .X(_11275_));
 sky130_fd_sc_hd__buf_1 _15280_ (.A(_11275_),
    .X(_11276_));
 sky130_fd_sc_hd__and3_2 _15281_ (.A(_11035_),
    .B(_11043_),
    .C(_11143_),
    .X(_11277_));
 sky130_fd_sc_hd__buf_1 _15282_ (.A(_11277_),
    .X(_11278_));
 sky130_fd_sc_hd__a22oi_2 _15283_ (.A1(\decode.regfile.registers_13[1] ),
    .A2(_11276_),
    .B1(_11278_),
    .B2(\decode.regfile.registers_12[1] ),
    .Y(_11279_));
 sky130_fd_sc_hd__buf_1 _15284_ (.A(_11192_),
    .X(_11280_));
 sky130_fd_sc_hd__buf_1 _15285_ (.A(_11133_),
    .X(_11281_));
 sky130_fd_sc_hd__a31o_2 _15286_ (.A1(\decode.regfile.registers_9[1] ),
    .A2(_11280_),
    .A3(_11281_),
    .B1(_11183_),
    .X(_11282_));
 sky130_fd_sc_hd__or4b_2 _15287_ (.A(_10645_),
    .B(_10627_),
    .C(_10635_),
    .D_N(_11069_),
    .X(_11283_));
 sky130_fd_sc_hd__buf_1 _15288_ (.A(_11283_),
    .X(_11284_));
 sky130_fd_sc_hd__buf_1 _15289_ (.A(_11284_),
    .X(_11285_));
 sky130_fd_sc_hd__or4b_2 _15290_ (.A(_11129_),
    .B(_10627_),
    .C(_11042_),
    .D_N(_11069_),
    .X(_11286_));
 sky130_fd_sc_hd__buf_1 _15291_ (.A(_11286_),
    .X(_11287_));
 sky130_fd_sc_hd__and3_2 _15292_ (.A(_11091_),
    .B(_11057_),
    .C(_10628_),
    .X(_11288_));
 sky130_fd_sc_hd__buf_1 _15293_ (.A(_11288_),
    .X(_11289_));
 sky130_fd_sc_hd__and3_2 _15294_ (.A(_11116_),
    .B(_11091_),
    .C(_11137_),
    .X(_11290_));
 sky130_fd_sc_hd__buf_1 _15295_ (.A(_11290_),
    .X(_11291_));
 sky130_fd_sc_hd__and4_2 _15296_ (.A(_10627_),
    .B(\decode.immGen._imm_T_24[11] ),
    .C(_11108_),
    .D(_11056_),
    .X(_11292_));
 sky130_fd_sc_hd__or4b_2 _15297_ (.A(_10645_),
    .B(\decode.immGen._imm_T_24[3] ),
    .C(\decode.immGen._imm_T_24[1] ),
    .D_N(\decode.immGen._imm_T_24[2] ),
    .X(_11293_));
 sky130_fd_sc_hd__o2bb2a_2 _15298_ (.A1_N(\decode.regfile.registers_3[1] ),
    .A2_N(_11292_),
    .B1(_11293_),
    .B2(_10635_),
    .X(_11294_));
 sky130_fd_sc_hd__nand4_2 _15299_ (.A(_10627_),
    .B(_11107_),
    .C(_11041_),
    .D(_11055_),
    .Y(_11295_));
 sky130_fd_sc_hd__buf_1 _15300_ (.A(_11295_),
    .X(_11296_));
 sky130_fd_sc_hd__buf_1 _15301_ (.A(_11150_),
    .X(_11297_));
 sky130_fd_sc_hd__buf_1 _15302_ (.A(_11147_),
    .X(_11298_));
 sky130_fd_sc_hd__nand4_2 _15303_ (.A(\decode.regfile.registers_1[1] ),
    .B(_11116_),
    .C(_11137_),
    .D(_11157_),
    .Y(_11299_));
 sky130_fd_sc_hd__buf_1 _15304_ (.A(_11153_),
    .X(_11300_));
 sky130_fd_sc_hd__nand2_2 _15305_ (.A(_11300_),
    .B(\decode.regfile.registers_0[1] ),
    .Y(_11301_));
 sky130_fd_sc_hd__o211ai_2 _15306_ (.A1(_11298_),
    .A2(_10646_),
    .B1(_11299_),
    .C1(_11301_),
    .Y(_11302_));
 sky130_fd_sc_hd__o221ai_2 _15307_ (.A1(\decode.regfile.registers_2[1] ),
    .A2(_11296_),
    .B1(_11297_),
    .B2(_11121_),
    .C1(_11302_),
    .Y(_11303_));
 sky130_fd_sc_hd__nand2_2 _15308_ (.A(_11294_),
    .B(_11303_),
    .Y(_11304_));
 sky130_fd_sc_hd__a2111o_2 _15309_ (.A1(_11043_),
    .A2(\decode.regfile.registers_4[1] ),
    .B1(_11190_),
    .C1(_10628_),
    .D1(_11083_),
    .X(_11305_));
 sky130_fd_sc_hd__a22oi_2 _15310_ (.A1(\decode.regfile.registers_5[1] ),
    .A2(_11291_),
    .B1(_11304_),
    .B2(_11305_),
    .Y(_11306_));
 sky130_fd_sc_hd__and4_2 _15311_ (.A(_10627_),
    .B(\decode.immGen._imm_T_24[11] ),
    .C(_11091_),
    .D(_11056_),
    .X(_11307_));
 sky130_fd_sc_hd__buf_1 _15312_ (.A(_11307_),
    .X(_11308_));
 sky130_fd_sc_hd__a221oi_2 _15313_ (.A1(\decode.regfile.registers_7[1] ),
    .A2(_11308_),
    .B1(_11169_),
    .B2(\decode.regfile.registers_6[1] ),
    .C1(_11165_),
    .Y(_11309_));
 sky130_fd_sc_hd__o21ai_2 _15314_ (.A1(_11289_),
    .A2(_11306_),
    .B1(_11309_),
    .Y(_11310_));
 sky130_fd_sc_hd__o211a_2 _15315_ (.A1(\decode.regfile.registers_8[1] ),
    .A2(_11285_),
    .B1(_11287_),
    .C1(_11310_),
    .X(_11311_));
 sky130_fd_sc_hd__o32a_2 _15316_ (.A1(\decode.regfile.registers_10[1] ),
    .A2(_10638_),
    .A3(_11132_),
    .B1(_11282_),
    .B2(_11311_),
    .X(_11312_));
 sky130_fd_sc_hd__buf_1 _15317_ (.A(_11042_),
    .X(_11313_));
 sky130_fd_sc_hd__nand2_2 _15318_ (.A(_11057_),
    .B(_10628_),
    .Y(_11314_));
 sky130_fd_sc_hd__or4b_2 _15319_ (.A(_10655_),
    .B(_11313_),
    .C(_11314_),
    .D_N(_10660_),
    .X(_11315_));
 sky130_fd_sc_hd__o32a_2 _15320_ (.A1(_10649_),
    .A2(_10631_),
    .A3(_11052_),
    .B1(\decode.regfile.registers_11[1] ),
    .B2(_11315_),
    .X(_11316_));
 sky130_fd_sc_hd__o21ai_2 _15321_ (.A1(_11181_),
    .A2(_11312_),
    .B1(_11316_),
    .Y(_11317_));
 sky130_fd_sc_hd__buf_1 _15322_ (.A(_11314_),
    .X(_11318_));
 sky130_fd_sc_hd__o2bb2a_2 _15323_ (.A1_N(_11279_),
    .A2_N(_11317_),
    .B1(_11318_),
    .B2(_11053_),
    .X(_11319_));
 sky130_fd_sc_hd__a221o_2 _15324_ (.A1(\decode.regfile.registers_14[1] ),
    .A2(_11208_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[1] ),
    .C1(_11319_),
    .X(_11320_));
 sky130_fd_sc_hd__a32o_2 _15325_ (.A1(_10651_),
    .A2(_11111_),
    .A3(_11118_),
    .B1(_11202_),
    .B2(\decode.regfile.registers_16[1] ),
    .X(_11321_));
 sky130_fd_sc_hd__a21o_2 _15326_ (.A1(_11124_),
    .A2(_11320_),
    .B1(_11321_),
    .X(_11322_));
 sky130_fd_sc_hd__o221a_2 _15327_ (.A1(_11059_),
    .A2(_11149_),
    .B1(_11127_),
    .B2(\decode.regfile.registers_17[1] ),
    .C1(_11322_),
    .X(_11323_));
 sky130_fd_sc_hd__a211o_2 _15328_ (.A1(\decode.regfile.registers_18[1] ),
    .A2(_11269_),
    .B1(_11271_),
    .C1(_11323_),
    .X(_11324_));
 sky130_fd_sc_hd__buf_1 _15329_ (.A(_11218_),
    .X(_11325_));
 sky130_fd_sc_hd__o41a_2 _15330_ (.A1(\decode.regfile.registers_19[1] ),
    .A2(_11048_),
    .A3(_11215_),
    .A4(_11216_),
    .B1(_11325_),
    .X(_11326_));
 sky130_fd_sc_hd__buf_1 _15331_ (.A(_11221_),
    .X(_11327_));
 sky130_fd_sc_hd__a221o_2 _15332_ (.A1(\decode.regfile.registers_20[1] ),
    .A2(_11102_),
    .B1(_11324_),
    .B2(_11326_),
    .C1(_11327_),
    .X(_11328_));
 sky130_fd_sc_hd__o311a_2 _15333_ (.A1(\decode.regfile.registers_21[1] ),
    .A2(_11267_),
    .A3(_11099_),
    .B1(_11228_),
    .C1(_11328_),
    .X(_11329_));
 sky130_fd_sc_hd__o22a_2 _15334_ (.A1(\decode.regfile.registers_23[1] ),
    .A2(_11262_),
    .B1(_11266_),
    .B2(_11329_),
    .X(_11330_));
 sky130_fd_sc_hd__a31o_2 _15335_ (.A1(_10992_),
    .A2(_11244_),
    .A3(_11261_),
    .B1(_11330_),
    .X(_11331_));
 sky130_fd_sc_hd__or4b_2 _15336_ (.A(_11060_),
    .B(_10977_),
    .C(_11049_),
    .D_N(_11072_),
    .X(_11332_));
 sky130_fd_sc_hd__buf_1 _15337_ (.A(_11332_),
    .X(_11333_));
 sky130_fd_sc_hd__or4b_2 _15338_ (.A(_11059_),
    .B(_10977_),
    .C(_10955_),
    .D_N(_11072_),
    .X(_11334_));
 sky130_fd_sc_hd__buf_1 _15339_ (.A(_11334_),
    .X(_11335_));
 sky130_fd_sc_hd__buf_1 _15340_ (.A(_11335_),
    .X(_11336_));
 sky130_fd_sc_hd__o22a_2 _15341_ (.A1(\decode.regfile.registers_25[1] ),
    .A2(_11333_),
    .B1(_11336_),
    .B2(\decode.regfile.registers_24[1] ),
    .X(_11337_));
 sky130_fd_sc_hd__buf_1 _15342_ (.A(_10978_),
    .X(_11338_));
 sky130_fd_sc_hd__o2111a_2 _15343_ (.A1(_10958_),
    .A2(\decode.regfile.registers_26[1] ),
    .B1(_11261_),
    .C1(_11338_),
    .D1(_10992_),
    .X(_11339_));
 sky130_fd_sc_hd__a31o_2 _15344_ (.A1(_11260_),
    .A2(_11331_),
    .A3(_11337_),
    .B1(_11339_),
    .X(_11340_));
 sky130_fd_sc_hd__o311a_2 _15345_ (.A1(_11250_),
    .A2(\decode.regfile.registers_27[1] ),
    .A3(_11259_),
    .B1(_11238_),
    .C1(_11340_),
    .X(_11341_));
 sky130_fd_sc_hd__o221ai_2 _15346_ (.A1(\decode.regfile.registers_29[1] ),
    .A2(_11255_),
    .B1(_11256_),
    .B2(_11341_),
    .C1(_11246_),
    .Y(_11342_));
 sky130_fd_sc_hd__o21ai_2 _15347_ (.A1(_11253_),
    .A2(_11254_),
    .B1(_11342_),
    .Y(_11343_));
 sky130_fd_sc_hd__o311a_2 _15348_ (.A1(_11251_),
    .A2(\decode.regfile.registers_31[1] ),
    .A3(_11253_),
    .B1(_11248_),
    .C1(_11343_),
    .X(_00389_));
 sky130_fd_sc_hd__buf_1 _15349_ (.A(_11243_),
    .X(_11344_));
 sky130_fd_sc_hd__o2111a_2 _15350_ (.A1(_10962_),
    .A2(\decode.regfile.registers_30[2] ),
    .B1(_11039_),
    .C1(_11032_),
    .D1(_11033_),
    .X(_11345_));
 sky130_fd_sc_hd__buf_1 _15351_ (.A(_10961_),
    .X(_11346_));
 sky130_fd_sc_hd__buf_1 _15352_ (.A(_11079_),
    .X(_11347_));
 sky130_fd_sc_hd__buf_1 _15353_ (.A(_11338_),
    .X(_11348_));
 sky130_fd_sc_hd__buf_1 _15354_ (.A(_11080_),
    .X(_11349_));
 sky130_fd_sc_hd__and4_2 _15355_ (.A(_11079_),
    .B(_10979_),
    .C(_10958_),
    .D(_11080_),
    .X(_11350_));
 sky130_fd_sc_hd__a41o_2 _15356_ (.A1(_11347_),
    .A2(_11348_),
    .A3(\decode.regfile.registers_26[2] ),
    .A4(_11349_),
    .B1(_11350_),
    .X(_11351_));
 sky130_fd_sc_hd__and4_2 _15357_ (.A(_10990_),
    .B(_11072_),
    .C(_11065_),
    .D(_10957_),
    .X(_11352_));
 sky130_fd_sc_hd__o2111a_2 _15358_ (.A1(_10956_),
    .A2(\decode.regfile.registers_22[2] ),
    .B1(_11093_),
    .C1(_11264_),
    .D1(_10989_),
    .X(_11353_));
 sky130_fd_sc_hd__or4_2 _15359_ (.A(_10662_),
    .B(_10657_),
    .C(_11048_),
    .D(_11104_),
    .X(_11354_));
 sky130_fd_sc_hd__and3_2 _15360_ (.A(_10650_),
    .B(_11111_),
    .C(_11117_),
    .X(_11355_));
 sky130_fd_sc_hd__buf_1 _15361_ (.A(_11355_),
    .X(_11356_));
 sky130_fd_sc_hd__buf_1 _15362_ (.A(_11356_),
    .X(_11357_));
 sky130_fd_sc_hd__nand2_2 _15363_ (.A(\decode.regfile.registers_17[2] ),
    .B(_11357_),
    .Y(_11358_));
 sky130_fd_sc_hd__buf_1 _15364_ (.A(_11123_),
    .X(_11359_));
 sky130_fd_sc_hd__buf_1 _15365_ (.A(_11207_),
    .X(_11360_));
 sky130_fd_sc_hd__buf_1 _15366_ (.A(_11201_),
    .X(_11361_));
 sky130_fd_sc_hd__a221o_2 _15367_ (.A1(\decode.regfile.registers_14[2] ),
    .A2(_11360_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[2] ),
    .C1(_11361_),
    .X(_11362_));
 sky130_fd_sc_hd__a31o_2 _15368_ (.A1(\decode.regfile.registers_11[2] ),
    .A2(_11071_),
    .A3(_11204_),
    .B1(_11187_),
    .X(_11363_));
 sky130_fd_sc_hd__buf_1 _15369_ (.A(_11315_),
    .X(_11364_));
 sky130_fd_sc_hd__buf_1 _15370_ (.A(_11287_),
    .X(_11365_));
 sky130_fd_sc_hd__o22ai_2 _15371_ (.A1(\decode.regfile.registers_8[2] ),
    .A2(_11285_),
    .B1(_11365_),
    .B2(\decode.regfile.registers_9[2] ),
    .Y(_11366_));
 sky130_fd_sc_hd__buf_1 _15372_ (.A(_11293_),
    .X(_11367_));
 sky130_fd_sc_hd__o2bb2a_2 _15373_ (.A1_N(\decode.regfile.registers_3[2] ),
    .A2_N(_11292_),
    .B1(_11367_),
    .B2(_11178_),
    .X(_11368_));
 sky130_fd_sc_hd__buf_1 _15374_ (.A(_11295_),
    .X(_11369_));
 sky130_fd_sc_hd__a31oi_2 _15375_ (.A1(_11117_),
    .A2(_11137_),
    .A3(_11157_),
    .B1(\decode.regfile.registers_0[2] ),
    .Y(_11370_));
 sky130_fd_sc_hd__buf_1 _15376_ (.A(_11153_),
    .X(_11371_));
 sky130_fd_sc_hd__nor2_2 _15377_ (.A(\decode.regfile.registers_1[2] ),
    .B(_11371_),
    .Y(_11372_));
 sky130_fd_sc_hd__o21ai_2 _15378_ (.A1(_11370_),
    .A2(_11372_),
    .B1(_11296_),
    .Y(_11373_));
 sky130_fd_sc_hd__o221ai_2 _15379_ (.A1(\decode.regfile.registers_2[2] ),
    .A2(_11369_),
    .B1(_11297_),
    .B2(_11121_),
    .C1(_11373_),
    .Y(_11374_));
 sky130_fd_sc_hd__or4_2 _15380_ (.A(_10645_),
    .B(_10627_),
    .C(\decode.immGen._imm_T_24[11] ),
    .D(_11082_),
    .X(_11375_));
 sky130_fd_sc_hd__o2bb2a_2 _15381_ (.A1_N(_11368_),
    .A2_N(_11374_),
    .B1(_11375_),
    .B2(\decode.regfile.registers_4[2] ),
    .X(_11376_));
 sky130_fd_sc_hd__mux2_2 _15382_ (.A0(_11376_),
    .A1(\decode.regfile.registers_5[2] ),
    .S(_11291_),
    .X(_11377_));
 sky130_fd_sc_hd__buf_1 _15383_ (.A(_11308_),
    .X(_11378_));
 sky130_fd_sc_hd__a221o_2 _15384_ (.A1(\decode.regfile.registers_7[2] ),
    .A2(_11378_),
    .B1(_11170_),
    .B2(\decode.regfile.registers_6[2] ),
    .C1(_11281_),
    .X(_11379_));
 sky130_fd_sc_hd__a21oi_2 _15385_ (.A1(_11136_),
    .A2(_11377_),
    .B1(_11379_),
    .Y(_11380_));
 sky130_fd_sc_hd__or4b_2 _15386_ (.A(_10655_),
    .B(_10636_),
    .C(_11314_),
    .D_N(_10660_),
    .X(_11381_));
 sky130_fd_sc_hd__buf_1 _15387_ (.A(_11381_),
    .X(_11382_));
 sky130_fd_sc_hd__o21ai_2 _15388_ (.A1(_11366_),
    .A2(_11380_),
    .B1(_11382_),
    .Y(_11383_));
 sky130_fd_sc_hd__o311a_2 _15389_ (.A1(\decode.regfile.registers_10[2] ),
    .A2(_10639_),
    .A3(_11132_),
    .B1(_11364_),
    .C1(_11383_),
    .X(_11384_));
 sky130_fd_sc_hd__o22a_2 _15390_ (.A1(_11194_),
    .A2(\decode.regfile.registers_12[2] ),
    .B1(\decode.regfile.registers_13[2] ),
    .B2(_11196_),
    .X(_11385_));
 sky130_fd_sc_hd__o211a_2 _15391_ (.A1(_11363_),
    .A2(_11384_),
    .B1(_11385_),
    .C1(_11199_),
    .X(_11386_));
 sky130_fd_sc_hd__o221ai_2 _15392_ (.A1(\decode.regfile.registers_16[2] ),
    .A2(_11359_),
    .B1(_11362_),
    .B2(_11386_),
    .C1(_11126_),
    .Y(_11387_));
 sky130_fd_sc_hd__a21oi_2 _15393_ (.A1(_11358_),
    .A2(_11387_),
    .B1(_11268_),
    .Y(_11388_));
 sky130_fd_sc_hd__a211o_2 _15394_ (.A1(\decode.regfile.registers_18[2] ),
    .A2(_11268_),
    .B1(_11271_),
    .C1(_11388_),
    .X(_11389_));
 sky130_fd_sc_hd__o211a_2 _15395_ (.A1(\decode.regfile.registers_19[2] ),
    .A2(_11354_),
    .B1(_11218_),
    .C1(_11389_),
    .X(_11390_));
 sky130_fd_sc_hd__a211o_2 _15396_ (.A1(\decode.regfile.registers_20[2] ),
    .A2(_11102_),
    .B1(_11327_),
    .C1(_11390_),
    .X(_11391_));
 sky130_fd_sc_hd__o311a_2 _15397_ (.A1(\decode.regfile.registers_21[2] ),
    .A2(_11060_),
    .A3(_11098_),
    .B1(_11227_),
    .C1(_11391_),
    .X(_11392_));
 sky130_fd_sc_hd__o221a_2 _15398_ (.A1(\decode.regfile.registers_23[2] ),
    .A2(_11086_),
    .B1(_11353_),
    .B2(_11392_),
    .C1(_11335_),
    .X(_11393_));
 sky130_fd_sc_hd__a211o_2 _15399_ (.A1(\decode.regfile.registers_24[2] ),
    .A2(_11074_),
    .B1(_11352_),
    .C1(_11393_),
    .X(_11394_));
 sky130_fd_sc_hd__o311a_2 _15400_ (.A1(_11076_),
    .A2(\decode.regfile.registers_25[2] ),
    .A3(_11090_),
    .B1(_11235_),
    .C1(_11394_),
    .X(_11395_));
 sky130_fd_sc_hd__buf_1 _15401_ (.A(_11238_),
    .X(_11396_));
 sky130_fd_sc_hd__o221ai_2 _15402_ (.A1(\decode.regfile.registers_27[2] ),
    .A2(_11237_),
    .B1(_11351_),
    .B2(_11395_),
    .C1(_11396_),
    .Y(_11397_));
 sky130_fd_sc_hd__and3_2 _15403_ (.A(_11347_),
    .B(_11037_),
    .C(_11066_),
    .X(_11398_));
 sky130_fd_sc_hd__o21ai_2 _15404_ (.A1(_10960_),
    .A2(\decode.regfile.registers_28[2] ),
    .B1(_11398_),
    .Y(_11399_));
 sky130_fd_sc_hd__nand2_2 _15405_ (.A(_11397_),
    .B(_11399_),
    .Y(_11400_));
 sky130_fd_sc_hd__o221a_2 _15406_ (.A1(_11346_),
    .A2(_11253_),
    .B1(_11064_),
    .B2(\decode.regfile.registers_29[2] ),
    .C1(_11400_),
    .X(_11401_));
 sky130_fd_sc_hd__o221a_2 _15407_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[2] ),
    .B1(_11345_),
    .B2(_11401_),
    .C1(_11249_),
    .X(_00390_));
 sky130_fd_sc_hd__o2111a_2 _15408_ (.A1(_10962_),
    .A2(\decode.regfile.registers_30[3] ),
    .B1(_11039_),
    .C1(_11032_),
    .D1(_11033_),
    .X(_11402_));
 sky130_fd_sc_hd__buf_1 _15409_ (.A(_11238_),
    .X(_11403_));
 sky130_fd_sc_hd__buf_1 _15410_ (.A(_11093_),
    .X(_11404_));
 sky130_fd_sc_hd__o2111a_2 _15411_ (.A1(_10957_),
    .A2(\decode.regfile.registers_22[3] ),
    .B1(_11404_),
    .C1(_10978_),
    .D1(_10990_),
    .X(_11405_));
 sky130_fd_sc_hd__buf_1 _15412_ (.A(_11354_),
    .X(_11406_));
 sky130_fd_sc_hd__buf_1 _15413_ (.A(_11278_),
    .X(_11407_));
 sky130_fd_sc_hd__a221o_2 _15414_ (.A1(\decode.regfile.registers_7[3] ),
    .A2(_11378_),
    .B1(_11170_),
    .B2(\decode.regfile.registers_6[3] ),
    .C1(_11134_),
    .X(_11408_));
 sky130_fd_sc_hd__and3_2 _15415_ (.A(\decode.regfile.registers_5[3] ),
    .B(_10637_),
    .C(_11139_),
    .X(_11409_));
 sky130_fd_sc_hd__buf_1 _15416_ (.A(_11367_),
    .X(_11410_));
 sky130_fd_sc_hd__and4_2 _15417_ (.A(\decode.regfile.registers_1[3] ),
    .B(_11116_),
    .C(_11137_),
    .D(_11157_),
    .X(_11411_));
 sky130_fd_sc_hd__a211o_2 _15418_ (.A1(_11154_),
    .A2(\decode.regfile.registers_0[3] ),
    .B1(_11156_),
    .C1(_11411_),
    .X(_11412_));
 sky130_fd_sc_hd__or3_2 _15419_ (.A(\decode.regfile.registers_2[3] ),
    .B(_10646_),
    .C(_11298_),
    .X(_11413_));
 sky130_fd_sc_hd__a31o_2 _15420_ (.A1(\decode.regfile.registers_3[3] ),
    .A2(_11109_),
    .A3(_11141_),
    .B1(_11145_),
    .X(_11414_));
 sky130_fd_sc_hd__a31o_2 _15421_ (.A1(_11152_),
    .A2(_11412_),
    .A3(_11413_),
    .B1(_11414_),
    .X(_11415_));
 sky130_fd_sc_hd__o221a_2 _15422_ (.A1(\decode.regfile.registers_4[3] ),
    .A2(_11410_),
    .B1(_11097_),
    .B2(_10648_),
    .C1(_11415_),
    .X(_11416_));
 sky130_fd_sc_hd__o32a_2 _15423_ (.A1(_10648_),
    .A2(_10624_),
    .A3(_11085_),
    .B1(_11409_),
    .B2(_11416_),
    .X(_11417_));
 sky130_fd_sc_hd__o221a_2 _15424_ (.A1(\decode.regfile.registers_8[3] ),
    .A2(_11285_),
    .B1(_11365_),
    .B2(\decode.regfile.registers_9[3] ),
    .C1(_11132_),
    .X(_11418_));
 sky130_fd_sc_hd__o21ai_2 _15425_ (.A1(_11408_),
    .A2(_11417_),
    .B1(_11418_),
    .Y(_11419_));
 sky130_fd_sc_hd__a22oi_2 _15426_ (.A1(\decode.regfile.registers_11[3] ),
    .A2(_11181_),
    .B1(_11184_),
    .B2(\decode.regfile.registers_10[3] ),
    .Y(_11420_));
 sky130_fd_sc_hd__a21oi_2 _15427_ (.A1(_11419_),
    .A2(_11420_),
    .B1(_11186_),
    .Y(_11421_));
 sky130_fd_sc_hd__a221o_2 _15428_ (.A1(\decode.regfile.registers_13[3] ),
    .A2(_11276_),
    .B1(_11407_),
    .B2(\decode.regfile.registers_12[3] ),
    .C1(_11421_),
    .X(_11422_));
 sky130_fd_sc_hd__a31o_2 _15429_ (.A1(\decode.regfile.registers_15[3] ),
    .A2(_11036_),
    .A3(_11204_),
    .B1(_11361_),
    .X(_11423_));
 sky130_fd_sc_hd__a221o_2 _15430_ (.A1(\decode.regfile.registers_14[3] ),
    .A2(_11208_),
    .B1(_11422_),
    .B2(_11199_),
    .C1(_11423_),
    .X(_11424_));
 sky130_fd_sc_hd__o211a_2 _15431_ (.A1(_11124_),
    .A2(\decode.regfile.registers_16[3] ),
    .B1(_11127_),
    .C1(_11424_),
    .X(_11425_));
 sky130_fd_sc_hd__a21oi_2 _15432_ (.A1(\decode.regfile.registers_17[3] ),
    .A2(_11357_),
    .B1(_11425_),
    .Y(_11426_));
 sky130_fd_sc_hd__a21oi_2 _15433_ (.A1(\decode.regfile.registers_18[3] ),
    .A2(_11269_),
    .B1(_11271_),
    .Y(_11427_));
 sky130_fd_sc_hd__o21ai_2 _15434_ (.A1(_11269_),
    .A2(_11426_),
    .B1(_11427_),
    .Y(_11428_));
 sky130_fd_sc_hd__o211a_2 _15435_ (.A1(\decode.regfile.registers_19[3] ),
    .A2(_11406_),
    .B1(_11325_),
    .C1(_11428_),
    .X(_11429_));
 sky130_fd_sc_hd__a211o_2 _15436_ (.A1(\decode.regfile.registers_20[3] ),
    .A2(_11103_),
    .B1(_11222_),
    .C1(_11429_),
    .X(_11430_));
 sky130_fd_sc_hd__o311a_2 _15437_ (.A1(\decode.regfile.registers_21[3] ),
    .A2(_11267_),
    .A3(_11099_),
    .B1(_11228_),
    .C1(_11430_),
    .X(_11431_));
 sky130_fd_sc_hd__o22a_2 _15438_ (.A1(\decode.regfile.registers_23[3] ),
    .A2(_11087_),
    .B1(_11405_),
    .B2(_11431_),
    .X(_11432_));
 sky130_fd_sc_hd__a31o_2 _15439_ (.A1(_10992_),
    .A2(_11066_),
    .A3(_11261_),
    .B1(_11432_),
    .X(_11433_));
 sky130_fd_sc_hd__o22a_2 _15440_ (.A1(\decode.regfile.registers_25[3] ),
    .A2(_11333_),
    .B1(_11336_),
    .B2(\decode.regfile.registers_24[3] ),
    .X(_11434_));
 sky130_fd_sc_hd__buf_1 _15441_ (.A(_10957_),
    .X(_11435_));
 sky130_fd_sc_hd__buf_1 _15442_ (.A(_11435_),
    .X(_11436_));
 sky130_fd_sc_hd__o2111a_2 _15443_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[3] ),
    .B1(_11349_),
    .C1(_10980_),
    .D1(_11347_),
    .X(_11437_));
 sky130_fd_sc_hd__a31o_2 _15444_ (.A1(_11236_),
    .A2(_11433_),
    .A3(_11434_),
    .B1(_11437_),
    .X(_11438_));
 sky130_fd_sc_hd__or3_2 _15445_ (.A(_11250_),
    .B(\decode.regfile.registers_27[3] ),
    .C(_11258_),
    .X(_11439_));
 sky130_fd_sc_hd__buf_1 _15446_ (.A(_11347_),
    .X(_11440_));
 sky130_fd_sc_hd__o2111a_2 _15447_ (.A1(_10960_),
    .A2(\decode.regfile.registers_28[3] ),
    .B1(_11067_),
    .C1(_11038_),
    .D1(_11440_),
    .X(_11441_));
 sky130_fd_sc_hd__a31o_2 _15448_ (.A1(_11403_),
    .A2(_11438_),
    .A3(_11439_),
    .B1(_11441_),
    .X(_11442_));
 sky130_fd_sc_hd__o221a_2 _15449_ (.A1(_11346_),
    .A2(_11253_),
    .B1(_11064_),
    .B2(\decode.regfile.registers_29[3] ),
    .C1(_11442_),
    .X(_11443_));
 sky130_fd_sc_hd__o221a_2 _15450_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[3] ),
    .B1(_11402_),
    .B2(_11443_),
    .C1(_11249_),
    .X(_00391_));
 sky130_fd_sc_hd__o2111a_2 _15451_ (.A1(_10962_),
    .A2(\decode.regfile.registers_30[4] ),
    .B1(_11039_),
    .C1(_11032_),
    .D1(_11033_),
    .X(_11444_));
 sky130_fd_sc_hd__buf_1 _15452_ (.A(_11398_),
    .X(_11445_));
 sky130_fd_sc_hd__buf_1 _15453_ (.A(_10959_),
    .X(_11446_));
 sky130_fd_sc_hd__buf_1 _15454_ (.A(_11349_),
    .X(_11447_));
 sky130_fd_sc_hd__buf_1 _15455_ (.A(_11347_),
    .X(_11448_));
 sky130_fd_sc_hd__o2111a_2 _15456_ (.A1(_11446_),
    .A2(\decode.regfile.registers_26[4] ),
    .B1(_11447_),
    .C1(_10981_),
    .D1(_11448_),
    .X(_11449_));
 sky130_fd_sc_hd__buf_1 _15457_ (.A(_11404_),
    .X(_11450_));
 sky130_fd_sc_hd__o2111a_2 _15458_ (.A1(_11435_),
    .A2(\decode.regfile.registers_22[4] ),
    .B1(_11450_),
    .C1(_10979_),
    .D1(_10991_),
    .X(_11451_));
 sky130_fd_sc_hd__buf_1 _15459_ (.A(_11103_),
    .X(_11452_));
 sky130_fd_sc_hd__buf_1 _15460_ (.A(_11406_),
    .X(_11453_));
 sky130_fd_sc_hd__buf_1 _15461_ (.A(_11219_),
    .X(_11454_));
 sky130_fd_sc_hd__buf_1 _15462_ (.A(_11269_),
    .X(_11455_));
 sky130_fd_sc_hd__buf_1 _15463_ (.A(_11271_),
    .X(_11456_));
 sky130_fd_sc_hd__a221o_2 _15464_ (.A1(\decode.regfile.registers_14[4] ),
    .A2(_11360_),
    .B1(_11273_),
    .B2(\decode.regfile.registers_15[4] ),
    .C1(_11361_),
    .X(_11457_));
 sky130_fd_sc_hd__and4_2 _15465_ (.A(\decode.regfile.registers_1[4] ),
    .B(_11115_),
    .C(_11056_),
    .D(_11108_),
    .X(_11458_));
 sky130_fd_sc_hd__a211o_2 _15466_ (.A1(_11300_),
    .A2(\decode.regfile.registers_0[4] ),
    .B1(_11155_),
    .C1(_11458_),
    .X(_11459_));
 sky130_fd_sc_hd__o311a_2 _15467_ (.A1(\decode.regfile.registers_2[4] ),
    .A2(_11190_),
    .A3(_11148_),
    .B1(_11151_),
    .C1(_11459_),
    .X(_11460_));
 sky130_fd_sc_hd__a311o_2 _15468_ (.A1(\decode.regfile.registers_3[4] ),
    .A2(_11110_),
    .A3(_11142_),
    .B1(_11146_),
    .C1(_11460_),
    .X(_11461_));
 sky130_fd_sc_hd__buf_1 _15469_ (.A(_11082_),
    .X(_11462_));
 sky130_fd_sc_hd__a2111o_2 _15470_ (.A1(_11313_),
    .A2(\decode.regfile.registers_4[4] ),
    .B1(_11191_),
    .C1(_10630_),
    .D1(_11462_),
    .X(_11463_));
 sky130_fd_sc_hd__a32o_2 _15471_ (.A1(\decode.regfile.registers_5[4] ),
    .A2(_10637_),
    .A3(_11139_),
    .B1(_11461_),
    .B2(_11463_),
    .X(_11464_));
 sky130_fd_sc_hd__buf_1 _15472_ (.A(_11308_),
    .X(_11465_));
 sky130_fd_sc_hd__buf_1 _15473_ (.A(_11169_),
    .X(_11466_));
 sky130_fd_sc_hd__a221o_2 _15474_ (.A1(\decode.regfile.registers_7[4] ),
    .A2(_11465_),
    .B1(_11466_),
    .B2(\decode.regfile.registers_6[4] ),
    .C1(_11281_),
    .X(_11467_));
 sky130_fd_sc_hd__a21o_2 _15475_ (.A1(_11136_),
    .A2(_11464_),
    .B1(_11467_),
    .X(_11468_));
 sky130_fd_sc_hd__o221a_2 _15476_ (.A1(\decode.regfile.registers_8[4] ),
    .A2(_11285_),
    .B1(_11365_),
    .B2(\decode.regfile.registers_9[4] ),
    .C1(_11132_),
    .X(_11469_));
 sky130_fd_sc_hd__buf_1 _15477_ (.A(_11167_),
    .X(_11470_));
 sky130_fd_sc_hd__a31o_2 _15478_ (.A1(\decode.regfile.registers_11[4] ),
    .A2(_11070_),
    .A3(_11470_),
    .B1(_11186_),
    .X(_11471_));
 sky130_fd_sc_hd__a221o_2 _15479_ (.A1(\decode.regfile.registers_10[4] ),
    .A2(_11184_),
    .B1(_11468_),
    .B2(_11469_),
    .C1(_11471_),
    .X(_11472_));
 sky130_fd_sc_hd__o221a_2 _15480_ (.A1(_11194_),
    .A2(\decode.regfile.registers_12[4] ),
    .B1(\decode.regfile.registers_13[4] ),
    .B2(_11195_),
    .C1(_11198_),
    .X(_11473_));
 sky130_fd_sc_hd__and2_2 _15481_ (.A(_11472_),
    .B(_11473_),
    .X(_11474_));
 sky130_fd_sc_hd__o221a_2 _15482_ (.A1(\decode.regfile.registers_16[4] ),
    .A2(_11359_),
    .B1(_11457_),
    .B2(_11474_),
    .C1(_11126_),
    .X(_11475_));
 sky130_fd_sc_hd__a41o_2 _15483_ (.A1(\decode.regfile.registers_17[4] ),
    .A2(_10652_),
    .A3(_11112_),
    .A4(_11118_),
    .B1(_11475_),
    .X(_11476_));
 sky130_fd_sc_hd__o31a_2 _15484_ (.A1(_10955_),
    .A2(_11215_),
    .A3(_11216_),
    .B1(_11476_),
    .X(_11477_));
 sky130_fd_sc_hd__a211o_2 _15485_ (.A1(\decode.regfile.registers_18[4] ),
    .A2(_11455_),
    .B1(_11456_),
    .C1(_11477_),
    .X(_11478_));
 sky130_fd_sc_hd__o211a_2 _15486_ (.A1(\decode.regfile.registers_19[4] ),
    .A2(_11453_),
    .B1(_11454_),
    .C1(_11478_),
    .X(_11479_));
 sky130_fd_sc_hd__a211o_2 _15487_ (.A1(\decode.regfile.registers_20[4] ),
    .A2(_11452_),
    .B1(_11223_),
    .C1(_11479_),
    .X(_11480_));
 sky130_fd_sc_hd__o311a_2 _15488_ (.A1(\decode.regfile.registers_21[4] ),
    .A2(_11062_),
    .A3(_11100_),
    .B1(_11229_),
    .C1(_11480_),
    .X(_11481_));
 sky130_fd_sc_hd__o22a_2 _15489_ (.A1(\decode.regfile.registers_23[4] ),
    .A2(_11088_),
    .B1(_11451_),
    .B2(_11481_),
    .X(_11482_));
 sky130_fd_sc_hd__buf_1 _15490_ (.A(_11333_),
    .X(_11483_));
 sky130_fd_sc_hd__buf_1 _15491_ (.A(_11335_),
    .X(_11484_));
 sky130_fd_sc_hd__o22a_2 _15492_ (.A1(\decode.regfile.registers_25[4] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[4] ),
    .X(_11485_));
 sky130_fd_sc_hd__buf_1 _15493_ (.A(_11235_),
    .X(_11486_));
 sky130_fd_sc_hd__o211a_2 _15494_ (.A1(_11075_),
    .A2(_11482_),
    .B1(_11485_),
    .C1(_11486_),
    .X(_11487_));
 sky130_fd_sc_hd__o32a_2 _15495_ (.A1(_11251_),
    .A2(_11259_),
    .A3(\decode.regfile.registers_27[4] ),
    .B1(_11449_),
    .B2(_11487_),
    .X(_11488_));
 sky130_fd_sc_hd__buf_1 _15496_ (.A(_11238_),
    .X(_11489_));
 sky130_fd_sc_hd__o221a_2 _15497_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[4] ),
    .B1(\decode.regfile.registers_29[4] ),
    .B2(_11255_),
    .C1(_11246_),
    .X(_11490_));
 sky130_fd_sc_hd__o21a_2 _15498_ (.A1(_11445_),
    .A2(_11488_),
    .B1(_11490_),
    .X(_11491_));
 sky130_fd_sc_hd__o221a_2 _15499_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[4] ),
    .B1(_11444_),
    .B2(_11491_),
    .C1(_11249_),
    .X(_00392_));
 sky130_fd_sc_hd__o2111a_2 _15500_ (.A1(_10962_),
    .A2(\decode.regfile.registers_30[5] ),
    .B1(_11039_),
    .C1(_11032_),
    .D1(_11033_),
    .X(_11492_));
 sky130_fd_sc_hd__buf_1 _15501_ (.A(_10956_),
    .X(_11493_));
 sky130_fd_sc_hd__o2111a_2 _15502_ (.A1(_11493_),
    .A2(\decode.regfile.registers_24[5] ),
    .B1(_11065_),
    .C1(_11072_),
    .D1(_10990_),
    .X(_11494_));
 sky130_fd_sc_hd__o2111a_2 _15503_ (.A1(_10956_),
    .A2(\decode.regfile.registers_22[5] ),
    .B1(_11093_),
    .C1(_10977_),
    .D1(_10989_),
    .X(_11495_));
 sky130_fd_sc_hd__a221o_2 _15504_ (.A1(\decode.regfile.registers_14[5] ),
    .A2(_11206_),
    .B1(_11272_),
    .B2(\decode.regfile.registers_15[5] ),
    .C1(_11201_),
    .X(_11496_));
 sky130_fd_sc_hd__a221o_2 _15505_ (.A1(\decode.regfile.registers_7[5] ),
    .A2(_11465_),
    .B1(_11466_),
    .B2(\decode.regfile.registers_6[5] ),
    .C1(_11281_),
    .X(_11497_));
 sky130_fd_sc_hd__and4_2 _15506_ (.A(\decode.regfile.registers_1[5] ),
    .B(_11115_),
    .C(_11056_),
    .D(_11108_),
    .X(_11498_));
 sky130_fd_sc_hd__a211o_2 _15507_ (.A1(_11371_),
    .A2(\decode.regfile.registers_0[5] ),
    .B1(_11155_),
    .C1(_11498_),
    .X(_11499_));
 sky130_fd_sc_hd__o221ai_2 _15508_ (.A1(\decode.regfile.registers_2[5] ),
    .A2(_11369_),
    .B1(_11297_),
    .B2(_11121_),
    .C1(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__o2bb2a_2 _15509_ (.A1_N(\decode.regfile.registers_3[5] ),
    .A2_N(_11292_),
    .B1(_11293_),
    .B2(_10635_),
    .X(_11501_));
 sky130_fd_sc_hd__nand2_2 _15510_ (.A(_11500_),
    .B(_11501_),
    .Y(_11502_));
 sky130_fd_sc_hd__buf_1 _15511_ (.A(_11129_),
    .X(_11503_));
 sky130_fd_sc_hd__a2111o_2 _15512_ (.A1(_11043_),
    .A2(\decode.regfile.registers_4[5] ),
    .B1(_11503_),
    .C1(_10629_),
    .D1(_11083_),
    .X(_11504_));
 sky130_fd_sc_hd__a32o_2 _15513_ (.A1(\decode.regfile.registers_5[5] ),
    .A2(_11192_),
    .A3(_11139_),
    .B1(_11502_),
    .B2(_11504_),
    .X(_11505_));
 sky130_fd_sc_hd__o31a_2 _15514_ (.A1(_10648_),
    .A2(_10624_),
    .A3(_11084_),
    .B1(_11505_),
    .X(_11506_));
 sky130_fd_sc_hd__o221a_2 _15515_ (.A1(\decode.regfile.registers_8[5] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(\decode.regfile.registers_9[5] ),
    .C1(_11131_),
    .X(_11507_));
 sky130_fd_sc_hd__o21ai_2 _15516_ (.A1(_11497_),
    .A2(_11506_),
    .B1(_11507_),
    .Y(_11508_));
 sky130_fd_sc_hd__buf_1 _15517_ (.A(_11183_),
    .X(_11509_));
 sky130_fd_sc_hd__a221oi_2 _15518_ (.A1(\decode.regfile.registers_11[5] ),
    .A2(_11180_),
    .B1(_11509_),
    .B2(\decode.regfile.registers_10[5] ),
    .C1(_11186_),
    .Y(_11510_));
 sky130_fd_sc_hd__nand2_2 _15519_ (.A(_11508_),
    .B(_11510_),
    .Y(_11511_));
 sky130_fd_sc_hd__o221a_2 _15520_ (.A1(_11193_),
    .A2(\decode.regfile.registers_12[5] ),
    .B1(\decode.regfile.registers_13[5] ),
    .B2(_11195_),
    .C1(_11198_),
    .X(_11512_));
 sky130_fd_sc_hd__and2_2 _15521_ (.A(_11511_),
    .B(_11512_),
    .X(_11513_));
 sky130_fd_sc_hd__o22a_2 _15522_ (.A1(\decode.regfile.registers_16[5] ),
    .A2(_11122_),
    .B1(_11496_),
    .B2(_11513_),
    .X(_11514_));
 sky130_fd_sc_hd__a31o_2 _15523_ (.A1(_10651_),
    .A2(_11111_),
    .A3(_11118_),
    .B1(_11514_),
    .X(_11515_));
 sky130_fd_sc_hd__o211a_2 _15524_ (.A1(_11127_),
    .A2(\decode.regfile.registers_17[5] ),
    .B1(_11105_),
    .C1(_11515_),
    .X(_11516_));
 sky130_fd_sc_hd__a211o_2 _15525_ (.A1(\decode.regfile.registers_18[5] ),
    .A2(_11268_),
    .B1(_11271_),
    .C1(_11516_),
    .X(_11517_));
 sky130_fd_sc_hd__o211a_2 _15526_ (.A1(\decode.regfile.registers_19[5] ),
    .A2(_11354_),
    .B1(_11218_),
    .C1(_11517_),
    .X(_11518_));
 sky130_fd_sc_hd__a211o_2 _15527_ (.A1(\decode.regfile.registers_20[5] ),
    .A2(_11102_),
    .B1(_11221_),
    .C1(_11518_),
    .X(_11519_));
 sky130_fd_sc_hd__o311a_2 _15528_ (.A1(\decode.regfile.registers_21[5] ),
    .A2(_11060_),
    .A3(_11098_),
    .B1(_11227_),
    .C1(_11519_),
    .X(_11520_));
 sky130_fd_sc_hd__o221a_2 _15529_ (.A1(\decode.regfile.registers_23[5] ),
    .A2(_11086_),
    .B1(_11495_),
    .B2(_11520_),
    .C1(_11335_),
    .X(_11521_));
 sky130_fd_sc_hd__o32a_2 _15530_ (.A1(_11050_),
    .A2(_11089_),
    .A3(\decode.regfile.registers_25[5] ),
    .B1(_11494_),
    .B2(_11521_),
    .X(_11522_));
 sky130_fd_sc_hd__a221o_2 _15531_ (.A1(\decode.regfile.registers_26[5] ),
    .A2(_11081_),
    .B1(_11522_),
    .B2(_11235_),
    .C1(_11350_),
    .X(_11523_));
 sky130_fd_sc_hd__or3_2 _15532_ (.A(_11250_),
    .B(\decode.regfile.registers_27[5] ),
    .C(_11258_),
    .X(_11524_));
 sky130_fd_sc_hd__o2111a_2 _15533_ (.A1(_10960_),
    .A2(\decode.regfile.registers_28[5] ),
    .B1(_11067_),
    .C1(_11038_),
    .D1(_11440_),
    .X(_11525_));
 sky130_fd_sc_hd__a31o_2 _15534_ (.A1(_11403_),
    .A2(_11523_),
    .A3(_11524_),
    .B1(_11525_),
    .X(_11526_));
 sky130_fd_sc_hd__o221a_2 _15535_ (.A1(_11346_),
    .A2(_11253_),
    .B1(_11064_),
    .B2(\decode.regfile.registers_29[5] ),
    .C1(_11526_),
    .X(_11527_));
 sky130_fd_sc_hd__o221a_2 _15536_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[5] ),
    .B1(_11492_),
    .B2(_11527_),
    .C1(_11249_),
    .X(_00393_));
 sky130_fd_sc_hd__o2111a_2 _15537_ (.A1(_10962_),
    .A2(\decode.regfile.registers_30[6] ),
    .B1(_11039_),
    .C1(_11032_),
    .D1(_11033_),
    .X(_11528_));
 sky130_fd_sc_hd__or2_2 _15538_ (.A(_11493_),
    .B(\decode.regfile.registers_24[6] ),
    .X(_11529_));
 sky130_fd_sc_hd__o2111a_2 _15539_ (.A1(_10956_),
    .A2(\decode.regfile.registers_22[6] ),
    .B1(_11093_),
    .C1(_11264_),
    .D1(_11265_),
    .X(_11530_));
 sky130_fd_sc_hd__a221o_2 _15540_ (.A1(\decode.regfile.registers_14[6] ),
    .A2(_11207_),
    .B1(_11273_),
    .B2(\decode.regfile.registers_15[6] ),
    .C1(_11201_),
    .X(_11531_));
 sky130_fd_sc_hd__a22o_2 _15541_ (.A1(\decode.regfile.registers_13[6] ),
    .A2(_11275_),
    .B1(_11278_),
    .B2(\decode.regfile.registers_12[6] ),
    .X(_11532_));
 sky130_fd_sc_hd__or4_2 _15542_ (.A(_11503_),
    .B(_10624_),
    .C(_11043_),
    .D(_11083_),
    .X(_11533_));
 sky130_fd_sc_hd__or4_2 _15543_ (.A(_10646_),
    .B(_10624_),
    .C(_10635_),
    .D(_11082_),
    .X(_11534_));
 sky130_fd_sc_hd__o221ai_2 _15544_ (.A1(\decode.regfile.registers_7[6] ),
    .A2(_11533_),
    .B1(\decode.regfile.registers_6[6] ),
    .B2(_11534_),
    .C1(_11174_),
    .Y(_11535_));
 sky130_fd_sc_hd__or3_2 _15545_ (.A(\decode.regfile.registers_5[6] ),
    .B(_11313_),
    .C(_11410_),
    .X(_11536_));
 sky130_fd_sc_hd__o2bb2a_2 _15546_ (.A1_N(\decode.regfile.registers_2[6] ),
    .A2_N(_11155_),
    .B1(_11150_),
    .B2(_11120_),
    .X(_11537_));
 sky130_fd_sc_hd__and3_2 _15547_ (.A(_11115_),
    .B(_11055_),
    .C(_11107_),
    .X(_11538_));
 sky130_fd_sc_hd__buf_1 _15548_ (.A(_11538_),
    .X(_11539_));
 sky130_fd_sc_hd__o22a_2 _15549_ (.A1(_11129_),
    .A2(_11147_),
    .B1(_11300_),
    .B2(\decode.regfile.registers_1[6] ),
    .X(_11540_));
 sky130_fd_sc_hd__o21ai_2 _15550_ (.A1(\decode.regfile.registers_0[6] ),
    .A2(_11539_),
    .B1(_11540_),
    .Y(_11541_));
 sky130_fd_sc_hd__a2bb2o_2 _15551_ (.A1_N(\decode.regfile.registers_3[6] ),
    .A2_N(_11152_),
    .B1(_11537_),
    .B2(_11541_),
    .X(_11542_));
 sky130_fd_sc_hd__o21ai_2 _15552_ (.A1(\decode.regfile.registers_4[6] ),
    .A2(_10636_),
    .B1(_11138_),
    .Y(_11543_));
 sky130_fd_sc_hd__o21ai_2 _15553_ (.A1(_11146_),
    .A2(_11542_),
    .B1(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__a21oi_2 _15554_ (.A1(_11536_),
    .A2(_11544_),
    .B1(_11289_),
    .Y(_11545_));
 sky130_fd_sc_hd__and3_2 _15555_ (.A(_10635_),
    .B(_11143_),
    .C(_11069_),
    .X(_11546_));
 sky130_fd_sc_hd__buf_1 _15556_ (.A(_11546_),
    .X(_11547_));
 sky130_fd_sc_hd__a221oi_2 _15557_ (.A1(\decode.regfile.registers_8[6] ),
    .A2(_11166_),
    .B1(_11547_),
    .B2(\decode.regfile.registers_9[6] ),
    .C1(_11183_),
    .Y(_11548_));
 sky130_fd_sc_hd__o21ai_2 _15558_ (.A1(_11535_),
    .A2(_11545_),
    .B1(_11548_),
    .Y(_11549_));
 sky130_fd_sc_hd__o31a_2 _15559_ (.A1(\decode.regfile.registers_10[6] ),
    .A2(_10637_),
    .A3(_11131_),
    .B1(_11315_),
    .X(_11550_));
 sky130_fd_sc_hd__a32o_2 _15560_ (.A1(\decode.regfile.registers_11[6] ),
    .A2(_11070_),
    .A3(_11470_),
    .B1(_11549_),
    .B2(_11550_),
    .X(_11551_));
 sky130_fd_sc_hd__o31a_2 _15561_ (.A1(_10649_),
    .A2(_10632_),
    .A3(_11052_),
    .B1(_11551_),
    .X(_11552_));
 sky130_fd_sc_hd__o32a_2 _15562_ (.A1(_10650_),
    .A2(_10625_),
    .A3(_11053_),
    .B1(_11532_),
    .B2(_11552_),
    .X(_11553_));
 sky130_fd_sc_hd__o22a_2 _15563_ (.A1(\decode.regfile.registers_16[6] ),
    .A2(_11123_),
    .B1(_11531_),
    .B2(_11553_),
    .X(_11554_));
 sky130_fd_sc_hd__mux2_2 _15564_ (.A0(_11554_),
    .A1(\decode.regfile.registers_17[6] ),
    .S(_11356_),
    .X(_11555_));
 sky130_fd_sc_hd__o2111a_2 _15565_ (.A1(\decode.regfile.registers_18[6] ),
    .A2(_10642_),
    .B1(_11112_),
    .C1(_10652_),
    .D1(_10633_),
    .X(_11556_));
 sky130_fd_sc_hd__a21o_2 _15566_ (.A1(_11106_),
    .A2(_11555_),
    .B1(_11556_),
    .X(_11557_));
 sky130_fd_sc_hd__o211a_2 _15567_ (.A1(\decode.regfile.registers_19[6] ),
    .A2(_11354_),
    .B1(_11325_),
    .C1(_11557_),
    .X(_11558_));
 sky130_fd_sc_hd__a211o_2 _15568_ (.A1(\decode.regfile.registers_20[6] ),
    .A2(_11102_),
    .B1(_11327_),
    .C1(_11558_),
    .X(_11559_));
 sky130_fd_sc_hd__o311a_2 _15569_ (.A1(\decode.regfile.registers_21[6] ),
    .A2(_11267_),
    .A3(_11098_),
    .B1(_11227_),
    .C1(_11559_),
    .X(_11560_));
 sky130_fd_sc_hd__o221a_2 _15570_ (.A1(\decode.regfile.registers_23[6] ),
    .A2(_11262_),
    .B1(_11530_),
    .B2(_11560_),
    .C1(_11335_),
    .X(_11561_));
 sky130_fd_sc_hd__a41o_2 _15571_ (.A1(_11079_),
    .A2(_11244_),
    .A3(_11261_),
    .A4(_11529_),
    .B1(_11561_),
    .X(_11562_));
 sky130_fd_sc_hd__or3_2 _15572_ (.A(_11050_),
    .B(\decode.regfile.registers_25[6] ),
    .C(_11090_),
    .X(_11563_));
 sky130_fd_sc_hd__buf_1 _15573_ (.A(_11079_),
    .X(_11564_));
 sky130_fd_sc_hd__o2111a_2 _15574_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[6] ),
    .B1(_11349_),
    .C1(_10980_),
    .D1(_11564_),
    .X(_11565_));
 sky130_fd_sc_hd__a31o_2 _15575_ (.A1(_11236_),
    .A2(_11562_),
    .A3(_11563_),
    .B1(_11565_),
    .X(_11566_));
 sky130_fd_sc_hd__or3_2 _15576_ (.A(_11250_),
    .B(\decode.regfile.registers_27[6] ),
    .C(_11258_),
    .X(_11567_));
 sky130_fd_sc_hd__o2111a_2 _15577_ (.A1(_10960_),
    .A2(\decode.regfile.registers_28[6] ),
    .B1(_11067_),
    .C1(_11038_),
    .D1(_11440_),
    .X(_11568_));
 sky130_fd_sc_hd__a31o_2 _15578_ (.A1(_11403_),
    .A2(_11566_),
    .A3(_11567_),
    .B1(_11568_),
    .X(_11569_));
 sky130_fd_sc_hd__o221a_2 _15579_ (.A1(_11346_),
    .A2(_11253_),
    .B1(_11064_),
    .B2(\decode.regfile.registers_29[6] ),
    .C1(_11569_),
    .X(_11570_));
 sky130_fd_sc_hd__o221a_2 _15580_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[6] ),
    .B1(_11528_),
    .B2(_11570_),
    .C1(_11249_),
    .X(_00394_));
 sky130_fd_sc_hd__buf_1 _15581_ (.A(_10961_),
    .X(_11571_));
 sky130_fd_sc_hd__o2111a_2 _15582_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[7] ),
    .B1(_11039_),
    .C1(_11032_),
    .D1(_11033_),
    .X(_11572_));
 sky130_fd_sc_hd__o2111a_2 _15583_ (.A1(_11263_),
    .A2(\decode.regfile.registers_22[7] ),
    .B1(_11404_),
    .C1(_10978_),
    .D1(_10990_),
    .X(_11573_));
 sky130_fd_sc_hd__a221o_2 _15584_ (.A1(\decode.regfile.registers_14[7] ),
    .A2(_11360_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[7] ),
    .C1(_11202_),
    .X(_11574_));
 sky130_fd_sc_hd__a31o_2 _15585_ (.A1(\decode.regfile.registers_9[7] ),
    .A2(_11280_),
    .A3(_11281_),
    .B1(_11183_),
    .X(_11575_));
 sky130_fd_sc_hd__a31o_2 _15586_ (.A1(\decode.regfile.registers_7[7] ),
    .A2(_11092_),
    .A3(_11142_),
    .B1(_11165_),
    .X(_11576_));
 sky130_fd_sc_hd__a31o_2 _15587_ (.A1(\decode.regfile.registers_3[7] ),
    .A2(_11157_),
    .A3(_11140_),
    .B1(_11145_),
    .X(_11577_));
 sky130_fd_sc_hd__nand4_2 _15588_ (.A(\decode.regfile.registers_1[7] ),
    .B(_11115_),
    .C(_11056_),
    .D(_11108_),
    .Y(_11578_));
 sky130_fd_sc_hd__nand2_2 _15589_ (.A(_11153_),
    .B(\decode.regfile.registers_0[7] ),
    .Y(_11579_));
 sky130_fd_sc_hd__o211ai_2 _15590_ (.A1(_11147_),
    .A2(_10645_),
    .B1(_11578_),
    .C1(_11579_),
    .Y(_11580_));
 sky130_fd_sc_hd__o311a_2 _15591_ (.A1(\decode.regfile.registers_2[7] ),
    .A2(_11129_),
    .A3(_11147_),
    .B1(_11151_),
    .C1(_11580_),
    .X(_11581_));
 sky130_fd_sc_hd__o22ai_2 _15592_ (.A1(\decode.regfile.registers_4[7] ),
    .A2(_11375_),
    .B1(_11577_),
    .B2(_11581_),
    .Y(_11582_));
 sky130_fd_sc_hd__o2bb2a_2 _15593_ (.A1_N(\decode.regfile.registers_5[7] ),
    .A2_N(_11290_),
    .B1(_10635_),
    .B2(_11135_),
    .X(_11583_));
 sky130_fd_sc_hd__o21ai_2 _15594_ (.A1(_11290_),
    .A2(_11582_),
    .B1(_11583_),
    .Y(_11584_));
 sky130_fd_sc_hd__o221a_2 _15595_ (.A1(_11084_),
    .A2(_11297_),
    .B1(_11534_),
    .B2(\decode.regfile.registers_6[7] ),
    .C1(_11584_),
    .X(_11585_));
 sky130_fd_sc_hd__a21o_2 _15596_ (.A1(\decode.regfile.registers_8[7] ),
    .A2(_11044_),
    .B1(_11174_),
    .X(_11586_));
 sky130_fd_sc_hd__o21a_2 _15597_ (.A1(_11576_),
    .A2(_11585_),
    .B1(_11586_),
    .X(_11587_));
 sky130_fd_sc_hd__o32a_2 _15598_ (.A1(\decode.regfile.registers_10[7] ),
    .A2(_10638_),
    .A3(_11132_),
    .B1(_11575_),
    .B2(_11587_),
    .X(_11588_));
 sky130_fd_sc_hd__a31o_2 _15599_ (.A1(\decode.regfile.registers_11[7] ),
    .A2(_11070_),
    .A3(_11470_),
    .B1(_11278_),
    .X(_11589_));
 sky130_fd_sc_hd__a21o_2 _15600_ (.A1(_11588_),
    .A2(_11315_),
    .B1(_11589_),
    .X(_11590_));
 sky130_fd_sc_hd__a2111o_2 _15601_ (.A1(_11046_),
    .A2(\decode.regfile.registers_12[7] ),
    .B1(_10649_),
    .C1(_11052_),
    .D1(_10632_),
    .X(_11591_));
 sky130_fd_sc_hd__a32o_2 _15602_ (.A1(\decode.regfile.registers_13[7] ),
    .A2(_10639_),
    .A3(_11187_),
    .B1(_11590_),
    .B2(_11591_),
    .X(_11592_));
 sky130_fd_sc_hd__o31a_2 _15603_ (.A1(_10651_),
    .A2(_10625_),
    .A3(_11054_),
    .B1(_11592_),
    .X(_11593_));
 sky130_fd_sc_hd__o221a_2 _15604_ (.A1(\decode.regfile.registers_16[7] ),
    .A2(_11359_),
    .B1(_11574_),
    .B2(_11593_),
    .C1(_11127_),
    .X(_11594_));
 sky130_fd_sc_hd__a21oi_2 _15605_ (.A1(\decode.regfile.registers_17[7] ),
    .A2(_11357_),
    .B1(_11594_),
    .Y(_11595_));
 sky130_fd_sc_hd__a21oi_2 _15606_ (.A1(\decode.regfile.registers_18[7] ),
    .A2(_11269_),
    .B1(_11271_),
    .Y(_11596_));
 sky130_fd_sc_hd__o21ai_2 _15607_ (.A1(_11269_),
    .A2(_11595_),
    .B1(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__o211a_2 _15608_ (.A1(\decode.regfile.registers_19[7] ),
    .A2(_11406_),
    .B1(_11325_),
    .C1(_11597_),
    .X(_11598_));
 sky130_fd_sc_hd__a211o_2 _15609_ (.A1(\decode.regfile.registers_20[7] ),
    .A2(_11103_),
    .B1(_11222_),
    .C1(_11598_),
    .X(_11599_));
 sky130_fd_sc_hd__o311a_2 _15610_ (.A1(\decode.regfile.registers_21[7] ),
    .A2(_11267_),
    .A3(_11099_),
    .B1(_11228_),
    .C1(_11599_),
    .X(_11600_));
 sky130_fd_sc_hd__o22a_2 _15611_ (.A1(\decode.regfile.registers_23[7] ),
    .A2(_11087_),
    .B1(_11573_),
    .B2(_11600_),
    .X(_11601_));
 sky130_fd_sc_hd__a31o_2 _15612_ (.A1(_10992_),
    .A2(_11066_),
    .A3(_11261_),
    .B1(_11601_),
    .X(_11602_));
 sky130_fd_sc_hd__o22a_2 _15613_ (.A1(\decode.regfile.registers_25[7] ),
    .A2(_11333_),
    .B1(_11336_),
    .B2(\decode.regfile.registers_24[7] ),
    .X(_11603_));
 sky130_fd_sc_hd__o2111a_2 _15614_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[7] ),
    .B1(_11349_),
    .C1(_10980_),
    .D1(_11564_),
    .X(_11604_));
 sky130_fd_sc_hd__a31o_2 _15615_ (.A1(_11236_),
    .A2(_11602_),
    .A3(_11603_),
    .B1(_11604_),
    .X(_11605_));
 sky130_fd_sc_hd__or3_2 _15616_ (.A(_11250_),
    .B(\decode.regfile.registers_27[7] ),
    .C(_11258_),
    .X(_11606_));
 sky130_fd_sc_hd__o2111a_2 _15617_ (.A1(_10960_),
    .A2(\decode.regfile.registers_28[7] ),
    .B1(_11067_),
    .C1(_11038_),
    .D1(_11440_),
    .X(_11607_));
 sky130_fd_sc_hd__a31o_2 _15618_ (.A1(_11403_),
    .A2(_11605_),
    .A3(_11606_),
    .B1(_11607_),
    .X(_11608_));
 sky130_fd_sc_hd__o221a_2 _15619_ (.A1(_11346_),
    .A2(_11253_),
    .B1(_11064_),
    .B2(\decode.regfile.registers_29[7] ),
    .C1(_11608_),
    .X(_11609_));
 sky130_fd_sc_hd__o221a_2 _15620_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[7] ),
    .B1(_11572_),
    .B2(_11609_),
    .C1(_11249_),
    .X(_00395_));
 sky130_fd_sc_hd__o2111a_2 _15621_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[8] ),
    .B1(_11039_),
    .C1(_11032_),
    .D1(_11033_),
    .X(_11610_));
 sky130_fd_sc_hd__o2111a_2 _15622_ (.A1(_10959_),
    .A2(\decode.regfile.registers_26[8] ),
    .B1(_11447_),
    .C1(_11348_),
    .D1(_10993_),
    .X(_11611_));
 sky130_fd_sc_hd__o2111a_2 _15623_ (.A1(_10957_),
    .A2(\decode.regfile.registers_22[8] ),
    .B1(_11450_),
    .C1(_10978_),
    .D1(_10990_),
    .X(_11612_));
 sky130_fd_sc_hd__o21ai_2 _15624_ (.A1(\decode.regfile.registers_17[8] ),
    .A2(_11128_),
    .B1(_11106_),
    .Y(_11613_));
 sky130_fd_sc_hd__buf_1 _15625_ (.A(_11292_),
    .X(_11614_));
 sky130_fd_sc_hd__o2bb2ai_2 _15626_ (.A1_N(\decode.regfile.registers_0[8] ),
    .A2_N(_11154_),
    .B1(_11503_),
    .B2(_11148_),
    .Y(_11615_));
 sky130_fd_sc_hd__and4_2 _15627_ (.A(\decode.regfile.registers_1[8] ),
    .B(_11117_),
    .C(_11057_),
    .D(_11109_),
    .X(_11616_));
 sky130_fd_sc_hd__o22ai_2 _15628_ (.A1(\decode.regfile.registers_2[8] ),
    .A2(_11369_),
    .B1(_11615_),
    .B2(_11616_),
    .Y(_11617_));
 sky130_fd_sc_hd__o2bb2a_2 _15629_ (.A1_N(\decode.regfile.registers_3[8] ),
    .A2_N(_11614_),
    .B1(_11367_),
    .B2(_10636_),
    .X(_11618_));
 sky130_fd_sc_hd__o21ai_2 _15630_ (.A1(_11614_),
    .A2(_11617_),
    .B1(_11618_),
    .Y(_11619_));
 sky130_fd_sc_hd__a2111o_2 _15631_ (.A1(_11313_),
    .A2(\decode.regfile.registers_4[8] ),
    .B1(_11191_),
    .C1(_10630_),
    .D1(_11462_),
    .X(_11620_));
 sky130_fd_sc_hd__a32o_2 _15632_ (.A1(\decode.regfile.registers_5[8] ),
    .A2(_10637_),
    .A3(_11139_),
    .B1(_11619_),
    .B2(_11620_),
    .X(_11621_));
 sky130_fd_sc_hd__a32o_2 _15633_ (.A1(\decode.regfile.registers_7[8] ),
    .A2(_11092_),
    .A3(_11167_),
    .B1(_11170_),
    .B2(\decode.regfile.registers_6[8] ),
    .X(_11622_));
 sky130_fd_sc_hd__a211o_2 _15634_ (.A1(_11136_),
    .A2(_11621_),
    .B1(_11622_),
    .C1(_11166_),
    .X(_11623_));
 sky130_fd_sc_hd__a21o_2 _15635_ (.A1(\decode.regfile.registers_8[8] ),
    .A2(_11045_),
    .B1(_11175_),
    .X(_11624_));
 sky130_fd_sc_hd__a221o_2 _15636_ (.A1(\decode.regfile.registers_9[8] ),
    .A2(_11547_),
    .B1(_11623_),
    .B2(_11624_),
    .C1(_11184_),
    .X(_11625_));
 sky130_fd_sc_hd__o211a_2 _15637_ (.A1(_11382_),
    .A2(\decode.regfile.registers_10[8] ),
    .B1(_11364_),
    .C1(_11625_),
    .X(_11626_));
 sky130_fd_sc_hd__a311o_2 _15638_ (.A1(\decode.regfile.registers_11[8] ),
    .A2(_11072_),
    .A3(_11205_),
    .B1(_11407_),
    .C1(_11626_),
    .X(_11627_));
 sky130_fd_sc_hd__a2111o_2 _15639_ (.A1(_11048_),
    .A2(\decode.regfile.registers_12[8] ),
    .B1(_10651_),
    .C1(_11054_),
    .D1(_10633_),
    .X(_11628_));
 sky130_fd_sc_hd__a32o_2 _15640_ (.A1(\decode.regfile.registers_13[8] ),
    .A2(_11225_),
    .A3(_11187_),
    .B1(_11627_),
    .B2(_11628_),
    .X(_11629_));
 sky130_fd_sc_hd__and3_2 _15641_ (.A(\decode.regfile.registers_15[8] ),
    .B(_11037_),
    .C(_11205_),
    .X(_11630_));
 sky130_fd_sc_hd__a221o_2 _15642_ (.A1(\decode.regfile.registers_14[8] ),
    .A2(_11208_),
    .B1(_11629_),
    .B2(_11199_),
    .C1(_11630_),
    .X(_11631_));
 sky130_fd_sc_hd__a32o_2 _15643_ (.A1(_11094_),
    .A2(_11114_),
    .A3(_11119_),
    .B1(_11203_),
    .B2(\decode.regfile.registers_16[8] ),
    .X(_11632_));
 sky130_fd_sc_hd__a21oi_2 _15644_ (.A1(_11124_),
    .A2(_11631_),
    .B1(_11632_),
    .Y(_11633_));
 sky130_fd_sc_hd__a21oi_2 _15645_ (.A1(\decode.regfile.registers_18[8] ),
    .A2(_11455_),
    .B1(_11456_),
    .Y(_11634_));
 sky130_fd_sc_hd__o21ai_2 _15646_ (.A1(_11613_),
    .A2(_11633_),
    .B1(_11634_),
    .Y(_11635_));
 sky130_fd_sc_hd__o41a_2 _15647_ (.A1(\decode.regfile.registers_19[8] ),
    .A2(_11049_),
    .A3(_11215_),
    .A4(_11217_),
    .B1(_11219_),
    .X(_11636_));
 sky130_fd_sc_hd__a221o_2 _15648_ (.A1(\decode.regfile.registers_20[8] ),
    .A2(_11103_),
    .B1(_11635_),
    .B2(_11636_),
    .C1(_11222_),
    .X(_11637_));
 sky130_fd_sc_hd__o311a_2 _15649_ (.A1(\decode.regfile.registers_21[8] ),
    .A2(_11061_),
    .A3(_11100_),
    .B1(_11229_),
    .C1(_11637_),
    .X(_11638_));
 sky130_fd_sc_hd__o22a_2 _15650_ (.A1(\decode.regfile.registers_23[8] ),
    .A2(_11088_),
    .B1(_11612_),
    .B2(_11638_),
    .X(_11639_));
 sky130_fd_sc_hd__o22a_2 _15651_ (.A1(\decode.regfile.registers_25[8] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[8] ),
    .X(_11640_));
 sky130_fd_sc_hd__o211a_2 _15652_ (.A1(_11075_),
    .A2(_11639_),
    .B1(_11640_),
    .C1(_11236_),
    .X(_11641_));
 sky130_fd_sc_hd__o32a_2 _15653_ (.A1(_11251_),
    .A2(_11259_),
    .A3(\decode.regfile.registers_27[8] ),
    .B1(_11611_),
    .B2(_11641_),
    .X(_11642_));
 sky130_fd_sc_hd__o22a_2 _15654_ (.A1(_11396_),
    .A2(\decode.regfile.registers_28[8] ),
    .B1(\decode.regfile.registers_29[8] ),
    .B2(_11255_),
    .X(_11643_));
 sky130_fd_sc_hd__o211a_2 _15655_ (.A1(_11445_),
    .A2(_11642_),
    .B1(_11643_),
    .C1(_11246_),
    .X(_11644_));
 sky130_fd_sc_hd__o221a_2 _15656_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[8] ),
    .B1(_11610_),
    .B2(_11644_),
    .C1(_11249_),
    .X(_00396_));
 sky130_fd_sc_hd__o2111a_2 _15657_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[9] ),
    .B1(_11039_),
    .C1(_11032_),
    .D1(_11033_),
    .X(_11645_));
 sky130_fd_sc_hd__buf_1 _15658_ (.A(_10961_),
    .X(_11646_));
 sky130_fd_sc_hd__or2_2 _15659_ (.A(_11493_),
    .B(\decode.regfile.registers_24[9] ),
    .X(_11647_));
 sky130_fd_sc_hd__or4_2 _15660_ (.A(_11059_),
    .B(_10976_),
    .C(_11048_),
    .D(_11085_),
    .X(_11648_));
 sky130_fd_sc_hd__a32o_2 _15661_ (.A1(_11094_),
    .A2(_11119_),
    .A3(_11093_),
    .B1(_11101_),
    .B2(\decode.regfile.registers_20[9] ),
    .X(_11649_));
 sky130_fd_sc_hd__a221o_2 _15662_ (.A1(\decode.regfile.registers_11[9] ),
    .A2(_11180_),
    .B1(_11509_),
    .B2(\decode.regfile.registers_10[9] ),
    .C1(_11186_),
    .X(_11650_));
 sky130_fd_sc_hd__a221o_2 _15663_ (.A1(\decode.regfile.registers_7[9] ),
    .A2(_11465_),
    .B1(_11466_),
    .B2(\decode.regfile.registers_6[9] ),
    .C1(_11281_),
    .X(_11651_));
 sky130_fd_sc_hd__or3b_2 _15664_ (.A(_10647_),
    .B(_11097_),
    .C_N(\decode.regfile.registers_5[9] ),
    .X(_11652_));
 sky130_fd_sc_hd__mux2_2 _15665_ (.A0(\decode.regfile.registers_1[9] ),
    .A1(\decode.regfile.registers_0[9] ),
    .S(_11300_),
    .X(_11653_));
 sky130_fd_sc_hd__o32a_2 _15666_ (.A1(_10659_),
    .A2(_10654_),
    .A3(_11150_),
    .B1(\decode.regfile.registers_2[9] ),
    .B2(_11296_),
    .X(_11654_));
 sky130_fd_sc_hd__o21ai_2 _15667_ (.A1(_11156_),
    .A2(_11653_),
    .B1(_11654_),
    .Y(_11655_));
 sky130_fd_sc_hd__or4b_2 _15668_ (.A(_10659_),
    .B(_10654_),
    .C(_11150_),
    .D_N(\decode.regfile.registers_3[9] ),
    .X(_11656_));
 sky130_fd_sc_hd__nand2_2 _15669_ (.A(_11313_),
    .B(\decode.regfile.registers_4[9] ),
    .Y(_11657_));
 sky130_fd_sc_hd__a32o_2 _15670_ (.A1(_11375_),
    .A2(_11655_),
    .A3(_11656_),
    .B1(_11657_),
    .B2(_11138_),
    .X(_11658_));
 sky130_fd_sc_hd__o2bb2a_2 _15671_ (.A1_N(_11652_),
    .A2_N(_11658_),
    .B1(_11318_),
    .B2(_11084_),
    .X(_11659_));
 sky130_fd_sc_hd__o221a_2 _15672_ (.A1(\decode.regfile.registers_8[9] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(\decode.regfile.registers_9[9] ),
    .C1(_11131_),
    .X(_11660_));
 sky130_fd_sc_hd__o21a_2 _15673_ (.A1(_11651_),
    .A2(_11659_),
    .B1(_11660_),
    .X(_11661_));
 sky130_fd_sc_hd__or2_2 _15674_ (.A(_11650_),
    .B(_11661_),
    .X(_11662_));
 sky130_fd_sc_hd__o22a_2 _15675_ (.A1(_11194_),
    .A2(\decode.regfile.registers_12[9] ),
    .B1(\decode.regfile.registers_13[9] ),
    .B2(_11196_),
    .X(_11663_));
 sky130_fd_sc_hd__a221o_2 _15676_ (.A1(\decode.regfile.registers_14[9] ),
    .A2(_11207_),
    .B1(_11273_),
    .B2(\decode.regfile.registers_15[9] ),
    .C1(_11201_),
    .X(_11664_));
 sky130_fd_sc_hd__a31o_2 _15677_ (.A1(_11198_),
    .A2(_11662_),
    .A3(_11663_),
    .B1(_11664_),
    .X(_11665_));
 sky130_fd_sc_hd__o211a_2 _15678_ (.A1(_11123_),
    .A2(\decode.regfile.registers_16[9] ),
    .B1(_11126_),
    .C1(_11665_),
    .X(_11666_));
 sky130_fd_sc_hd__a41o_2 _15679_ (.A1(\decode.regfile.registers_17[9] ),
    .A2(_10652_),
    .A3(_11112_),
    .A4(_11118_),
    .B1(_11666_),
    .X(_11667_));
 sky130_fd_sc_hd__o2111a_2 _15680_ (.A1(\decode.regfile.registers_18[9] ),
    .A2(_10642_),
    .B1(_11112_),
    .C1(_10652_),
    .D1(_10633_),
    .X(_11668_));
 sky130_fd_sc_hd__a21o_2 _15681_ (.A1(_11106_),
    .A2(_11667_),
    .B1(_11668_),
    .X(_11669_));
 sky130_fd_sc_hd__o211a_2 _15682_ (.A1(\decode.regfile.registers_19[9] ),
    .A2(_11354_),
    .B1(_11218_),
    .C1(_11669_),
    .X(_11670_));
 sky130_fd_sc_hd__o221a_2 _15683_ (.A1(\decode.regfile.registers_21[9] ),
    .A2(_11648_),
    .B1(_11649_),
    .B2(_11670_),
    .C1(_11227_),
    .X(_11671_));
 sky130_fd_sc_hd__a211o_2 _15684_ (.A1(\decode.regfile.registers_22[9] ),
    .A2(_11096_),
    .B1(_11232_),
    .C1(_11671_),
    .X(_11672_));
 sky130_fd_sc_hd__o221a_2 _15685_ (.A1(\decode.regfile.registers_23[9] ),
    .A2(_11262_),
    .B1(_11089_),
    .B2(_11493_),
    .C1(_11672_),
    .X(_11673_));
 sky130_fd_sc_hd__a41o_2 _15686_ (.A1(_11079_),
    .A2(_11244_),
    .A3(_11261_),
    .A4(_11647_),
    .B1(_11673_),
    .X(_11674_));
 sky130_fd_sc_hd__or3_2 _15687_ (.A(_11050_),
    .B(\decode.regfile.registers_25[9] ),
    .C(_11090_),
    .X(_11675_));
 sky130_fd_sc_hd__buf_1 _15688_ (.A(_11080_),
    .X(_11676_));
 sky130_fd_sc_hd__o2111a_2 _15689_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[9] ),
    .B1(_11676_),
    .C1(_10980_),
    .D1(_11564_),
    .X(_11677_));
 sky130_fd_sc_hd__a31o_2 _15690_ (.A1(_11236_),
    .A2(_11674_),
    .A3(_11675_),
    .B1(_11677_),
    .X(_11678_));
 sky130_fd_sc_hd__buf_1 _15691_ (.A(_11050_),
    .X(_11679_));
 sky130_fd_sc_hd__or3_2 _15692_ (.A(_11679_),
    .B(\decode.regfile.registers_27[9] ),
    .C(_11258_),
    .X(_11680_));
 sky130_fd_sc_hd__buf_1 _15693_ (.A(_11037_),
    .X(_11681_));
 sky130_fd_sc_hd__o2111a_2 _15694_ (.A1(_10960_),
    .A2(\decode.regfile.registers_28[9] ),
    .B1(_11067_),
    .C1(_11681_),
    .D1(_11440_),
    .X(_11682_));
 sky130_fd_sc_hd__a31o_2 _15695_ (.A1(_11403_),
    .A2(_11678_),
    .A3(_11680_),
    .B1(_11682_),
    .X(_11683_));
 sky130_fd_sc_hd__o221a_2 _15696_ (.A1(_11646_),
    .A2(_11253_),
    .B1(_11064_),
    .B2(\decode.regfile.registers_29[9] ),
    .C1(_11683_),
    .X(_11684_));
 sky130_fd_sc_hd__o221a_2 _15697_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[9] ),
    .B1(_11645_),
    .B2(_11684_),
    .C1(_11249_),
    .X(_00397_));
 sky130_fd_sc_hd__o2111a_2 _15698_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[10] ),
    .B1(_11039_),
    .C1(_11032_),
    .D1(_11033_),
    .X(_11685_));
 sky130_fd_sc_hd__o2111a_2 _15699_ (.A1(_11446_),
    .A2(\decode.regfile.registers_26[10] ),
    .B1(_11447_),
    .C1(_10981_),
    .D1(_11448_),
    .X(_11686_));
 sky130_fd_sc_hd__or2_2 _15700_ (.A(_11435_),
    .B(\decode.regfile.registers_24[10] ),
    .X(_11687_));
 sky130_fd_sc_hd__o2111a_2 _15701_ (.A1(\decode.regfile.registers_18[10] ),
    .A2(_10955_),
    .B1(_11114_),
    .C1(_11094_),
    .D1(_10977_),
    .X(_11688_));
 sky130_fd_sc_hd__or3_2 _15702_ (.A(_11191_),
    .B(_10630_),
    .C(_11051_),
    .X(_11689_));
 sky130_fd_sc_hd__buf_1 _15703_ (.A(_11689_),
    .X(_11690_));
 sky130_fd_sc_hd__a31o_2 _15704_ (.A1(\decode.regfile.registers_11[10] ),
    .A2(_11071_),
    .A3(_11204_),
    .B1(_11407_),
    .X(_11691_));
 sky130_fd_sc_hd__and2_2 _15705_ (.A(_11046_),
    .B(\decode.regfile.registers_10[10] ),
    .X(_11692_));
 sky130_fd_sc_hd__a21oi_2 _15706_ (.A1(\decode.regfile.registers_8[10] ),
    .A2(_11046_),
    .B1(_11175_),
    .Y(_11693_));
 sky130_fd_sc_hd__a31o_2 _15707_ (.A1(\decode.regfile.registers_3[10] ),
    .A2(_11110_),
    .A3(_11141_),
    .B1(_11146_),
    .X(_11694_));
 sky130_fd_sc_hd__and4_2 _15708_ (.A(\decode.regfile.registers_1[10] ),
    .B(_11117_),
    .C(_11057_),
    .D(_11157_),
    .X(_11695_));
 sky130_fd_sc_hd__a2bb2o_2 _15709_ (.A1_N(_11129_),
    .A2_N(_11298_),
    .B1(_11300_),
    .B2(\decode.regfile.registers_0[10] ),
    .X(_11696_));
 sky130_fd_sc_hd__o221a_2 _15710_ (.A1(\decode.regfile.registers_2[10] ),
    .A2(_11369_),
    .B1(_11695_),
    .B2(_11696_),
    .C1(_11152_),
    .X(_11697_));
 sky130_fd_sc_hd__o32a_2 _15711_ (.A1(\decode.regfile.registers_4[10] ),
    .A2(_11192_),
    .A3(_11410_),
    .B1(_11694_),
    .B2(_11697_),
    .X(_11698_));
 sky130_fd_sc_hd__mux2_2 _15712_ (.A0(_11698_),
    .A1(\decode.regfile.registers_5[10] ),
    .S(_11291_),
    .X(_11699_));
 sky130_fd_sc_hd__a221o_2 _15713_ (.A1(\decode.regfile.registers_7[10] ),
    .A2(_11378_),
    .B1(_11170_),
    .B2(\decode.regfile.registers_6[10] ),
    .C1(_11166_),
    .X(_11700_));
 sky130_fd_sc_hd__a21oi_2 _15714_ (.A1(_11136_),
    .A2(_11699_),
    .B1(_11700_),
    .Y(_11701_));
 sky130_fd_sc_hd__o2bb2a_2 _15715_ (.A1_N(\decode.regfile.registers_9[10] ),
    .A2_N(_11547_),
    .B1(_10638_),
    .B2(_11132_),
    .X(_11702_));
 sky130_fd_sc_hd__o21ai_2 _15716_ (.A1(_11693_),
    .A2(_11701_),
    .B1(_11702_),
    .Y(_11703_));
 sky130_fd_sc_hd__o21a_2 _15717_ (.A1(_11132_),
    .A2(_11692_),
    .B1(_11703_),
    .X(_11704_));
 sky130_fd_sc_hd__o32a_2 _15718_ (.A1(\decode.regfile.registers_12[10] ),
    .A2(_10640_),
    .A3(_11690_),
    .B1(_11691_),
    .B2(_11704_),
    .X(_11705_));
 sky130_fd_sc_hd__mux2_2 _15719_ (.A0(_11705_),
    .A1(\decode.regfile.registers_13[10] ),
    .S(_11276_),
    .X(_11706_));
 sky130_fd_sc_hd__a32o_2 _15720_ (.A1(\decode.regfile.registers_15[10] ),
    .A2(_11037_),
    .A3(_11205_),
    .B1(_11208_),
    .B2(\decode.regfile.registers_14[10] ),
    .X(_11707_));
 sky130_fd_sc_hd__a21oi_2 _15721_ (.A1(_11199_),
    .A2(_11706_),
    .B1(_11707_),
    .Y(_11708_));
 sky130_fd_sc_hd__a21oi_2 _15722_ (.A1(\decode.regfile.registers_16[10] ),
    .A2(_11203_),
    .B1(_11357_),
    .Y(_11709_));
 sky130_fd_sc_hd__o21ai_2 _15723_ (.A1(_11203_),
    .A2(_11708_),
    .B1(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__o221a_2 _15724_ (.A1(_11059_),
    .A2(_11149_),
    .B1(_11128_),
    .B2(\decode.regfile.registers_17[10] ),
    .C1(_11710_),
    .X(_11711_));
 sky130_fd_sc_hd__o221a_2 _15725_ (.A1(\decode.regfile.registers_19[10] ),
    .A2(_11453_),
    .B1(_11688_),
    .B2(_11711_),
    .C1(_11454_),
    .X(_11712_));
 sky130_fd_sc_hd__a211o_2 _15726_ (.A1(\decode.regfile.registers_20[10] ),
    .A2(_11452_),
    .B1(_11223_),
    .C1(_11712_),
    .X(_11713_));
 sky130_fd_sc_hd__o32a_2 _15727_ (.A1(_10956_),
    .A2(_11217_),
    .A3(_11085_),
    .B1(\decode.regfile.registers_21[10] ),
    .B2(_11648_),
    .X(_11714_));
 sky130_fd_sc_hd__a221o_2 _15728_ (.A1(\decode.regfile.registers_22[10] ),
    .A2(_11096_),
    .B1(_11713_),
    .B2(_11714_),
    .C1(_11232_),
    .X(_11715_));
 sky130_fd_sc_hd__o22a_2 _15729_ (.A1(_11435_),
    .A2(_11089_),
    .B1(\decode.regfile.registers_23[10] ),
    .B2(_11087_),
    .X(_11716_));
 sky130_fd_sc_hd__a22o_2 _15730_ (.A1(_11074_),
    .A2(_11687_),
    .B1(_11715_),
    .B2(_11716_),
    .X(_11717_));
 sky130_fd_sc_hd__o311a_2 _15731_ (.A1(_11250_),
    .A2(\decode.regfile.registers_25[10] ),
    .A3(_11090_),
    .B1(_11486_),
    .C1(_11717_),
    .X(_11718_));
 sky130_fd_sc_hd__o32a_2 _15732_ (.A1(_11251_),
    .A2(_11259_),
    .A3(\decode.regfile.registers_27[10] ),
    .B1(_11686_),
    .B2(_11718_),
    .X(_11719_));
 sky130_fd_sc_hd__o221a_2 _15733_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[10] ),
    .B1(\decode.regfile.registers_29[10] ),
    .B2(_11255_),
    .C1(_11246_),
    .X(_11720_));
 sky130_fd_sc_hd__o21a_2 _15734_ (.A1(_11445_),
    .A2(_11719_),
    .B1(_11720_),
    .X(_11721_));
 sky130_fd_sc_hd__o221a_2 _15735_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[10] ),
    .B1(_11685_),
    .B2(_11721_),
    .C1(_11249_),
    .X(_00398_));
 sky130_fd_sc_hd__buf_1 _15736_ (.A(_11038_),
    .X(_11722_));
 sky130_fd_sc_hd__buf_1 _15737_ (.A(_10981_),
    .X(_11723_));
 sky130_fd_sc_hd__buf_1 _15738_ (.A(_10994_),
    .X(_11724_));
 sky130_fd_sc_hd__o2111a_2 _15739_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[11] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_11725_));
 sky130_fd_sc_hd__a21o_2 _15740_ (.A1(\decode.regfile.registers_19[11] ),
    .A2(_11271_),
    .B1(_11101_),
    .X(_11726_));
 sky130_fd_sc_hd__a221o_2 _15741_ (.A1(\decode.regfile.registers_14[11] ),
    .A2(_11360_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[11] ),
    .C1(_11202_),
    .X(_11727_));
 sky130_fd_sc_hd__a31o_2 _15742_ (.A1(\decode.regfile.registers_11[11] ),
    .A2(_11071_),
    .A3(_11470_),
    .B1(_11278_),
    .X(_11728_));
 sky130_fd_sc_hd__a2bb2o_2 _15743_ (.A1_N(\decode.regfile.registers_2[11] ),
    .A2_N(_11296_),
    .B1(_11141_),
    .B2(_11109_),
    .X(_11729_));
 sky130_fd_sc_hd__and4_2 _15744_ (.A(\decode.regfile.registers_1[11] ),
    .B(_11117_),
    .C(_11057_),
    .D(_11109_),
    .X(_11730_));
 sky130_fd_sc_hd__a211oi_2 _15745_ (.A1(_11154_),
    .A2(\decode.regfile.registers_0[11] ),
    .B1(_11156_),
    .C1(_11730_),
    .Y(_11731_));
 sky130_fd_sc_hd__o2bb2a_2 _15746_ (.A1_N(\decode.regfile.registers_3[11] ),
    .A2_N(_11614_),
    .B1(_11367_),
    .B2(_11178_),
    .X(_11732_));
 sky130_fd_sc_hd__o21ai_2 _15747_ (.A1(_11729_),
    .A2(_11731_),
    .B1(_11732_),
    .Y(_11733_));
 sky130_fd_sc_hd__a2111o_2 _15748_ (.A1(_11043_),
    .A2(\decode.regfile.registers_4[11] ),
    .B1(_11503_),
    .C1(_10629_),
    .D1(_11083_),
    .X(_11734_));
 sky130_fd_sc_hd__a22oi_2 _15749_ (.A1(\decode.regfile.registers_5[11] ),
    .A2(_11291_),
    .B1(_11733_),
    .B2(_11734_),
    .Y(_11735_));
 sky130_fd_sc_hd__a221oi_2 _15750_ (.A1(\decode.regfile.registers_7[11] ),
    .A2(_11465_),
    .B1(_11466_),
    .B2(\decode.regfile.registers_6[11] ),
    .C1(_11166_),
    .Y(_11736_));
 sky130_fd_sc_hd__o21ai_2 _15751_ (.A1(_11289_),
    .A2(_11735_),
    .B1(_11736_),
    .Y(_11737_));
 sky130_fd_sc_hd__a21o_2 _15752_ (.A1(\decode.regfile.registers_8[11] ),
    .A2(_11044_),
    .B1(_11174_),
    .X(_11738_));
 sky130_fd_sc_hd__a221o_2 _15753_ (.A1(\decode.regfile.registers_9[11] ),
    .A2(_11547_),
    .B1(_11737_),
    .B2(_11738_),
    .C1(_11509_),
    .X(_11739_));
 sky130_fd_sc_hd__o211a_2 _15754_ (.A1(_11382_),
    .A2(\decode.regfile.registers_10[11] ),
    .B1(_11315_),
    .C1(_11739_),
    .X(_11740_));
 sky130_fd_sc_hd__a2111o_2 _15755_ (.A1(_11046_),
    .A2(\decode.regfile.registers_12[11] ),
    .B1(_10649_),
    .C1(_11052_),
    .D1(_10631_),
    .X(_11741_));
 sky130_fd_sc_hd__o21a_2 _15756_ (.A1(_11728_),
    .A2(_11740_),
    .B1(_11741_),
    .X(_11742_));
 sky130_fd_sc_hd__and3_2 _15757_ (.A(\decode.regfile.registers_13[11] ),
    .B(_10639_),
    .C(_11187_),
    .X(_11743_));
 sky130_fd_sc_hd__o32a_2 _15758_ (.A1(_10650_),
    .A2(_10625_),
    .A3(_11053_),
    .B1(_11742_),
    .B2(_11743_),
    .X(_11744_));
 sky130_fd_sc_hd__o221a_2 _15759_ (.A1(\decode.regfile.registers_16[11] ),
    .A2(_11359_),
    .B1(_11727_),
    .B2(_11744_),
    .C1(_11127_),
    .X(_11745_));
 sky130_fd_sc_hd__a211o_2 _15760_ (.A1(\decode.regfile.registers_17[11] ),
    .A2(_11357_),
    .B1(_11745_),
    .C1(_11268_),
    .X(_11746_));
 sky130_fd_sc_hd__o311a_2 _15761_ (.A1(\decode.regfile.registers_18[11] ),
    .A2(_11059_),
    .A3(_11149_),
    .B1(_11406_),
    .C1(_11746_),
    .X(_11747_));
 sky130_fd_sc_hd__o221a_2 _15762_ (.A1(\decode.regfile.registers_20[11] ),
    .A2(_11219_),
    .B1(_11726_),
    .B2(_11747_),
    .C1(_11648_),
    .X(_11748_));
 sky130_fd_sc_hd__a211o_2 _15763_ (.A1(\decode.regfile.registers_21[11] ),
    .A2(_11222_),
    .B1(_11096_),
    .C1(_11748_),
    .X(_11749_));
 sky130_fd_sc_hd__o211a_2 _15764_ (.A1(\decode.regfile.registers_22[11] ),
    .A2(_11228_),
    .B1(_11262_),
    .C1(_11749_),
    .X(_11750_));
 sky130_fd_sc_hd__a211o_2 _15765_ (.A1(\decode.regfile.registers_23[11] ),
    .A2(_11232_),
    .B1(_11074_),
    .C1(_11750_),
    .X(_11751_));
 sky130_fd_sc_hd__o22a_2 _15766_ (.A1(\decode.regfile.registers_25[11] ),
    .A2(_11333_),
    .B1(_11336_),
    .B2(\decode.regfile.registers_24[11] ),
    .X(_11752_));
 sky130_fd_sc_hd__o2111a_2 _15767_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[11] ),
    .B1(_11676_),
    .C1(_10980_),
    .D1(_11564_),
    .X(_11753_));
 sky130_fd_sc_hd__a31o_2 _15768_ (.A1(_11260_),
    .A2(_11751_),
    .A3(_11752_),
    .B1(_11753_),
    .X(_11754_));
 sky130_fd_sc_hd__or3_2 _15769_ (.A(_11679_),
    .B(\decode.regfile.registers_27[11] ),
    .C(_11258_),
    .X(_11755_));
 sky130_fd_sc_hd__buf_1 _15770_ (.A(_10959_),
    .X(_11756_));
 sky130_fd_sc_hd__o2111a_2 _15771_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[11] ),
    .B1(_11067_),
    .C1(_11681_),
    .D1(_11440_),
    .X(_11757_));
 sky130_fd_sc_hd__a31o_2 _15772_ (.A1(_11403_),
    .A2(_11754_),
    .A3(_11755_),
    .B1(_11757_),
    .X(_11758_));
 sky130_fd_sc_hd__o221a_2 _15773_ (.A1(_11646_),
    .A2(_11253_),
    .B1(_11064_),
    .B2(\decode.regfile.registers_29[11] ),
    .C1(_11758_),
    .X(_11759_));
 sky130_fd_sc_hd__buf_1 _15774_ (.A(_11248_),
    .X(_11760_));
 sky130_fd_sc_hd__o221a_2 _15775_ (.A1(_11344_),
    .A2(\decode.regfile.registers_31[11] ),
    .B1(_11725_),
    .B2(_11759_),
    .C1(_11760_),
    .X(_00399_));
 sky130_fd_sc_hd__buf_1 _15776_ (.A(_11243_),
    .X(_11761_));
 sky130_fd_sc_hd__o2111a_2 _15777_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[12] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_11762_));
 sky130_fd_sc_hd__o2111a_2 _15778_ (.A1(_11446_),
    .A2(\decode.regfile.registers_26[12] ),
    .B1(_11447_),
    .C1(_11348_),
    .D1(_10993_),
    .X(_11763_));
 sky130_fd_sc_hd__o2111a_2 _15779_ (.A1(_11435_),
    .A2(\decode.regfile.registers_22[12] ),
    .B1(_11450_),
    .C1(_10979_),
    .D1(_10991_),
    .X(_11764_));
 sky130_fd_sc_hd__nor2_2 _15780_ (.A(\decode.regfile.registers_10[12] ),
    .B(_11382_),
    .Y(_11765_));
 sky130_fd_sc_hd__o2bb2ai_2 _15781_ (.A1_N(\decode.regfile.registers_0[12] ),
    .A2_N(_11154_),
    .B1(_11190_),
    .B2(_11298_),
    .Y(_11766_));
 sky130_fd_sc_hd__a21o_2 _15782_ (.A1(\decode.regfile.registers_1[12] ),
    .A2(_11539_),
    .B1(_11766_),
    .X(_11767_));
 sky130_fd_sc_hd__o311a_2 _15783_ (.A1(\decode.regfile.registers_2[12] ),
    .A2(_10647_),
    .A3(_11149_),
    .B1(_11152_),
    .C1(_11767_),
    .X(_11768_));
 sky130_fd_sc_hd__a311o_2 _15784_ (.A1(\decode.regfile.registers_3[12] ),
    .A2(_11111_),
    .A3(_11167_),
    .B1(_11146_),
    .C1(_11768_),
    .X(_11769_));
 sky130_fd_sc_hd__a2111o_2 _15785_ (.A1(_11044_),
    .A2(\decode.regfile.registers_4[12] ),
    .B1(_10648_),
    .C1(_10631_),
    .D1(_11084_),
    .X(_11770_));
 sky130_fd_sc_hd__a22oi_2 _15786_ (.A1(\decode.regfile.registers_5[12] ),
    .A2(_11291_),
    .B1(_11769_),
    .B2(_11770_),
    .Y(_11771_));
 sky130_fd_sc_hd__a221oi_2 _15787_ (.A1(\decode.regfile.registers_7[12] ),
    .A2(_11378_),
    .B1(_11170_),
    .B2(\decode.regfile.registers_6[12] ),
    .C1(_11166_),
    .Y(_11772_));
 sky130_fd_sc_hd__o21ai_2 _15788_ (.A1(_11289_),
    .A2(_11771_),
    .B1(_11772_),
    .Y(_11773_));
 sky130_fd_sc_hd__a21o_2 _15789_ (.A1(\decode.regfile.registers_8[12] ),
    .A2(_11046_),
    .B1(_11175_),
    .X(_11774_));
 sky130_fd_sc_hd__a221oi_2 _15790_ (.A1(\decode.regfile.registers_9[12] ),
    .A2(_11547_),
    .B1(_11773_),
    .B2(_11774_),
    .C1(_11184_),
    .Y(_11775_));
 sky130_fd_sc_hd__a41o_2 _15791_ (.A1(_11058_),
    .A2(_10632_),
    .A3(_10640_),
    .A4(_11071_),
    .B1(_11775_),
    .X(_11776_));
 sky130_fd_sc_hd__o2bb2a_2 _15792_ (.A1_N(\decode.regfile.registers_11[12] ),
    .A2_N(_11181_),
    .B1(_11690_),
    .B2(_10640_),
    .X(_11777_));
 sky130_fd_sc_hd__o21ai_2 _15793_ (.A1(_11765_),
    .A2(_11776_),
    .B1(_11777_),
    .Y(_11778_));
 sky130_fd_sc_hd__a2111o_2 _15794_ (.A1(_11047_),
    .A2(\decode.regfile.registers_12[12] ),
    .B1(_10651_),
    .C1(_11053_),
    .D1(_10633_),
    .X(_11779_));
 sky130_fd_sc_hd__a32o_2 _15795_ (.A1(\decode.regfile.registers_13[12] ),
    .A2(_10642_),
    .A3(_11187_),
    .B1(_11778_),
    .B2(_11779_),
    .X(_11780_));
 sky130_fd_sc_hd__a32o_2 _15796_ (.A1(\decode.regfile.registers_15[12] ),
    .A2(_11037_),
    .A3(_11205_),
    .B1(_11208_),
    .B2(\decode.regfile.registers_14[12] ),
    .X(_11781_));
 sky130_fd_sc_hd__a21oi_2 _15797_ (.A1(_11199_),
    .A2(_11780_),
    .B1(_11781_),
    .Y(_11782_));
 sky130_fd_sc_hd__a21oi_2 _15798_ (.A1(\decode.regfile.registers_16[12] ),
    .A2(_11203_),
    .B1(_11357_),
    .Y(_11783_));
 sky130_fd_sc_hd__o21ai_2 _15799_ (.A1(_11203_),
    .A2(_11782_),
    .B1(_11783_),
    .Y(_11784_));
 sky130_fd_sc_hd__o32a_2 _15800_ (.A1(_11225_),
    .A2(_11125_),
    .A3(_11216_),
    .B1(\decode.regfile.registers_17[12] ),
    .B2(_11128_),
    .X(_11785_));
 sky130_fd_sc_hd__a221o_2 _15801_ (.A1(\decode.regfile.registers_18[12] ),
    .A2(_11455_),
    .B1(_11784_),
    .B2(_11785_),
    .C1(_11456_),
    .X(_11786_));
 sky130_fd_sc_hd__o211a_2 _15802_ (.A1(\decode.regfile.registers_19[12] ),
    .A2(_11453_),
    .B1(_11454_),
    .C1(_11786_),
    .X(_11787_));
 sky130_fd_sc_hd__a211o_2 _15803_ (.A1(\decode.regfile.registers_20[12] ),
    .A2(_11452_),
    .B1(_11223_),
    .C1(_11787_),
    .X(_11788_));
 sky130_fd_sc_hd__o311a_2 _15804_ (.A1(\decode.regfile.registers_21[12] ),
    .A2(_11062_),
    .A3(_11100_),
    .B1(_11229_),
    .C1(_11788_),
    .X(_11789_));
 sky130_fd_sc_hd__o22a_2 _15805_ (.A1(\decode.regfile.registers_23[12] ),
    .A2(_11088_),
    .B1(_11764_),
    .B2(_11789_),
    .X(_11790_));
 sky130_fd_sc_hd__o22a_2 _15806_ (.A1(\decode.regfile.registers_25[12] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[12] ),
    .X(_11791_));
 sky130_fd_sc_hd__o211a_2 _15807_ (.A1(_11075_),
    .A2(_11790_),
    .B1(_11791_),
    .C1(_11486_),
    .X(_11792_));
 sky130_fd_sc_hd__o32a_2 _15808_ (.A1(_11251_),
    .A2(_11259_),
    .A3(\decode.regfile.registers_27[12] ),
    .B1(_11763_),
    .B2(_11792_),
    .X(_11793_));
 sky130_fd_sc_hd__o221a_2 _15809_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[12] ),
    .B1(\decode.regfile.registers_29[12] ),
    .B2(_11255_),
    .C1(_11246_),
    .X(_11794_));
 sky130_fd_sc_hd__o21a_2 _15810_ (.A1(_11445_),
    .A2(_11793_),
    .B1(_11794_),
    .X(_11795_));
 sky130_fd_sc_hd__o221a_2 _15811_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[12] ),
    .B1(_11762_),
    .B2(_11795_),
    .C1(_11760_),
    .X(_00400_));
 sky130_fd_sc_hd__o2111a_2 _15812_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[13] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_11796_));
 sky130_fd_sc_hd__o2111a_2 _15813_ (.A1(_11263_),
    .A2(\decode.regfile.registers_22[13] ),
    .B1(_11404_),
    .C1(_10978_),
    .D1(_11265_),
    .X(_11797_));
 sky130_fd_sc_hd__o2111a_2 _15814_ (.A1(\decode.regfile.registers_18[13] ),
    .A2(_11225_),
    .B1(_11113_),
    .C1(_10988_),
    .D1(_10976_),
    .X(_11798_));
 sky130_fd_sc_hd__a221o_2 _15815_ (.A1(\decode.regfile.registers_14[13] ),
    .A2(_11207_),
    .B1(_11273_),
    .B2(\decode.regfile.registers_15[13] ),
    .C1(_11361_),
    .X(_11799_));
 sky130_fd_sc_hd__o2bb2a_2 _15816_ (.A1_N(_11069_),
    .A2_N(_11167_),
    .B1(\decode.regfile.registers_10[13] ),
    .B2(_11381_),
    .X(_11800_));
 sky130_fd_sc_hd__a221o_2 _15817_ (.A1(\decode.regfile.registers_7[13] ),
    .A2(_11308_),
    .B1(_11169_),
    .B2(\decode.regfile.registers_6[13] ),
    .C1(_11165_),
    .X(_11801_));
 sky130_fd_sc_hd__and3_2 _15818_ (.A(\decode.regfile.registers_5[13] ),
    .B(_11178_),
    .C(_11138_),
    .X(_11802_));
 sky130_fd_sc_hd__a31o_2 _15819_ (.A1(\decode.regfile.registers_3[13] ),
    .A2(_11157_),
    .A3(_11140_),
    .B1(_11145_),
    .X(_11803_));
 sky130_fd_sc_hd__nand4_2 _15820_ (.A(\decode.regfile.registers_1[13] ),
    .B(_11115_),
    .C(_11056_),
    .D(_11108_),
    .Y(_11804_));
 sky130_fd_sc_hd__nand2_2 _15821_ (.A(_11153_),
    .B(\decode.regfile.registers_0[13] ),
    .Y(_11805_));
 sky130_fd_sc_hd__o211ai_2 _15822_ (.A1(_10645_),
    .A2(_11147_),
    .B1(_11804_),
    .C1(_11805_),
    .Y(_11806_));
 sky130_fd_sc_hd__o211a_2 _15823_ (.A1(\decode.regfile.registers_2[13] ),
    .A2(_11295_),
    .B1(_11151_),
    .C1(_11806_),
    .X(_11807_));
 sky130_fd_sc_hd__a2111o_2 _15824_ (.A1(_11042_),
    .A2(\decode.regfile.registers_4[13] ),
    .B1(_11129_),
    .C1(_10628_),
    .D1(_11082_),
    .X(_11808_));
 sky130_fd_sc_hd__o21a_2 _15825_ (.A1(_11803_),
    .A2(_11807_),
    .B1(_11808_),
    .X(_11809_));
 sky130_fd_sc_hd__o32a_2 _15826_ (.A1(_10647_),
    .A2(_10624_),
    .A3(_11462_),
    .B1(_11802_),
    .B2(_11809_),
    .X(_11810_));
 sky130_fd_sc_hd__o22ai_2 _15827_ (.A1(\decode.regfile.registers_8[13] ),
    .A2(_11284_),
    .B1(_11801_),
    .B2(_11810_),
    .Y(_11811_));
 sky130_fd_sc_hd__o2bb2a_2 _15828_ (.A1_N(\decode.regfile.registers_9[13] ),
    .A2_N(_11547_),
    .B1(_11192_),
    .B2(_11131_),
    .X(_11812_));
 sky130_fd_sc_hd__o21ai_2 _15829_ (.A1(_11547_),
    .A2(_11811_),
    .B1(_11812_),
    .Y(_11813_));
 sky130_fd_sc_hd__a32o_2 _15830_ (.A1(\decode.regfile.registers_11[13] ),
    .A2(_11070_),
    .A3(_11470_),
    .B1(_11800_),
    .B2(_11813_),
    .X(_11814_));
 sky130_fd_sc_hd__o22a_2 _15831_ (.A1(\decode.regfile.registers_12[13] ),
    .A2(_11689_),
    .B1(_11278_),
    .B2(_11814_),
    .X(_11815_));
 sky130_fd_sc_hd__o32a_2 _15832_ (.A1(\decode.regfile.registers_13[13] ),
    .A2(_11046_),
    .A3(_11689_),
    .B1(_11318_),
    .B2(_11052_),
    .X(_11816_));
 sky130_fd_sc_hd__o21a_2 _15833_ (.A1(_11276_),
    .A2(_11815_),
    .B1(_11816_),
    .X(_11817_));
 sky130_fd_sc_hd__o22a_2 _15834_ (.A1(\decode.regfile.registers_16[13] ),
    .A2(_11123_),
    .B1(_11799_),
    .B2(_11817_),
    .X(_11818_));
 sky130_fd_sc_hd__mux2_2 _15835_ (.A0(_11818_),
    .A1(\decode.regfile.registers_17[13] ),
    .S(_11356_),
    .X(_11819_));
 sky130_fd_sc_hd__o31a_2 _15836_ (.A1(_11225_),
    .A2(_11125_),
    .A3(_11216_),
    .B1(_11819_),
    .X(_11820_));
 sky130_fd_sc_hd__o221a_2 _15837_ (.A1(\decode.regfile.registers_19[13] ),
    .A2(_11406_),
    .B1(_11798_),
    .B2(_11820_),
    .C1(_11219_),
    .X(_11821_));
 sky130_fd_sc_hd__a211o_2 _15838_ (.A1(\decode.regfile.registers_20[13] ),
    .A2(_11103_),
    .B1(_11327_),
    .C1(_11821_),
    .X(_11822_));
 sky130_fd_sc_hd__o311a_2 _15839_ (.A1(\decode.regfile.registers_21[13] ),
    .A2(_11267_),
    .A3(_11099_),
    .B1(_11228_),
    .C1(_11822_),
    .X(_11823_));
 sky130_fd_sc_hd__o22a_2 _15840_ (.A1(\decode.regfile.registers_23[13] ),
    .A2(_11087_),
    .B1(_11797_),
    .B2(_11823_),
    .X(_11824_));
 sky130_fd_sc_hd__a31o_2 _15841_ (.A1(_10992_),
    .A2(_11066_),
    .A3(_11261_),
    .B1(_11824_),
    .X(_11825_));
 sky130_fd_sc_hd__o22a_2 _15842_ (.A1(\decode.regfile.registers_25[13] ),
    .A2(_11333_),
    .B1(_11336_),
    .B2(\decode.regfile.registers_24[13] ),
    .X(_11826_));
 sky130_fd_sc_hd__o2111a_2 _15843_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[13] ),
    .B1(_11676_),
    .C1(_11338_),
    .D1(_11564_),
    .X(_11827_));
 sky130_fd_sc_hd__a31o_2 _15844_ (.A1(_11260_),
    .A2(_11825_),
    .A3(_11826_),
    .B1(_11827_),
    .X(_11828_));
 sky130_fd_sc_hd__or3_2 _15845_ (.A(_11679_),
    .B(\decode.regfile.registers_27[13] ),
    .C(_11258_),
    .X(_11829_));
 sky130_fd_sc_hd__o2111a_2 _15846_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[13] ),
    .B1(_11067_),
    .C1(_11681_),
    .D1(_11440_),
    .X(_11830_));
 sky130_fd_sc_hd__a31o_2 _15847_ (.A1(_11403_),
    .A2(_11828_),
    .A3(_11829_),
    .B1(_11830_),
    .X(_11831_));
 sky130_fd_sc_hd__o221a_2 _15848_ (.A1(_11646_),
    .A2(_11253_),
    .B1(_11064_),
    .B2(\decode.regfile.registers_29[13] ),
    .C1(_11831_),
    .X(_11832_));
 sky130_fd_sc_hd__o221a_2 _15849_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[13] ),
    .B1(_11796_),
    .B2(_11832_),
    .C1(_11760_),
    .X(_00401_));
 sky130_fd_sc_hd__o2111a_2 _15850_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[14] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_11833_));
 sky130_fd_sc_hd__buf_1 _15851_ (.A(_11252_),
    .X(_11834_));
 sky130_fd_sc_hd__or2_2 _15852_ (.A(_11493_),
    .B(\decode.regfile.registers_24[14] ),
    .X(_11835_));
 sky130_fd_sc_hd__o2111a_2 _15853_ (.A1(_10956_),
    .A2(\decode.regfile.registers_22[14] ),
    .B1(_11093_),
    .C1(_11264_),
    .D1(_11265_),
    .X(_11836_));
 sky130_fd_sc_hd__o2111a_2 _15854_ (.A1(\decode.regfile.registers_18[14] ),
    .A2(_11225_),
    .B1(_11113_),
    .C1(_10988_),
    .D1(_10976_),
    .X(_11837_));
 sky130_fd_sc_hd__a221o_2 _15855_ (.A1(\decode.regfile.registers_14[14] ),
    .A2(_11207_),
    .B1(_11273_),
    .B2(\decode.regfile.registers_15[14] ),
    .C1(_11201_),
    .X(_11838_));
 sky130_fd_sc_hd__a31o_2 _15856_ (.A1(\decode.regfile.registers_11[14] ),
    .A2(_11070_),
    .A3(_11470_),
    .B1(_11278_),
    .X(_11839_));
 sky130_fd_sc_hd__a31o_2 _15857_ (.A1(\decode.regfile.registers_9[14] ),
    .A2(_11280_),
    .A3(_11134_),
    .B1(_11183_),
    .X(_11840_));
 sky130_fd_sc_hd__and3_2 _15858_ (.A(\decode.regfile.registers_5[14] ),
    .B(_10636_),
    .C(_11138_),
    .X(_11841_));
 sky130_fd_sc_hd__inv_2 _15859_ (.A(\decode.regfile.registers_0[14] ),
    .Y(_11842_));
 sky130_fd_sc_hd__nand2_2 _15860_ (.A(\decode.regfile.registers_1[14] ),
    .B(_11539_),
    .Y(_11843_));
 sky130_fd_sc_hd__o211ai_2 _15861_ (.A1(_11842_),
    .A2(_11539_),
    .B1(_11843_),
    .C1(_11296_),
    .Y(_11844_));
 sky130_fd_sc_hd__o211ai_2 _15862_ (.A1(\decode.regfile.registers_2[14] ),
    .A2(_11369_),
    .B1(_11152_),
    .C1(_11844_),
    .Y(_11845_));
 sky130_fd_sc_hd__o2bb2a_2 _15863_ (.A1_N(\decode.regfile.registers_3[14] ),
    .A2_N(_11614_),
    .B1(_11367_),
    .B2(_11178_),
    .X(_11846_));
 sky130_fd_sc_hd__a2111o_2 _15864_ (.A1(_11042_),
    .A2(\decode.regfile.registers_4[14] ),
    .B1(_10646_),
    .C1(_10628_),
    .D1(_11082_),
    .X(_11847_));
 sky130_fd_sc_hd__a21boi_2 _15865_ (.A1(_11845_),
    .A2(_11846_),
    .B1_N(_11847_),
    .Y(_11848_));
 sky130_fd_sc_hd__o21ai_2 _15866_ (.A1(_11841_),
    .A2(_11848_),
    .B1(_11136_),
    .Y(_11849_));
 sky130_fd_sc_hd__a221oi_2 _15867_ (.A1(\decode.regfile.registers_7[14] ),
    .A2(_11465_),
    .B1(_11169_),
    .B2(\decode.regfile.registers_6[14] ),
    .C1(_11165_),
    .Y(_11850_));
 sky130_fd_sc_hd__nand2_2 _15868_ (.A(_11849_),
    .B(_11850_),
    .Y(_11851_));
 sky130_fd_sc_hd__o211a_2 _15869_ (.A1(\decode.regfile.registers_8[14] ),
    .A2(_11175_),
    .B1(_11365_),
    .C1(_11851_),
    .X(_11852_));
 sky130_fd_sc_hd__o2bb2a_2 _15870_ (.A1_N(_11070_),
    .A2_N(_11167_),
    .B1(\decode.regfile.registers_10[14] ),
    .B2(_11381_),
    .X(_11853_));
 sky130_fd_sc_hd__o21a_2 _15871_ (.A1(_11840_),
    .A2(_11852_),
    .B1(_11853_),
    .X(_11854_));
 sky130_fd_sc_hd__o22ai_2 _15872_ (.A1(\decode.regfile.registers_12[14] ),
    .A2(_11194_),
    .B1(_11839_),
    .B2(_11854_),
    .Y(_11855_));
 sky130_fd_sc_hd__o21ai_2 _15873_ (.A1(\decode.regfile.registers_13[14] ),
    .A2(_11196_),
    .B1(_11198_),
    .Y(_11856_));
 sky130_fd_sc_hd__a21oi_2 _15874_ (.A1(_11196_),
    .A2(_11855_),
    .B1(_11856_),
    .Y(_11857_));
 sky130_fd_sc_hd__o22a_2 _15875_ (.A1(\decode.regfile.registers_16[14] ),
    .A2(_11123_),
    .B1(_11838_),
    .B2(_11857_),
    .X(_11858_));
 sky130_fd_sc_hd__mux2_2 _15876_ (.A0(_11858_),
    .A1(\decode.regfile.registers_17[14] ),
    .S(_11356_),
    .X(_11859_));
 sky130_fd_sc_hd__o31a_2 _15877_ (.A1(_11225_),
    .A2(_11125_),
    .A3(_11104_),
    .B1(_11859_),
    .X(_11860_));
 sky130_fd_sc_hd__o221a_2 _15878_ (.A1(\decode.regfile.registers_19[14] ),
    .A2(_11354_),
    .B1(_11837_),
    .B2(_11860_),
    .C1(_11325_),
    .X(_11861_));
 sky130_fd_sc_hd__a211o_2 _15879_ (.A1(\decode.regfile.registers_20[14] ),
    .A2(_11102_),
    .B1(_11327_),
    .C1(_11861_),
    .X(_11862_));
 sky130_fd_sc_hd__o311a_2 _15880_ (.A1(\decode.regfile.registers_21[14] ),
    .A2(_11060_),
    .A3(_11098_),
    .B1(_11227_),
    .C1(_11862_),
    .X(_11863_));
 sky130_fd_sc_hd__o221a_2 _15881_ (.A1(\decode.regfile.registers_23[14] ),
    .A2(_11262_),
    .B1(_11836_),
    .B2(_11863_),
    .C1(_11335_),
    .X(_11864_));
 sky130_fd_sc_hd__a41o_2 _15882_ (.A1(_11079_),
    .A2(_11244_),
    .A3(_11261_),
    .A4(_11835_),
    .B1(_11864_),
    .X(_11865_));
 sky130_fd_sc_hd__or3_2 _15883_ (.A(_11050_),
    .B(\decode.regfile.registers_25[14] ),
    .C(_11090_),
    .X(_11866_));
 sky130_fd_sc_hd__o2111a_2 _15884_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[14] ),
    .B1(_11676_),
    .C1(_11338_),
    .D1(_11564_),
    .X(_11867_));
 sky130_fd_sc_hd__a31o_2 _15885_ (.A1(_11260_),
    .A2(_11865_),
    .A3(_11866_),
    .B1(_11867_),
    .X(_11868_));
 sky130_fd_sc_hd__buf_1 _15886_ (.A(_11257_),
    .X(_11869_));
 sky130_fd_sc_hd__or3_2 _15887_ (.A(_11679_),
    .B(\decode.regfile.registers_27[14] ),
    .C(_11869_),
    .X(_11870_));
 sky130_fd_sc_hd__buf_1 _15888_ (.A(_11066_),
    .X(_11871_));
 sky130_fd_sc_hd__o2111a_2 _15889_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[14] ),
    .B1(_11871_),
    .C1(_11681_),
    .D1(_11440_),
    .X(_11872_));
 sky130_fd_sc_hd__a31o_2 _15890_ (.A1(_11403_),
    .A2(_11868_),
    .A3(_11870_),
    .B1(_11872_),
    .X(_11873_));
 sky130_fd_sc_hd__o221a_2 _15891_ (.A1(_11646_),
    .A2(_11834_),
    .B1(_11064_),
    .B2(\decode.regfile.registers_29[14] ),
    .C1(_11873_),
    .X(_11874_));
 sky130_fd_sc_hd__o221a_2 _15892_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[14] ),
    .B1(_11833_),
    .B2(_11874_),
    .C1(_11760_),
    .X(_00402_));
 sky130_fd_sc_hd__o2111a_2 _15893_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[15] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_11875_));
 sky130_fd_sc_hd__o2111a_2 _15894_ (.A1(_11446_),
    .A2(\decode.regfile.registers_26[15] ),
    .B1(_11447_),
    .C1(_11348_),
    .D1(_10993_),
    .X(_11876_));
 sky130_fd_sc_hd__o2111a_2 _15895_ (.A1(_11435_),
    .A2(\decode.regfile.registers_22[15] ),
    .B1(_11450_),
    .C1(_10979_),
    .D1(_10991_),
    .X(_11877_));
 sky130_fd_sc_hd__a221o_2 _15896_ (.A1(\decode.regfile.registers_14[15] ),
    .A2(_11208_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[15] ),
    .C1(_11202_),
    .X(_11878_));
 sky130_fd_sc_hd__nand2_2 _15897_ (.A(\decode.regfile.registers_13[15] ),
    .B(_11276_),
    .Y(_11879_));
 sky130_fd_sc_hd__or3b_2 _15898_ (.A(_11191_),
    .B(_11097_),
    .C_N(\decode.regfile.registers_5[15] ),
    .X(_11880_));
 sky130_fd_sc_hd__a31o_2 _15899_ (.A1(\decode.regfile.registers_3[15] ),
    .A2(_11110_),
    .A3(_11141_),
    .B1(_11146_),
    .X(_11881_));
 sky130_fd_sc_hd__o2bb2ai_2 _15900_ (.A1_N(\decode.regfile.registers_0[15] ),
    .A2_N(_11300_),
    .B1(_11129_),
    .B2(_11298_),
    .Y(_11882_));
 sky130_fd_sc_hd__a21o_2 _15901_ (.A1(\decode.regfile.registers_1[15] ),
    .A2(_11539_),
    .B1(_11882_),
    .X(_11883_));
 sky130_fd_sc_hd__o311a_2 _15902_ (.A1(\decode.regfile.registers_2[15] ),
    .A2(_11503_),
    .A3(_11148_),
    .B1(_11152_),
    .C1(_11883_),
    .X(_11884_));
 sky130_fd_sc_hd__a2111o_2 _15903_ (.A1(_11043_),
    .A2(\decode.regfile.registers_4[15] ),
    .B1(_11503_),
    .C1(_10629_),
    .D1(_11462_),
    .X(_11885_));
 sky130_fd_sc_hd__o21ai_2 _15904_ (.A1(_11881_),
    .A2(_11884_),
    .B1(_11885_),
    .Y(_11886_));
 sky130_fd_sc_hd__nand2_2 _15905_ (.A(_11880_),
    .B(_11886_),
    .Y(_11887_));
 sky130_fd_sc_hd__a221o_2 _15906_ (.A1(\decode.regfile.registers_7[15] ),
    .A2(_11465_),
    .B1(_11466_),
    .B2(\decode.regfile.registers_6[15] ),
    .C1(_11165_),
    .X(_11888_));
 sky130_fd_sc_hd__a21o_2 _15907_ (.A1(_11136_),
    .A2(_11887_),
    .B1(_11888_),
    .X(_11889_));
 sky130_fd_sc_hd__a21o_2 _15908_ (.A1(\decode.regfile.registers_8[15] ),
    .A2(_11045_),
    .B1(_11175_),
    .X(_11890_));
 sky130_fd_sc_hd__a31o_2 _15909_ (.A1(\decode.regfile.registers_9[15] ),
    .A2(_11280_),
    .A3(_11281_),
    .B1(_11183_),
    .X(_11891_));
 sky130_fd_sc_hd__a21o_2 _15910_ (.A1(_11889_),
    .A2(_11890_),
    .B1(_11891_),
    .X(_11892_));
 sky130_fd_sc_hd__o2bb2a_2 _15911_ (.A1_N(_11070_),
    .A2_N(_11470_),
    .B1(\decode.regfile.registers_10[15] ),
    .B2(_11381_),
    .X(_11893_));
 sky130_fd_sc_hd__a221o_2 _15912_ (.A1(\decode.regfile.registers_11[15] ),
    .A2(_11181_),
    .B1(_11892_),
    .B2(_11893_),
    .C1(_11407_),
    .X(_11894_));
 sky130_fd_sc_hd__o211ai_2 _15913_ (.A1(_11194_),
    .A2(\decode.regfile.registers_12[15] ),
    .B1(_11196_),
    .C1(_11894_),
    .Y(_11895_));
 sky130_fd_sc_hd__o2bb2a_2 _15914_ (.A1_N(_11879_),
    .A2_N(_11895_),
    .B1(_11054_),
    .B2(_11318_),
    .X(_11896_));
 sky130_fd_sc_hd__o22a_2 _15915_ (.A1(\decode.regfile.registers_16[15] ),
    .A2(_11124_),
    .B1(_11878_),
    .B2(_11896_),
    .X(_11897_));
 sky130_fd_sc_hd__a31o_2 _15916_ (.A1(_11094_),
    .A2(_11113_),
    .A3(_11119_),
    .B1(_11897_),
    .X(_11898_));
 sky130_fd_sc_hd__o32a_2 _15917_ (.A1(_11225_),
    .A2(_11125_),
    .A3(_11216_),
    .B1(\decode.regfile.registers_17[15] ),
    .B2(_11128_),
    .X(_11899_));
 sky130_fd_sc_hd__a221o_2 _15918_ (.A1(\decode.regfile.registers_18[15] ),
    .A2(_11455_),
    .B1(_11898_),
    .B2(_11899_),
    .C1(_11456_),
    .X(_11900_));
 sky130_fd_sc_hd__o211a_2 _15919_ (.A1(\decode.regfile.registers_19[15] ),
    .A2(_11453_),
    .B1(_11454_),
    .C1(_11900_),
    .X(_11901_));
 sky130_fd_sc_hd__a211o_2 _15920_ (.A1(\decode.regfile.registers_20[15] ),
    .A2(_11452_),
    .B1(_11223_),
    .C1(_11901_),
    .X(_11902_));
 sky130_fd_sc_hd__o311a_2 _15921_ (.A1(\decode.regfile.registers_21[15] ),
    .A2(_11062_),
    .A3(_11100_),
    .B1(_11229_),
    .C1(_11902_),
    .X(_11903_));
 sky130_fd_sc_hd__o22a_2 _15922_ (.A1(\decode.regfile.registers_23[15] ),
    .A2(_11088_),
    .B1(_11877_),
    .B2(_11903_),
    .X(_11904_));
 sky130_fd_sc_hd__o22a_2 _15923_ (.A1(\decode.regfile.registers_25[15] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[15] ),
    .X(_11905_));
 sky130_fd_sc_hd__o211a_2 _15924_ (.A1(_11075_),
    .A2(_11904_),
    .B1(_11905_),
    .C1(_11486_),
    .X(_11906_));
 sky130_fd_sc_hd__o32a_2 _15925_ (.A1(_11251_),
    .A2(_11259_),
    .A3(\decode.regfile.registers_27[15] ),
    .B1(_11876_),
    .B2(_11906_),
    .X(_11907_));
 sky130_fd_sc_hd__o221a_2 _15926_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[15] ),
    .B1(\decode.regfile.registers_29[15] ),
    .B2(_11255_),
    .C1(_11246_),
    .X(_11908_));
 sky130_fd_sc_hd__o21a_2 _15927_ (.A1(_11445_),
    .A2(_11907_),
    .B1(_11908_),
    .X(_11909_));
 sky130_fd_sc_hd__o221a_2 _15928_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[15] ),
    .B1(_11875_),
    .B2(_11909_),
    .C1(_11760_),
    .X(_00403_));
 sky130_fd_sc_hd__o2111a_2 _15929_ (.A1(_11571_),
    .A2(\decode.regfile.registers_30[16] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_11910_));
 sky130_fd_sc_hd__o2111a_2 _15930_ (.A1(_10959_),
    .A2(\decode.regfile.registers_26[16] ),
    .B1(_11447_),
    .C1(_11348_),
    .D1(_10993_),
    .X(_11911_));
 sky130_fd_sc_hd__o2111a_2 _15931_ (.A1(_10957_),
    .A2(\decode.regfile.registers_22[16] ),
    .B1(_11450_),
    .C1(_10978_),
    .D1(_10990_),
    .X(_11912_));
 sky130_fd_sc_hd__a31o_2 _15932_ (.A1(\decode.regfile.registers_15[16] ),
    .A2(_11036_),
    .A3(_11204_),
    .B1(_11361_),
    .X(_11913_));
 sky130_fd_sc_hd__or4b_2 _15933_ (.A(_10660_),
    .B(_10655_),
    .C(_11297_),
    .D_N(\decode.regfile.registers_3[16] ),
    .X(_11914_));
 sky130_fd_sc_hd__and4_2 _15934_ (.A(\decode.regfile.registers_1[16] ),
    .B(_11116_),
    .C(_11137_),
    .D(_11157_),
    .X(_11915_));
 sky130_fd_sc_hd__a211o_2 _15935_ (.A1(_11154_),
    .A2(\decode.regfile.registers_0[16] ),
    .B1(_11156_),
    .C1(_11915_),
    .X(_11916_));
 sky130_fd_sc_hd__o221ai_2 _15936_ (.A1(\decode.regfile.registers_2[16] ),
    .A2(_11369_),
    .B1(_11297_),
    .B2(_11121_),
    .C1(_11916_),
    .Y(_11917_));
 sky130_fd_sc_hd__o211ai_2 _15937_ (.A1(_11410_),
    .A2(_11192_),
    .B1(_11914_),
    .C1(_11917_),
    .Y(_11918_));
 sky130_fd_sc_hd__a2111o_2 _15938_ (.A1(_11313_),
    .A2(\decode.regfile.registers_4[16] ),
    .B1(_10647_),
    .C1(_10630_),
    .D1(_11462_),
    .X(_11919_));
 sky130_fd_sc_hd__a22oi_2 _15939_ (.A1(\decode.regfile.registers_5[16] ),
    .A2(_11291_),
    .B1(_11918_),
    .B2(_11919_),
    .Y(_11920_));
 sky130_fd_sc_hd__a221oi_2 _15940_ (.A1(\decode.regfile.registers_7[16] ),
    .A2(_11465_),
    .B1(_11466_),
    .B2(\decode.regfile.registers_6[16] ),
    .C1(_11281_),
    .Y(_11921_));
 sky130_fd_sc_hd__o21ai_2 _15941_ (.A1(_11289_),
    .A2(_11920_),
    .B1(_11921_),
    .Y(_11922_));
 sky130_fd_sc_hd__o221a_2 _15942_ (.A1(\decode.regfile.registers_8[16] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(\decode.regfile.registers_9[16] ),
    .C1(_11131_),
    .X(_11923_));
 sky130_fd_sc_hd__a221o_2 _15943_ (.A1(\decode.regfile.registers_11[16] ),
    .A2(_11180_),
    .B1(_11183_),
    .B2(\decode.regfile.registers_10[16] ),
    .C1(_11278_),
    .X(_11924_));
 sky130_fd_sc_hd__a21o_2 _15944_ (.A1(_11922_),
    .A2(_11923_),
    .B1(_11924_),
    .X(_11925_));
 sky130_fd_sc_hd__a2111o_2 _15945_ (.A1(_11045_),
    .A2(\decode.regfile.registers_12[16] ),
    .B1(_10649_),
    .C1(_11051_),
    .D1(_10631_),
    .X(_11926_));
 sky130_fd_sc_hd__a32o_2 _15946_ (.A1(\decode.regfile.registers_13[16] ),
    .A2(_10639_),
    .A3(_11186_),
    .B1(_11925_),
    .B2(_11926_),
    .X(_11927_));
 sky130_fd_sc_hd__a22o_2 _15947_ (.A1(\decode.regfile.registers_14[16] ),
    .A2(_11360_),
    .B1(_11927_),
    .B2(_11198_),
    .X(_11928_));
 sky130_fd_sc_hd__o22a_2 _15948_ (.A1(_11123_),
    .A2(\decode.regfile.registers_16[16] ),
    .B1(_11913_),
    .B2(_11928_),
    .X(_11929_));
 sky130_fd_sc_hd__a31o_2 _15949_ (.A1(_10652_),
    .A2(_11112_),
    .A3(_11118_),
    .B1(_11929_),
    .X(_11930_));
 sky130_fd_sc_hd__o221a_2 _15950_ (.A1(_11059_),
    .A2(_11149_),
    .B1(_11128_),
    .B2(\decode.regfile.registers_17[16] ),
    .C1(_11930_),
    .X(_11931_));
 sky130_fd_sc_hd__a211o_2 _15951_ (.A1(\decode.regfile.registers_18[16] ),
    .A2(_11455_),
    .B1(_11456_),
    .C1(_11931_),
    .X(_11932_));
 sky130_fd_sc_hd__o211a_2 _15952_ (.A1(\decode.regfile.registers_19[16] ),
    .A2(_11453_),
    .B1(_11219_),
    .C1(_11932_),
    .X(_11933_));
 sky130_fd_sc_hd__a211o_2 _15953_ (.A1(\decode.regfile.registers_20[16] ),
    .A2(_11452_),
    .B1(_11222_),
    .C1(_11933_),
    .X(_11934_));
 sky130_fd_sc_hd__o311a_2 _15954_ (.A1(\decode.regfile.registers_21[16] ),
    .A2(_11061_),
    .A3(_11100_),
    .B1(_11229_),
    .C1(_11934_),
    .X(_11935_));
 sky130_fd_sc_hd__o22a_2 _15955_ (.A1(\decode.regfile.registers_23[16] ),
    .A2(_11088_),
    .B1(_11912_),
    .B2(_11935_),
    .X(_11936_));
 sky130_fd_sc_hd__o22a_2 _15956_ (.A1(\decode.regfile.registers_25[16] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[16] ),
    .X(_11937_));
 sky130_fd_sc_hd__o211a_2 _15957_ (.A1(_11075_),
    .A2(_11936_),
    .B1(_11937_),
    .C1(_11236_),
    .X(_11938_));
 sky130_fd_sc_hd__o32a_2 _15958_ (.A1(_11250_),
    .A2(_11259_),
    .A3(\decode.regfile.registers_27[16] ),
    .B1(_11911_),
    .B2(_11938_),
    .X(_11939_));
 sky130_fd_sc_hd__o22a_2 _15959_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[16] ),
    .B1(\decode.regfile.registers_29[16] ),
    .B2(_11255_),
    .X(_11940_));
 sky130_fd_sc_hd__o211a_2 _15960_ (.A1(_11445_),
    .A2(_11939_),
    .B1(_11940_),
    .C1(_11246_),
    .X(_11941_));
 sky130_fd_sc_hd__o221a_2 _15961_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[16] ),
    .B1(_11910_),
    .B2(_11941_),
    .C1(_11760_),
    .X(_00404_));
 sky130_fd_sc_hd__buf_1 _15962_ (.A(_10961_),
    .X(_11942_));
 sky130_fd_sc_hd__o2111a_2 _15963_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[17] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_11943_));
 sky130_fd_sc_hd__buf_1 _15964_ (.A(_11063_),
    .X(_11944_));
 sky130_fd_sc_hd__o2111a_2 _15965_ (.A1(_11435_),
    .A2(\decode.regfile.registers_24[17] ),
    .B1(_11244_),
    .C1(_11080_),
    .D1(_11079_),
    .X(_11945_));
 sky130_fd_sc_hd__o2111a_2 _15966_ (.A1(_11263_),
    .A2(\decode.regfile.registers_22[17] ),
    .B1(_11404_),
    .C1(_11264_),
    .D1(_11265_),
    .X(_11946_));
 sky130_fd_sc_hd__nand2_2 _15967_ (.A(\decode.regfile.registers_21[17] ),
    .B(_11222_),
    .Y(_11947_));
 sky130_fd_sc_hd__nor2_2 _15968_ (.A(\decode.regfile.registers_19[17] ),
    .B(_11406_),
    .Y(_11948_));
 sky130_fd_sc_hd__a31o_2 _15969_ (.A1(\decode.regfile.registers_9[17] ),
    .A2(_11280_),
    .A3(_11134_),
    .B1(_11183_),
    .X(_11949_));
 sky130_fd_sc_hd__a32o_2 _15970_ (.A1(\decode.regfile.registers_7[17] ),
    .A2(_11092_),
    .A3(_11142_),
    .B1(_11169_),
    .B2(\decode.regfile.registers_6[17] ),
    .X(_11950_));
 sky130_fd_sc_hd__and3_2 _15971_ (.A(\decode.regfile.registers_5[17] ),
    .B(_10636_),
    .C(_11138_),
    .X(_11951_));
 sky130_fd_sc_hd__and2_2 _15972_ (.A(_11042_),
    .B(\decode.regfile.registers_4[17] ),
    .X(_11952_));
 sky130_fd_sc_hd__a31o_2 _15973_ (.A1(\decode.regfile.registers_3[17] ),
    .A2(_11109_),
    .A3(_11140_),
    .B1(_11145_),
    .X(_11953_));
 sky130_fd_sc_hd__nand4_2 _15974_ (.A(\decode.regfile.registers_1[17] ),
    .B(_11116_),
    .C(_11056_),
    .D(_11108_),
    .Y(_11954_));
 sky130_fd_sc_hd__nand2_2 _15975_ (.A(_11153_),
    .B(\decode.regfile.registers_0[17] ),
    .Y(_11955_));
 sky130_fd_sc_hd__o211ai_2 _15976_ (.A1(_11129_),
    .A2(_11147_),
    .B1(_11954_),
    .C1(_11955_),
    .Y(_11956_));
 sky130_fd_sc_hd__o221a_2 _15977_ (.A1(\decode.regfile.registers_2[17] ),
    .A2(_11295_),
    .B1(_11150_),
    .B2(_11121_),
    .C1(_11956_),
    .X(_11957_));
 sky130_fd_sc_hd__o22a_2 _15978_ (.A1(_11367_),
    .A2(_11952_),
    .B1(_11953_),
    .B2(_11957_),
    .X(_11958_));
 sky130_fd_sc_hd__o21ai_2 _15979_ (.A1(_11951_),
    .A2(_11958_),
    .B1(_11135_),
    .Y(_11959_));
 sky130_fd_sc_hd__nand3b_2 _15980_ (.A_N(_11950_),
    .B(_11959_),
    .C(_11284_),
    .Y(_11960_));
 sky130_fd_sc_hd__o211a_2 _15981_ (.A1(\decode.regfile.registers_8[17] ),
    .A2(_11285_),
    .B1(_11287_),
    .C1(_11960_),
    .X(_11961_));
 sky130_fd_sc_hd__o32a_2 _15982_ (.A1(\decode.regfile.registers_10[17] ),
    .A2(_10638_),
    .A3(_11132_),
    .B1(_11949_),
    .B2(_11961_),
    .X(_11962_));
 sky130_fd_sc_hd__o32a_2 _15983_ (.A1(_10649_),
    .A2(_10631_),
    .A3(_11052_),
    .B1(\decode.regfile.registers_11[17] ),
    .B2(_11315_),
    .X(_11963_));
 sky130_fd_sc_hd__o21a_2 _15984_ (.A1(_11181_),
    .A2(_11962_),
    .B1(_11963_),
    .X(_11964_));
 sky130_fd_sc_hd__a221o_2 _15985_ (.A1(\decode.regfile.registers_13[17] ),
    .A2(_11276_),
    .B1(_11407_),
    .B2(\decode.regfile.registers_12[17] ),
    .C1(_11964_),
    .X(_11965_));
 sky130_fd_sc_hd__a221o_2 _15986_ (.A1(\decode.regfile.registers_14[17] ),
    .A2(_11360_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[17] ),
    .C1(_11202_),
    .X(_11966_));
 sky130_fd_sc_hd__a21o_2 _15987_ (.A1(_11199_),
    .A2(_11965_),
    .B1(_11966_),
    .X(_11967_));
 sky130_fd_sc_hd__o211a_2 _15988_ (.A1(_11124_),
    .A2(\decode.regfile.registers_16[17] ),
    .B1(_11127_),
    .C1(_11967_),
    .X(_11968_));
 sky130_fd_sc_hd__a41o_2 _15989_ (.A1(\decode.regfile.registers_17[17] ),
    .A2(_11094_),
    .A3(_11114_),
    .A4(_11119_),
    .B1(_11968_),
    .X(_11969_));
 sky130_fd_sc_hd__o2111a_2 _15990_ (.A1(\decode.regfile.registers_18[17] ),
    .A2(_10955_),
    .B1(_11114_),
    .C1(_11094_),
    .D1(_10976_),
    .X(_11970_));
 sky130_fd_sc_hd__a21oi_2 _15991_ (.A1(_11106_),
    .A2(_11969_),
    .B1(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__o21ai_2 _15992_ (.A1(_11948_),
    .A2(_11971_),
    .B1(_11454_),
    .Y(_11972_));
 sky130_fd_sc_hd__o221ai_2 _15993_ (.A1(_11060_),
    .A2(_11098_),
    .B1(_11454_),
    .B2(\decode.regfile.registers_20[17] ),
    .C1(_11972_),
    .Y(_11973_));
 sky130_fd_sc_hd__a21oi_2 _15994_ (.A1(_11947_),
    .A2(_11973_),
    .B1(_11096_),
    .Y(_11974_));
 sky130_fd_sc_hd__o221a_2 _15995_ (.A1(\decode.regfile.registers_23[17] ),
    .A2(_11262_),
    .B1(_11946_),
    .B2(_11974_),
    .C1(_11336_),
    .X(_11975_));
 sky130_fd_sc_hd__o32a_2 _15996_ (.A1(_11076_),
    .A2(_11090_),
    .A3(\decode.regfile.registers_25[17] ),
    .B1(_11945_),
    .B2(_11975_),
    .X(_11976_));
 sky130_fd_sc_hd__o2111a_2 _15997_ (.A1(_10959_),
    .A2(\decode.regfile.registers_26[17] ),
    .B1(_11349_),
    .C1(_10980_),
    .D1(_11347_),
    .X(_11977_));
 sky130_fd_sc_hd__a21o_2 _15998_ (.A1(_11976_),
    .A2(_11486_),
    .B1(_11977_),
    .X(_11978_));
 sky130_fd_sc_hd__or3_2 _15999_ (.A(_11679_),
    .B(\decode.regfile.registers_27[17] ),
    .C(_11869_),
    .X(_11979_));
 sky130_fd_sc_hd__o2111a_2 _16000_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[17] ),
    .B1(_11871_),
    .C1(_11681_),
    .D1(_11440_),
    .X(_11980_));
 sky130_fd_sc_hd__a31o_2 _16001_ (.A1(_11403_),
    .A2(_11978_),
    .A3(_11979_),
    .B1(_11980_),
    .X(_11981_));
 sky130_fd_sc_hd__o221a_2 _16002_ (.A1(_11646_),
    .A2(_11834_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[17] ),
    .C1(_11981_),
    .X(_11982_));
 sky130_fd_sc_hd__o221a_2 _16003_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[17] ),
    .B1(_11943_),
    .B2(_11982_),
    .C1(_11760_),
    .X(_00405_));
 sky130_fd_sc_hd__o2111a_2 _16004_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[18] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_11983_));
 sky130_fd_sc_hd__o2111a_2 _16005_ (.A1(_11446_),
    .A2(\decode.regfile.registers_26[18] ),
    .B1(_11447_),
    .C1(_11348_),
    .D1(_10993_),
    .X(_11984_));
 sky130_fd_sc_hd__o2111a_2 _16006_ (.A1(_11493_),
    .A2(\decode.regfile.registers_22[18] ),
    .B1(_11450_),
    .C1(_10979_),
    .D1(_10991_),
    .X(_11985_));
 sky130_fd_sc_hd__a221o_2 _16007_ (.A1(\decode.regfile.registers_14[18] ),
    .A2(_11207_),
    .B1(_11273_),
    .B2(\decode.regfile.registers_15[18] ),
    .C1(_11361_),
    .X(_11986_));
 sky130_fd_sc_hd__a221o_2 _16008_ (.A1(\decode.regfile.registers_11[18] ),
    .A2(_11180_),
    .B1(_11509_),
    .B2(\decode.regfile.registers_10[18] ),
    .C1(_11186_),
    .X(_11987_));
 sky130_fd_sc_hd__a221o_2 _16009_ (.A1(\decode.regfile.registers_7[18] ),
    .A2(_11465_),
    .B1(_11466_),
    .B2(\decode.regfile.registers_6[18] ),
    .C1(_11281_),
    .X(_11988_));
 sky130_fd_sc_hd__and3_2 _16010_ (.A(\decode.regfile.registers_5[18] ),
    .B(_11192_),
    .C(_11139_),
    .X(_11989_));
 sky130_fd_sc_hd__nand2_2 _16011_ (.A(_11371_),
    .B(\decode.regfile.registers_0[18] ),
    .Y(_11990_));
 sky130_fd_sc_hd__nand2_2 _16012_ (.A(\decode.regfile.registers_1[18] ),
    .B(_11539_),
    .Y(_11991_));
 sky130_fd_sc_hd__nor2_2 _16013_ (.A(\decode.regfile.registers_2[18] ),
    .B(_11295_),
    .Y(_11992_));
 sky130_fd_sc_hd__a311o_2 _16014_ (.A1(_11296_),
    .A2(_11990_),
    .A3(_11991_),
    .B1(_11992_),
    .C1(_11614_),
    .X(_11993_));
 sky130_fd_sc_hd__o2bb2a_2 _16015_ (.A1_N(\decode.regfile.registers_3[18] ),
    .A2_N(_11292_),
    .B1(_11367_),
    .B2(_10635_),
    .X(_11994_));
 sky130_fd_sc_hd__nand2_2 _16016_ (.A(_11993_),
    .B(_11994_),
    .Y(_11995_));
 sky130_fd_sc_hd__o221a_2 _16017_ (.A1(_11191_),
    .A2(_11097_),
    .B1(_11375_),
    .B2(\decode.regfile.registers_4[18] ),
    .C1(_11995_),
    .X(_11996_));
 sky130_fd_sc_hd__o32a_2 _16018_ (.A1(_10648_),
    .A2(_10624_),
    .A3(_11084_),
    .B1(_11989_),
    .B2(_11996_),
    .X(_11997_));
 sky130_fd_sc_hd__o31a_2 _16019_ (.A1(\decode.regfile.registers_8[18] ),
    .A2(_11280_),
    .A3(_11175_),
    .B1(_11131_),
    .X(_11998_));
 sky130_fd_sc_hd__o221a_2 _16020_ (.A1(\decode.regfile.registers_9[18] ),
    .A2(_11365_),
    .B1(_11988_),
    .B2(_11997_),
    .C1(_11998_),
    .X(_11999_));
 sky130_fd_sc_hd__o32a_2 _16021_ (.A1(\decode.regfile.registers_13[18] ),
    .A2(_11046_),
    .A3(_11690_),
    .B1(_11987_),
    .B2(_11999_),
    .X(_12000_));
 sky130_fd_sc_hd__o311a_2 _16022_ (.A1(\decode.regfile.registers_12[18] ),
    .A2(_10639_),
    .A3(_11690_),
    .B1(_11198_),
    .C1(_12000_),
    .X(_12001_));
 sky130_fd_sc_hd__o221a_2 _16023_ (.A1(\decode.regfile.registers_16[18] ),
    .A2(_11359_),
    .B1(_11986_),
    .B2(_12001_),
    .C1(_11126_),
    .X(_12002_));
 sky130_fd_sc_hd__a41o_2 _16024_ (.A1(\decode.regfile.registers_17[18] ),
    .A2(_10652_),
    .A3(_11112_),
    .A4(_11118_),
    .B1(_12002_),
    .X(_12003_));
 sky130_fd_sc_hd__o31a_2 _16025_ (.A1(_10955_),
    .A2(_11215_),
    .A3(_11216_),
    .B1(_12003_),
    .X(_12004_));
 sky130_fd_sc_hd__a211o_2 _16026_ (.A1(\decode.regfile.registers_18[18] ),
    .A2(_11455_),
    .B1(_11456_),
    .C1(_12004_),
    .X(_12005_));
 sky130_fd_sc_hd__o211a_2 _16027_ (.A1(\decode.regfile.registers_19[18] ),
    .A2(_11453_),
    .B1(_11454_),
    .C1(_12005_),
    .X(_12006_));
 sky130_fd_sc_hd__a211o_2 _16028_ (.A1(\decode.regfile.registers_20[18] ),
    .A2(_11452_),
    .B1(_11223_),
    .C1(_12006_),
    .X(_12007_));
 sky130_fd_sc_hd__o311a_2 _16029_ (.A1(\decode.regfile.registers_21[18] ),
    .A2(_11062_),
    .A3(_11100_),
    .B1(_11229_),
    .C1(_12007_),
    .X(_12008_));
 sky130_fd_sc_hd__o22a_2 _16030_ (.A1(\decode.regfile.registers_23[18] ),
    .A2(_11088_),
    .B1(_11985_),
    .B2(_12008_),
    .X(_12009_));
 sky130_fd_sc_hd__o22a_2 _16031_ (.A1(\decode.regfile.registers_25[18] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[18] ),
    .X(_12010_));
 sky130_fd_sc_hd__o211a_2 _16032_ (.A1(_11075_),
    .A2(_12009_),
    .B1(_12010_),
    .C1(_11486_),
    .X(_12011_));
 sky130_fd_sc_hd__o32a_2 _16033_ (.A1(_11251_),
    .A2(_11259_),
    .A3(\decode.regfile.registers_27[18] ),
    .B1(_11984_),
    .B2(_12011_),
    .X(_12012_));
 sky130_fd_sc_hd__o221a_2 _16034_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[18] ),
    .B1(\decode.regfile.registers_29[18] ),
    .B2(_11255_),
    .C1(_11245_),
    .X(_12013_));
 sky130_fd_sc_hd__o21a_2 _16035_ (.A1(_11445_),
    .A2(_12012_),
    .B1(_12013_),
    .X(_12014_));
 sky130_fd_sc_hd__o221a_2 _16036_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[18] ),
    .B1(_11983_),
    .B2(_12014_),
    .C1(_11760_),
    .X(_00406_));
 sky130_fd_sc_hd__o2111a_2 _16037_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[19] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_12015_));
 sky130_fd_sc_hd__o2111a_2 _16038_ (.A1(_11263_),
    .A2(\decode.regfile.registers_22[19] ),
    .B1(_11404_),
    .C1(_11264_),
    .D1(_11265_),
    .X(_12016_));
 sky130_fd_sc_hd__a221o_2 _16039_ (.A1(\decode.regfile.registers_14[19] ),
    .A2(_11360_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[19] ),
    .C1(_11202_),
    .X(_12017_));
 sky130_fd_sc_hd__and3_2 _16040_ (.A(_11036_),
    .B(_11058_),
    .C(_10632_),
    .X(_12018_));
 sky130_fd_sc_hd__a31o_2 _16041_ (.A1(\decode.regfile.registers_9[19] ),
    .A2(_11280_),
    .A3(_11134_),
    .B1(_11509_),
    .X(_12019_));
 sky130_fd_sc_hd__a31o_2 _16042_ (.A1(\decode.regfile.registers_7[19] ),
    .A2(_11092_),
    .A3(_11142_),
    .B1(_11166_),
    .X(_12020_));
 sky130_fd_sc_hd__a31o_2 _16043_ (.A1(\decode.regfile.registers_3[19] ),
    .A2(_11109_),
    .A3(_11141_),
    .B1(_11145_),
    .X(_12021_));
 sky130_fd_sc_hd__nand4_2 _16044_ (.A(\decode.regfile.registers_1[19] ),
    .B(_11116_),
    .C(_11137_),
    .D(_11157_),
    .Y(_12022_));
 sky130_fd_sc_hd__nand2_2 _16045_ (.A(_11300_),
    .B(\decode.regfile.registers_0[19] ),
    .Y(_12023_));
 sky130_fd_sc_hd__o211ai_2 _16046_ (.A1(_11298_),
    .A2(_10646_),
    .B1(_12022_),
    .C1(_12023_),
    .Y(_12024_));
 sky130_fd_sc_hd__o311a_2 _16047_ (.A1(\decode.regfile.registers_2[19] ),
    .A2(_10646_),
    .A3(_11298_),
    .B1(_11151_),
    .C1(_12024_),
    .X(_12025_));
 sky130_fd_sc_hd__o22ai_2 _16048_ (.A1(\decode.regfile.registers_4[19] ),
    .A2(_11375_),
    .B1(_12021_),
    .B2(_12025_),
    .Y(_12026_));
 sky130_fd_sc_hd__o2bb2a_2 _16049_ (.A1_N(\decode.regfile.registers_5[19] ),
    .A2_N(_11290_),
    .B1(_10636_),
    .B2(_11135_),
    .X(_12027_));
 sky130_fd_sc_hd__o21ai_2 _16050_ (.A1(_11291_),
    .A2(_12026_),
    .B1(_12027_),
    .Y(_12028_));
 sky130_fd_sc_hd__o221a_2 _16051_ (.A1(_11084_),
    .A2(_11297_),
    .B1(_11534_),
    .B2(\decode.regfile.registers_6[19] ),
    .C1(_12028_),
    .X(_12029_));
 sky130_fd_sc_hd__a21o_2 _16052_ (.A1(\decode.regfile.registers_8[19] ),
    .A2(_11044_),
    .B1(_11174_),
    .X(_12030_));
 sky130_fd_sc_hd__o21a_2 _16053_ (.A1(_12020_),
    .A2(_12029_),
    .B1(_12030_),
    .X(_12031_));
 sky130_fd_sc_hd__o32a_2 _16054_ (.A1(\decode.regfile.registers_10[19] ),
    .A2(_10638_),
    .A3(_11132_),
    .B1(_12019_),
    .B2(_12031_),
    .X(_12032_));
 sky130_fd_sc_hd__a31o_2 _16055_ (.A1(\decode.regfile.registers_11[19] ),
    .A2(_11071_),
    .A3(_11470_),
    .B1(_11278_),
    .X(_12033_));
 sky130_fd_sc_hd__a21oi_2 _16056_ (.A1(_12032_),
    .A2(_11364_),
    .B1(_12033_),
    .Y(_12034_));
 sky130_fd_sc_hd__a21oi_2 _16057_ (.A1(\decode.regfile.registers_12[19] ),
    .A2(_11047_),
    .B1(_11690_),
    .Y(_12035_));
 sky130_fd_sc_hd__o2bb2a_2 _16058_ (.A1_N(\decode.regfile.registers_13[19] ),
    .A2_N(_11276_),
    .B1(_12034_),
    .B2(_12035_),
    .X(_12036_));
 sky130_fd_sc_hd__nor2_2 _16059_ (.A(_12018_),
    .B(_12036_),
    .Y(_12037_));
 sky130_fd_sc_hd__o221a_2 _16060_ (.A1(\decode.regfile.registers_16[19] ),
    .A2(_11359_),
    .B1(_12017_),
    .B2(_12037_),
    .C1(_11127_),
    .X(_12038_));
 sky130_fd_sc_hd__a41o_2 _16061_ (.A1(\decode.regfile.registers_17[19] ),
    .A2(_10988_),
    .A3(_11113_),
    .A4(_11119_),
    .B1(_12038_),
    .X(_12039_));
 sky130_fd_sc_hd__o2111a_2 _16062_ (.A1(\decode.regfile.registers_18[19] ),
    .A2(_10955_),
    .B1(_11113_),
    .C1(_11094_),
    .D1(_10976_),
    .X(_12040_));
 sky130_fd_sc_hd__a21o_2 _16063_ (.A1(_11106_),
    .A2(_12039_),
    .B1(_12040_),
    .X(_12041_));
 sky130_fd_sc_hd__o41a_2 _16064_ (.A1(\decode.regfile.registers_19[19] ),
    .A2(_11048_),
    .A3(_11215_),
    .A4(_11216_),
    .B1(_11325_),
    .X(_12042_));
 sky130_fd_sc_hd__a221o_2 _16065_ (.A1(\decode.regfile.registers_20[19] ),
    .A2(_11102_),
    .B1(_12041_),
    .B2(_12042_),
    .C1(_11327_),
    .X(_12043_));
 sky130_fd_sc_hd__o311a_2 _16066_ (.A1(\decode.regfile.registers_21[19] ),
    .A2(_11267_),
    .A3(_11099_),
    .B1(_11228_),
    .C1(_12043_),
    .X(_12044_));
 sky130_fd_sc_hd__o22a_2 _16067_ (.A1(\decode.regfile.registers_23[19] ),
    .A2(_11087_),
    .B1(_12016_),
    .B2(_12044_),
    .X(_12045_));
 sky130_fd_sc_hd__a31o_2 _16068_ (.A1(_10992_),
    .A2(_11066_),
    .A3(_11261_),
    .B1(_12045_),
    .X(_12046_));
 sky130_fd_sc_hd__o22a_2 _16069_ (.A1(\decode.regfile.registers_25[19] ),
    .A2(_11333_),
    .B1(_11336_),
    .B2(\decode.regfile.registers_24[19] ),
    .X(_12047_));
 sky130_fd_sc_hd__o2111a_2 _16070_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[19] ),
    .B1(_11676_),
    .C1(_11338_),
    .D1(_11564_),
    .X(_12048_));
 sky130_fd_sc_hd__a31o_2 _16071_ (.A1(_11260_),
    .A2(_12046_),
    .A3(_12047_),
    .B1(_12048_),
    .X(_12049_));
 sky130_fd_sc_hd__or3_2 _16072_ (.A(_11679_),
    .B(\decode.regfile.registers_27[19] ),
    .C(_11869_),
    .X(_12050_));
 sky130_fd_sc_hd__o2111a_2 _16073_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[19] ),
    .B1(_11871_),
    .C1(_11681_),
    .D1(_11440_),
    .X(_12051_));
 sky130_fd_sc_hd__a31o_2 _16074_ (.A1(_11403_),
    .A2(_12049_),
    .A3(_12050_),
    .B1(_12051_),
    .X(_12052_));
 sky130_fd_sc_hd__o221a_2 _16075_ (.A1(_11646_),
    .A2(_11834_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[19] ),
    .C1(_12052_),
    .X(_12053_));
 sky130_fd_sc_hd__o221a_2 _16076_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[19] ),
    .B1(_12015_),
    .B2(_12053_),
    .C1(_11760_),
    .X(_00407_));
 sky130_fd_sc_hd__o2111a_2 _16077_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[20] ),
    .B1(_11722_),
    .C1(_11723_),
    .D1(_11724_),
    .X(_12054_));
 sky130_fd_sc_hd__a2bb2o_2 _16078_ (.A1_N(\decode.regfile.registers_23[20] ),
    .A2_N(_11087_),
    .B1(_11074_),
    .B2(_11049_),
    .X(_12055_));
 sky130_fd_sc_hd__or2_2 _16079_ (.A(\decode.regfile.registers_14[20] ),
    .B(_10639_),
    .X(_12056_));
 sky130_fd_sc_hd__a21oi_2 _16080_ (.A1(\decode.regfile.registers_10[20] ),
    .A2(_11184_),
    .B1(_11181_),
    .Y(_12057_));
 sky130_fd_sc_hd__a31o_2 _16081_ (.A1(\decode.regfile.registers_3[20] ),
    .A2(_11110_),
    .A3(_11142_),
    .B1(_11146_),
    .X(_12058_));
 sky130_fd_sc_hd__a31oi_2 _16082_ (.A1(_11117_),
    .A2(_11057_),
    .A3(_11109_),
    .B1(\decode.regfile.registers_0[20] ),
    .Y(_12059_));
 sky130_fd_sc_hd__and4b_2 _16083_ (.A_N(\decode.regfile.registers_1[20] ),
    .B(_11117_),
    .C(_11057_),
    .D(_11109_),
    .X(_12060_));
 sky130_fd_sc_hd__o21ai_2 _16084_ (.A1(_12059_),
    .A2(_12060_),
    .B1(_11369_),
    .Y(_12061_));
 sky130_fd_sc_hd__o311a_2 _16085_ (.A1(\decode.regfile.registers_2[20] ),
    .A2(_10647_),
    .A3(_11148_),
    .B1(_11152_),
    .C1(_12061_),
    .X(_12062_));
 sky130_fd_sc_hd__o22ai_2 _16086_ (.A1(\decode.regfile.registers_4[20] ),
    .A2(_11410_),
    .B1(_12058_),
    .B2(_12062_),
    .Y(_12063_));
 sky130_fd_sc_hd__o21ai_2 _16087_ (.A1(_11045_),
    .A2(_11410_),
    .B1(_12063_),
    .Y(_12064_));
 sky130_fd_sc_hd__or4_2 _16088_ (.A(_11503_),
    .B(_10629_),
    .C(_11043_),
    .D(_11083_),
    .X(_12065_));
 sky130_fd_sc_hd__o32a_2 _16089_ (.A1(_11192_),
    .A2(_11318_),
    .A3(_11084_),
    .B1(\decode.regfile.registers_5[20] ),
    .B2(_12065_),
    .X(_12066_));
 sky130_fd_sc_hd__a22oi_2 _16090_ (.A1(\decode.regfile.registers_6[20] ),
    .A2(_11170_),
    .B1(_12064_),
    .B2(_12066_),
    .Y(_12067_));
 sky130_fd_sc_hd__a21oi_2 _16091_ (.A1(\decode.regfile.registers_7[20] ),
    .A2(_11378_),
    .B1(_11134_),
    .Y(_12068_));
 sky130_fd_sc_hd__o21ai_2 _16092_ (.A1(_11378_),
    .A2(_12067_),
    .B1(_12068_),
    .Y(_12069_));
 sky130_fd_sc_hd__o221a_2 _16093_ (.A1(\decode.regfile.registers_8[20] ),
    .A2(_11285_),
    .B1(_11365_),
    .B2(\decode.regfile.registers_9[20] ),
    .C1(_11381_),
    .X(_12070_));
 sky130_fd_sc_hd__nand2_2 _16094_ (.A(_12069_),
    .B(_12070_),
    .Y(_12071_));
 sky130_fd_sc_hd__a2bb2o_2 _16095_ (.A1_N(\decode.regfile.registers_11[20] ),
    .A2_N(_11364_),
    .B1(_12057_),
    .B2(_12071_),
    .X(_12072_));
 sky130_fd_sc_hd__nand2_2 _16096_ (.A(_11690_),
    .B(_12072_),
    .Y(_12073_));
 sky130_fd_sc_hd__or4_2 _16097_ (.A(_10649_),
    .B(_10638_),
    .C(_11052_),
    .D(_10625_),
    .X(_12074_));
 sky130_fd_sc_hd__o221a_2 _16098_ (.A1(_11194_),
    .A2(\decode.regfile.registers_12[20] ),
    .B1(\decode.regfile.registers_13[20] ),
    .B2(_11196_),
    .C1(_12074_),
    .X(_12075_));
 sky130_fd_sc_hd__a22o_2 _16099_ (.A1(_12018_),
    .A2(_12056_),
    .B1(_12073_),
    .B2(_12075_),
    .X(_12076_));
 sky130_fd_sc_hd__o31a_2 _16100_ (.A1(\decode.regfile.registers_15[20] ),
    .A2(_11047_),
    .A3(_11199_),
    .B1(_11359_),
    .X(_12077_));
 sky130_fd_sc_hd__a22o_2 _16101_ (.A1(\decode.regfile.registers_16[20] ),
    .A2(_11203_),
    .B1(_12076_),
    .B2(_12077_),
    .X(_12078_));
 sky130_fd_sc_hd__mux2_2 _16102_ (.A0(_12078_),
    .A1(\decode.regfile.registers_17[20] ),
    .S(_11357_),
    .X(_12079_));
 sky130_fd_sc_hd__mux2_2 _16103_ (.A0(_12079_),
    .A1(\decode.regfile.registers_18[20] ),
    .S(_11455_),
    .X(_12080_));
 sky130_fd_sc_hd__a41o_2 _16104_ (.A1(_10989_),
    .A2(_10977_),
    .A3(_10956_),
    .A4(_11114_),
    .B1(_12080_),
    .X(_12081_));
 sky130_fd_sc_hd__o41a_2 _16105_ (.A1(\decode.regfile.registers_19[20] ),
    .A2(_11049_),
    .A3(_11215_),
    .A4(_11217_),
    .B1(_11454_),
    .X(_12082_));
 sky130_fd_sc_hd__a221o_2 _16106_ (.A1(\decode.regfile.registers_20[20] ),
    .A2(_11452_),
    .B1(_12081_),
    .B2(_12082_),
    .C1(_11223_),
    .X(_12083_));
 sky130_fd_sc_hd__o32a_2 _16107_ (.A1(_10957_),
    .A2(_11217_),
    .A3(_11085_),
    .B1(\decode.regfile.registers_21[20] ),
    .B2(_11648_),
    .X(_12084_));
 sky130_fd_sc_hd__a221oi_2 _16108_ (.A1(\decode.regfile.registers_22[20] ),
    .A2(_11096_),
    .B1(_12083_),
    .B2(_12084_),
    .C1(_11232_),
    .Y(_12085_));
 sky130_fd_sc_hd__o21ai_2 _16109_ (.A1(_10958_),
    .A2(\decode.regfile.registers_24[20] ),
    .B1(_11074_),
    .Y(_12086_));
 sky130_fd_sc_hd__o21ai_2 _16110_ (.A1(_12055_),
    .A2(_12085_),
    .B1(_12086_),
    .Y(_12087_));
 sky130_fd_sc_hd__or3_2 _16111_ (.A(_11050_),
    .B(\decode.regfile.registers_25[20] ),
    .C(_11089_),
    .X(_12088_));
 sky130_fd_sc_hd__o2111a_2 _16112_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[20] ),
    .B1(_11676_),
    .C1(_11338_),
    .D1(_11564_),
    .X(_12089_));
 sky130_fd_sc_hd__a31o_2 _16113_ (.A1(_11260_),
    .A2(_12087_),
    .A3(_12088_),
    .B1(_12089_),
    .X(_12090_));
 sky130_fd_sc_hd__or3_2 _16114_ (.A(_11679_),
    .B(\decode.regfile.registers_27[20] ),
    .C(_11869_),
    .X(_12091_));
 sky130_fd_sc_hd__o2111a_2 _16115_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[20] ),
    .B1(_11871_),
    .C1(_11681_),
    .D1(_11448_),
    .X(_12092_));
 sky130_fd_sc_hd__a31o_2 _16116_ (.A1(_11396_),
    .A2(_12090_),
    .A3(_12091_),
    .B1(_12092_),
    .X(_12093_));
 sky130_fd_sc_hd__o221a_2 _16117_ (.A1(_11646_),
    .A2(_11834_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[20] ),
    .C1(_12093_),
    .X(_12094_));
 sky130_fd_sc_hd__o221a_2 _16118_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[20] ),
    .B1(_12054_),
    .B2(_12094_),
    .C1(_11760_),
    .X(_00408_));
 sky130_fd_sc_hd__buf_1 _16119_ (.A(_11038_),
    .X(_12095_));
 sky130_fd_sc_hd__buf_1 _16120_ (.A(_10981_),
    .X(_12096_));
 sky130_fd_sc_hd__buf_1 _16121_ (.A(_10994_),
    .X(_12097_));
 sky130_fd_sc_hd__o2111a_2 _16122_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[21] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12098_));
 sky130_fd_sc_hd__o2111a_2 _16123_ (.A1(_11446_),
    .A2(\decode.regfile.registers_26[21] ),
    .B1(_11447_),
    .C1(_11348_),
    .D1(_10993_),
    .X(_12099_));
 sky130_fd_sc_hd__o2111a_2 _16124_ (.A1(_11493_),
    .A2(\decode.regfile.registers_22[21] ),
    .B1(_11450_),
    .C1(_10979_),
    .D1(_10991_),
    .X(_12100_));
 sky130_fd_sc_hd__a221o_2 _16125_ (.A1(\decode.regfile.registers_14[21] ),
    .A2(_11208_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[21] ),
    .C1(_11202_),
    .X(_12101_));
 sky130_fd_sc_hd__a31o_2 _16126_ (.A1(\decode.regfile.registers_11[21] ),
    .A2(_11071_),
    .A3(_11204_),
    .B1(_11407_),
    .X(_12102_));
 sky130_fd_sc_hd__a2bb2o_2 _16127_ (.A1_N(\decode.regfile.registers_2[21] ),
    .A2_N(_11369_),
    .B1(_11142_),
    .B2(_11110_),
    .X(_12103_));
 sky130_fd_sc_hd__a2bb2o_2 _16128_ (.A1_N(_11190_),
    .A2_N(_11148_),
    .B1(_11154_),
    .B2(\decode.regfile.registers_0[21] ),
    .X(_12104_));
 sky130_fd_sc_hd__a21oi_2 _16129_ (.A1(\decode.regfile.registers_1[21] ),
    .A2(_11539_),
    .B1(_12104_),
    .Y(_12105_));
 sky130_fd_sc_hd__o2bb2a_2 _16130_ (.A1_N(\decode.regfile.registers_3[21] ),
    .A2_N(_11614_),
    .B1(_11410_),
    .B2(_10636_),
    .X(_12106_));
 sky130_fd_sc_hd__o21ai_2 _16131_ (.A1(_12103_),
    .A2(_12105_),
    .B1(_12106_),
    .Y(_12107_));
 sky130_fd_sc_hd__a2111o_2 _16132_ (.A1(_11313_),
    .A2(\decode.regfile.registers_4[21] ),
    .B1(_11191_),
    .C1(_10630_),
    .D1(_11462_),
    .X(_12108_));
 sky130_fd_sc_hd__a22oi_2 _16133_ (.A1(\decode.regfile.registers_5[21] ),
    .A2(_11291_),
    .B1(_12107_),
    .B2(_12108_),
    .Y(_12109_));
 sky130_fd_sc_hd__a221oi_2 _16134_ (.A1(\decode.regfile.registers_7[21] ),
    .A2(_11378_),
    .B1(_11170_),
    .B2(\decode.regfile.registers_6[21] ),
    .C1(_11166_),
    .Y(_12110_));
 sky130_fd_sc_hd__o21ai_2 _16135_ (.A1(_11289_),
    .A2(_12109_),
    .B1(_12110_),
    .Y(_12111_));
 sky130_fd_sc_hd__a21o_2 _16136_ (.A1(\decode.regfile.registers_8[21] ),
    .A2(_11045_),
    .B1(_11175_),
    .X(_12112_));
 sky130_fd_sc_hd__a221o_2 _16137_ (.A1(\decode.regfile.registers_9[21] ),
    .A2(_11547_),
    .B1(_12111_),
    .B2(_12112_),
    .C1(_11509_),
    .X(_12113_));
 sky130_fd_sc_hd__o211a_2 _16138_ (.A1(_11382_),
    .A2(\decode.regfile.registers_10[21] ),
    .B1(_11364_),
    .C1(_12113_),
    .X(_12114_));
 sky130_fd_sc_hd__a2111o_2 _16139_ (.A1(_11046_),
    .A2(\decode.regfile.registers_12[21] ),
    .B1(_10650_),
    .C1(_11052_),
    .D1(_10632_),
    .X(_12115_));
 sky130_fd_sc_hd__o21ai_2 _16140_ (.A1(_12102_),
    .A2(_12114_),
    .B1(_12115_),
    .Y(_12116_));
 sky130_fd_sc_hd__nand2_2 _16141_ (.A(\decode.regfile.registers_13[21] ),
    .B(_11276_),
    .Y(_12117_));
 sky130_fd_sc_hd__o2bb2a_2 _16142_ (.A1_N(_12116_),
    .A2_N(_12117_),
    .B1(_11054_),
    .B2(_11318_),
    .X(_12118_));
 sky130_fd_sc_hd__o22a_2 _16143_ (.A1(\decode.regfile.registers_16[21] ),
    .A2(_11124_),
    .B1(_12101_),
    .B2(_12118_),
    .X(_12119_));
 sky130_fd_sc_hd__a31o_2 _16144_ (.A1(_10988_),
    .A2(_11113_),
    .A3(_11119_),
    .B1(_12119_),
    .X(_12120_));
 sky130_fd_sc_hd__o32a_2 _16145_ (.A1(_11225_),
    .A2(_11125_),
    .A3(_11216_),
    .B1(\decode.regfile.registers_17[21] ),
    .B2(_11128_),
    .X(_12121_));
 sky130_fd_sc_hd__a221o_2 _16146_ (.A1(\decode.regfile.registers_18[21] ),
    .A2(_11455_),
    .B1(_12120_),
    .B2(_12121_),
    .C1(_11456_),
    .X(_12122_));
 sky130_fd_sc_hd__o211a_2 _16147_ (.A1(\decode.regfile.registers_19[21] ),
    .A2(_11453_),
    .B1(_11454_),
    .C1(_12122_),
    .X(_12123_));
 sky130_fd_sc_hd__a211o_2 _16148_ (.A1(\decode.regfile.registers_20[21] ),
    .A2(_11452_),
    .B1(_11223_),
    .C1(_12123_),
    .X(_12124_));
 sky130_fd_sc_hd__o311a_2 _16149_ (.A1(\decode.regfile.registers_21[21] ),
    .A2(_11061_),
    .A3(_11100_),
    .B1(_11229_),
    .C1(_12124_),
    .X(_12125_));
 sky130_fd_sc_hd__o22a_2 _16150_ (.A1(\decode.regfile.registers_23[21] ),
    .A2(_11088_),
    .B1(_12100_),
    .B2(_12125_),
    .X(_12126_));
 sky130_fd_sc_hd__o22a_2 _16151_ (.A1(\decode.regfile.registers_25[21] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[21] ),
    .X(_12127_));
 sky130_fd_sc_hd__o211a_2 _16152_ (.A1(_11075_),
    .A2(_12126_),
    .B1(_12127_),
    .C1(_11486_),
    .X(_12128_));
 sky130_fd_sc_hd__o32a_2 _16153_ (.A1(_11251_),
    .A2(_11259_),
    .A3(\decode.regfile.registers_27[21] ),
    .B1(_12099_),
    .B2(_12128_),
    .X(_12129_));
 sky130_fd_sc_hd__o221a_2 _16154_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[21] ),
    .B1(\decode.regfile.registers_29[21] ),
    .B2(_11063_),
    .C1(_11245_),
    .X(_12130_));
 sky130_fd_sc_hd__o21a_2 _16155_ (.A1(_11445_),
    .A2(_12129_),
    .B1(_12130_),
    .X(_12131_));
 sky130_fd_sc_hd__buf_1 _16156_ (.A(_11248_),
    .X(_12132_));
 sky130_fd_sc_hd__o221a_2 _16157_ (.A1(_11761_),
    .A2(\decode.regfile.registers_31[21] ),
    .B1(_12098_),
    .B2(_12131_),
    .C1(_12132_),
    .X(_00409_));
 sky130_fd_sc_hd__buf_1 _16158_ (.A(_11243_),
    .X(_12133_));
 sky130_fd_sc_hd__o2111a_2 _16159_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[22] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12134_));
 sky130_fd_sc_hd__o2111a_2 _16160_ (.A1(_10959_),
    .A2(\decode.regfile.registers_26[22] ),
    .B1(_11447_),
    .C1(_11348_),
    .D1(_10993_),
    .X(_12135_));
 sky130_fd_sc_hd__o2111a_2 _16161_ (.A1(_10957_),
    .A2(\decode.regfile.registers_22[22] ),
    .B1(_11450_),
    .C1(_10978_),
    .D1(_10990_),
    .X(_12136_));
 sky130_fd_sc_hd__o21ai_2 _16162_ (.A1(\decode.regfile.registers_17[22] ),
    .A2(_11128_),
    .B1(_11106_),
    .Y(_12137_));
 sky130_fd_sc_hd__inv_2 _16163_ (.A(\decode.regfile.registers_1[22] ),
    .Y(_12138_));
 sky130_fd_sc_hd__nand2_2 _16164_ (.A(_11371_),
    .B(\decode.regfile.registers_0[22] ),
    .Y(_12139_));
 sky130_fd_sc_hd__o221ai_2 _16165_ (.A1(_12138_),
    .A2(_11154_),
    .B1(_11190_),
    .B2(_11148_),
    .C1(_12139_),
    .Y(_12140_));
 sky130_fd_sc_hd__o32a_2 _16166_ (.A1(_10659_),
    .A2(_10654_),
    .A3(_11150_),
    .B1(\decode.regfile.registers_2[22] ),
    .B2(_11296_),
    .X(_12141_));
 sky130_fd_sc_hd__a221o_2 _16167_ (.A1(\decode.regfile.registers_3[22] ),
    .A2(_11614_),
    .B1(_12140_),
    .B2(_12141_),
    .C1(_11146_),
    .X(_12142_));
 sky130_fd_sc_hd__a2111o_2 _16168_ (.A1(_11313_),
    .A2(\decode.regfile.registers_4[22] ),
    .B1(_10647_),
    .C1(_10629_),
    .D1(_11462_),
    .X(_12143_));
 sky130_fd_sc_hd__a32o_2 _16169_ (.A1(\decode.regfile.registers_5[22] ),
    .A2(_10637_),
    .A3(_11139_),
    .B1(_12142_),
    .B2(_12143_),
    .X(_12144_));
 sky130_fd_sc_hd__a221o_2 _16170_ (.A1(\decode.regfile.registers_7[22] ),
    .A2(_11465_),
    .B1(_11466_),
    .B2(\decode.regfile.registers_6[22] ),
    .C1(_11166_),
    .X(_12145_));
 sky130_fd_sc_hd__a21o_2 _16171_ (.A1(_11136_),
    .A2(_12144_),
    .B1(_12145_),
    .X(_12146_));
 sky130_fd_sc_hd__a21o_2 _16172_ (.A1(\decode.regfile.registers_8[22] ),
    .A2(_11045_),
    .B1(_11175_),
    .X(_12147_));
 sky130_fd_sc_hd__a31o_2 _16173_ (.A1(\decode.regfile.registers_9[22] ),
    .A2(_11280_),
    .A3(_11134_),
    .B1(_11509_),
    .X(_12148_));
 sky130_fd_sc_hd__a21o_2 _16174_ (.A1(_12146_),
    .A2(_12147_),
    .B1(_12148_),
    .X(_12149_));
 sky130_fd_sc_hd__o211a_2 _16175_ (.A1(_11382_),
    .A2(\decode.regfile.registers_10[22] ),
    .B1(_11364_),
    .C1(_12149_),
    .X(_12150_));
 sky130_fd_sc_hd__a311o_2 _16176_ (.A1(\decode.regfile.registers_11[22] ),
    .A2(_11072_),
    .A3(_11204_),
    .B1(_11407_),
    .C1(_12150_),
    .X(_12151_));
 sky130_fd_sc_hd__a2111o_2 _16177_ (.A1(_11047_),
    .A2(\decode.regfile.registers_12[22] ),
    .B1(_10650_),
    .C1(_11053_),
    .D1(_10632_),
    .X(_12152_));
 sky130_fd_sc_hd__a32o_2 _16178_ (.A1(\decode.regfile.registers_13[22] ),
    .A2(_10642_),
    .A3(_11187_),
    .B1(_12151_),
    .B2(_12152_),
    .X(_12153_));
 sky130_fd_sc_hd__and3_2 _16179_ (.A(\decode.regfile.registers_15[22] ),
    .B(_11036_),
    .C(_11205_),
    .X(_12154_));
 sky130_fd_sc_hd__a221o_2 _16180_ (.A1(\decode.regfile.registers_14[22] ),
    .A2(_11208_),
    .B1(_12153_),
    .B2(_11199_),
    .C1(_12154_),
    .X(_12155_));
 sky130_fd_sc_hd__a32o_2 _16181_ (.A1(_10988_),
    .A2(_11113_),
    .A3(_11119_),
    .B1(_11203_),
    .B2(\decode.regfile.registers_16[22] ),
    .X(_12156_));
 sky130_fd_sc_hd__a21oi_2 _16182_ (.A1(_11124_),
    .A2(_12155_),
    .B1(_12156_),
    .Y(_12157_));
 sky130_fd_sc_hd__a21oi_2 _16183_ (.A1(\decode.regfile.registers_18[22] ),
    .A2(_11455_),
    .B1(_11456_),
    .Y(_12158_));
 sky130_fd_sc_hd__o21ai_2 _16184_ (.A1(_12137_),
    .A2(_12157_),
    .B1(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__o211a_2 _16185_ (.A1(\decode.regfile.registers_19[22] ),
    .A2(_11453_),
    .B1(_11219_),
    .C1(_12159_),
    .X(_12160_));
 sky130_fd_sc_hd__a211o_2 _16186_ (.A1(\decode.regfile.registers_20[22] ),
    .A2(_11103_),
    .B1(_11222_),
    .C1(_12160_),
    .X(_12161_));
 sky130_fd_sc_hd__o311a_2 _16187_ (.A1(\decode.regfile.registers_21[22] ),
    .A2(_11061_),
    .A3(_11099_),
    .B1(_11229_),
    .C1(_12161_),
    .X(_12162_));
 sky130_fd_sc_hd__o22a_2 _16188_ (.A1(\decode.regfile.registers_23[22] ),
    .A2(_11087_),
    .B1(_12136_),
    .B2(_12162_),
    .X(_12163_));
 sky130_fd_sc_hd__o22a_2 _16189_ (.A1(\decode.regfile.registers_25[22] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[22] ),
    .X(_12164_));
 sky130_fd_sc_hd__o211a_2 _16190_ (.A1(_11075_),
    .A2(_12163_),
    .B1(_12164_),
    .C1(_11236_),
    .X(_12165_));
 sky130_fd_sc_hd__o32a_2 _16191_ (.A1(_11250_),
    .A2(_11258_),
    .A3(\decode.regfile.registers_27[22] ),
    .B1(_12135_),
    .B2(_12165_),
    .X(_12166_));
 sky130_fd_sc_hd__o22a_2 _16192_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[22] ),
    .B1(\decode.regfile.registers_29[22] ),
    .B2(_11255_),
    .X(_12167_));
 sky130_fd_sc_hd__o211a_2 _16193_ (.A1(_11445_),
    .A2(_12166_),
    .B1(_12167_),
    .C1(_11246_),
    .X(_12168_));
 sky130_fd_sc_hd__o221a_2 _16194_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[22] ),
    .B1(_12134_),
    .B2(_12168_),
    .C1(_12132_),
    .X(_00410_));
 sky130_fd_sc_hd__o2111a_2 _16195_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[23] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12169_));
 sky130_fd_sc_hd__o2111a_2 _16196_ (.A1(_10959_),
    .A2(\decode.regfile.registers_26[23] ),
    .B1(_11349_),
    .C1(_11348_),
    .D1(_10993_),
    .X(_12170_));
 sky130_fd_sc_hd__o2111a_2 _16197_ (.A1(_10957_),
    .A2(\decode.regfile.registers_22[23] ),
    .B1(_11450_),
    .C1(_10978_),
    .D1(_10990_),
    .X(_12171_));
 sky130_fd_sc_hd__a221o_2 _16198_ (.A1(\decode.regfile.registers_14[23] ),
    .A2(_11360_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[23] ),
    .C1(_11202_),
    .X(_12172_));
 sky130_fd_sc_hd__a31o_2 _16199_ (.A1(\decode.regfile.registers_11[23] ),
    .A2(_11071_),
    .A3(_11204_),
    .B1(_11187_),
    .X(_12173_));
 sky130_fd_sc_hd__a31o_2 _16200_ (.A1(\decode.regfile.registers_5[23] ),
    .A2(_10637_),
    .A3(_11139_),
    .B1(_11170_),
    .X(_12174_));
 sky130_fd_sc_hd__a31o_2 _16201_ (.A1(\decode.regfile.registers_3[23] ),
    .A2(_11111_),
    .A3(_11142_),
    .B1(_11146_),
    .X(_12175_));
 sky130_fd_sc_hd__and4_2 _16202_ (.A(\decode.regfile.registers_1[23] ),
    .B(_11117_),
    .C(_11057_),
    .D(_11109_),
    .X(_12176_));
 sky130_fd_sc_hd__a211o_2 _16203_ (.A1(_11154_),
    .A2(\decode.regfile.registers_0[23] ),
    .B1(_11156_),
    .C1(_12176_),
    .X(_12177_));
 sky130_fd_sc_hd__o311a_2 _16204_ (.A1(\decode.regfile.registers_2[23] ),
    .A2(_11191_),
    .A3(_11149_),
    .B1(_11152_),
    .C1(_12177_),
    .X(_12178_));
 sky130_fd_sc_hd__a2111o_2 _16205_ (.A1(_11044_),
    .A2(\decode.regfile.registers_4[23] ),
    .B1(_11191_),
    .C1(_10630_),
    .D1(_11084_),
    .X(_12179_));
 sky130_fd_sc_hd__o21a_2 _16206_ (.A1(_12175_),
    .A2(_12178_),
    .B1(_12179_),
    .X(_12180_));
 sky130_fd_sc_hd__o32a_2 _16207_ (.A1(\decode.regfile.registers_6[23] ),
    .A2(_10638_),
    .A3(_11136_),
    .B1(_12174_),
    .B2(_12180_),
    .X(_12181_));
 sky130_fd_sc_hd__a31o_2 _16208_ (.A1(\decode.regfile.registers_7[23] ),
    .A2(_11092_),
    .A3(_11167_),
    .B1(_11134_),
    .X(_12182_));
 sky130_fd_sc_hd__a21o_2 _16209_ (.A1(_12181_),
    .A2(_11533_),
    .B1(_12182_),
    .X(_12183_));
 sky130_fd_sc_hd__o221a_2 _16210_ (.A1(\decode.regfile.registers_8[23] ),
    .A2(_11285_),
    .B1(_11365_),
    .B2(\decode.regfile.registers_9[23] ),
    .C1(_11382_),
    .X(_12184_));
 sky130_fd_sc_hd__a22oi_2 _16211_ (.A1(\decode.regfile.registers_10[23] ),
    .A2(_11184_),
    .B1(_12183_),
    .B2(_12184_),
    .Y(_12185_));
 sky130_fd_sc_hd__a21oi_2 _16212_ (.A1(_11072_),
    .A2(_11205_),
    .B1(_12185_),
    .Y(_12186_));
 sky130_fd_sc_hd__o221a_2 _16213_ (.A1(_11194_),
    .A2(\decode.regfile.registers_12[23] ),
    .B1(\decode.regfile.registers_13[23] ),
    .B2(_11196_),
    .C1(_11198_),
    .X(_12187_));
 sky130_fd_sc_hd__o21a_2 _16214_ (.A1(_12173_),
    .A2(_12186_),
    .B1(_12187_),
    .X(_12188_));
 sky130_fd_sc_hd__o22a_2 _16215_ (.A1(\decode.regfile.registers_16[23] ),
    .A2(_11359_),
    .B1(_12172_),
    .B2(_12188_),
    .X(_12189_));
 sky130_fd_sc_hd__mux2_2 _16216_ (.A0(_12189_),
    .A1(\decode.regfile.registers_17[23] ),
    .S(_11357_),
    .X(_12190_));
 sky130_fd_sc_hd__o2111a_2 _16217_ (.A1(\decode.regfile.registers_18[23] ),
    .A2(_10955_),
    .B1(_11114_),
    .C1(_11094_),
    .D1(_10976_),
    .X(_12191_));
 sky130_fd_sc_hd__a21o_2 _16218_ (.A1(_11106_),
    .A2(_12190_),
    .B1(_12191_),
    .X(_12192_));
 sky130_fd_sc_hd__o211a_2 _16219_ (.A1(\decode.regfile.registers_19[23] ),
    .A2(_11453_),
    .B1(_11219_),
    .C1(_12192_),
    .X(_12193_));
 sky130_fd_sc_hd__a211o_2 _16220_ (.A1(\decode.regfile.registers_20[23] ),
    .A2(_11103_),
    .B1(_11222_),
    .C1(_12193_),
    .X(_12194_));
 sky130_fd_sc_hd__o311a_2 _16221_ (.A1(\decode.regfile.registers_21[23] ),
    .A2(_11061_),
    .A3(_11099_),
    .B1(_11228_),
    .C1(_12194_),
    .X(_12195_));
 sky130_fd_sc_hd__o22a_2 _16222_ (.A1(\decode.regfile.registers_23[23] ),
    .A2(_11087_),
    .B1(_12171_),
    .B2(_12195_),
    .X(_12196_));
 sky130_fd_sc_hd__o22a_2 _16223_ (.A1(\decode.regfile.registers_25[23] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[23] ),
    .X(_12197_));
 sky130_fd_sc_hd__o211a_2 _16224_ (.A1(_11074_),
    .A2(_12196_),
    .B1(_12197_),
    .C1(_11236_),
    .X(_12198_));
 sky130_fd_sc_hd__o32a_2 _16225_ (.A1(_11250_),
    .A2(_11258_),
    .A3(\decode.regfile.registers_27[23] ),
    .B1(_12170_),
    .B2(_12198_),
    .X(_12199_));
 sky130_fd_sc_hd__o22a_2 _16226_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[23] ),
    .B1(\decode.regfile.registers_29[23] ),
    .B2(_11255_),
    .X(_12200_));
 sky130_fd_sc_hd__o211a_2 _16227_ (.A1(_11398_),
    .A2(_12199_),
    .B1(_12200_),
    .C1(_11246_),
    .X(_12201_));
 sky130_fd_sc_hd__o221a_2 _16228_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[23] ),
    .B1(_12169_),
    .B2(_12201_),
    .C1(_12132_),
    .X(_00411_));
 sky130_fd_sc_hd__o2111a_2 _16229_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[24] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12202_));
 sky130_fd_sc_hd__o2111a_2 _16230_ (.A1(_11435_),
    .A2(\decode.regfile.registers_24[24] ),
    .B1(_11244_),
    .C1(_11080_),
    .D1(_11079_),
    .X(_12203_));
 sky130_fd_sc_hd__o2111a_2 _16231_ (.A1(_11263_),
    .A2(\decode.regfile.registers_22[24] ),
    .B1(_11404_),
    .C1(_11264_),
    .D1(_11265_),
    .X(_12204_));
 sky130_fd_sc_hd__a221o_2 _16232_ (.A1(\decode.regfile.registers_14[24] ),
    .A2(_11207_),
    .B1(_11273_),
    .B2(\decode.regfile.registers_15[24] ),
    .C1(_11361_),
    .X(_12205_));
 sky130_fd_sc_hd__or4_2 _16233_ (.A(\decode.regfile.registers_12[24] ),
    .B(_10648_),
    .C(_10631_),
    .D(_11051_),
    .X(_12206_));
 sky130_fd_sc_hd__a32o_2 _16234_ (.A1(\decode.regfile.registers_7[24] ),
    .A2(_11092_),
    .A3(_11142_),
    .B1(_11169_),
    .B2(\decode.regfile.registers_6[24] ),
    .X(_12207_));
 sky130_fd_sc_hd__o2bb2a_2 _16235_ (.A1_N(\decode.regfile.registers_3[24] ),
    .A2_N(_11614_),
    .B1(_11367_),
    .B2(_11178_),
    .X(_12208_));
 sky130_fd_sc_hd__mux2_2 _16236_ (.A0(\decode.regfile.registers_1[24] ),
    .A1(\decode.regfile.registers_0[24] ),
    .S(_11371_),
    .X(_12209_));
 sky130_fd_sc_hd__o32a_2 _16237_ (.A1(_10660_),
    .A2(_10655_),
    .A3(_11150_),
    .B1(\decode.regfile.registers_2[24] ),
    .B2(_11296_),
    .X(_12210_));
 sky130_fd_sc_hd__o21ai_2 _16238_ (.A1(_11156_),
    .A2(_12209_),
    .B1(_12210_),
    .Y(_12211_));
 sky130_fd_sc_hd__a2bb2oi_2 _16239_ (.A1_N(\decode.regfile.registers_4[24] ),
    .A2_N(_11410_),
    .B1(_12208_),
    .B2(_12211_),
    .Y(_12212_));
 sky130_fd_sc_hd__o32a_2 _16240_ (.A1(\decode.regfile.registers_5[24] ),
    .A2(_11313_),
    .A3(_11410_),
    .B1(_11462_),
    .B2(_11314_),
    .X(_12213_));
 sky130_fd_sc_hd__o21ai_2 _16241_ (.A1(_11291_),
    .A2(_12212_),
    .B1(_12213_),
    .Y(_12214_));
 sky130_fd_sc_hd__nand3b_2 _16242_ (.A_N(_12207_),
    .B(_12214_),
    .C(_11175_),
    .Y(_12215_));
 sky130_fd_sc_hd__o221a_2 _16243_ (.A1(\decode.regfile.registers_8[24] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(\decode.regfile.registers_9[24] ),
    .C1(_11381_),
    .X(_12216_));
 sky130_fd_sc_hd__a22oi_2 _16244_ (.A1(\decode.regfile.registers_10[24] ),
    .A2(_11183_),
    .B1(_12215_),
    .B2(_12216_),
    .Y(_12217_));
 sky130_fd_sc_hd__o2bb2a_2 _16245_ (.A1_N(\decode.regfile.registers_11[24] ),
    .A2_N(_11180_),
    .B1(_11689_),
    .B2(_11280_),
    .X(_12218_));
 sky130_fd_sc_hd__o21ai_2 _16246_ (.A1(_11181_),
    .A2(_12217_),
    .B1(_12218_),
    .Y(_12219_));
 sky130_fd_sc_hd__a32o_2 _16247_ (.A1(_10639_),
    .A2(_11143_),
    .A3(_11036_),
    .B1(_12206_),
    .B2(_12219_),
    .X(_12220_));
 sky130_fd_sc_hd__o311a_2 _16248_ (.A1(\decode.regfile.registers_13[24] ),
    .A2(_11047_),
    .A3(_11690_),
    .B1(_11198_),
    .C1(_12220_),
    .X(_12221_));
 sky130_fd_sc_hd__o22a_2 _16249_ (.A1(\decode.regfile.registers_16[24] ),
    .A2(_11123_),
    .B1(_12205_),
    .B2(_12221_),
    .X(_12222_));
 sky130_fd_sc_hd__mux2_2 _16250_ (.A0(_12222_),
    .A1(\decode.regfile.registers_17[24] ),
    .S(_11357_),
    .X(_12223_));
 sky130_fd_sc_hd__o2111a_2 _16251_ (.A1(\decode.regfile.registers_18[24] ),
    .A2(_10642_),
    .B1(_11112_),
    .C1(_10988_),
    .D1(_10976_),
    .X(_12224_));
 sky130_fd_sc_hd__a21o_2 _16252_ (.A1(_11106_),
    .A2(_12223_),
    .B1(_12224_),
    .X(_12225_));
 sky130_fd_sc_hd__o211a_2 _16253_ (.A1(\decode.regfile.registers_19[24] ),
    .A2(_11406_),
    .B1(_11325_),
    .C1(_12225_),
    .X(_12226_));
 sky130_fd_sc_hd__a211o_2 _16254_ (.A1(\decode.regfile.registers_20[24] ),
    .A2(_11102_),
    .B1(_11327_),
    .C1(_12226_),
    .X(_12227_));
 sky130_fd_sc_hd__o311a_2 _16255_ (.A1(\decode.regfile.registers_21[24] ),
    .A2(_11267_),
    .A3(_11098_),
    .B1(_11227_),
    .C1(_12227_),
    .X(_12228_));
 sky130_fd_sc_hd__o221a_2 _16256_ (.A1(\decode.regfile.registers_23[24] ),
    .A2(_11262_),
    .B1(_12204_),
    .B2(_12228_),
    .C1(_11335_),
    .X(_12229_));
 sky130_fd_sc_hd__o32a_2 _16257_ (.A1(_11076_),
    .A2(_11090_),
    .A3(\decode.regfile.registers_25[24] ),
    .B1(_12203_),
    .B2(_12229_),
    .X(_12230_));
 sky130_fd_sc_hd__o2111a_2 _16258_ (.A1(_10959_),
    .A2(\decode.regfile.registers_26[24] ),
    .B1(_11349_),
    .C1(_10980_),
    .D1(_11347_),
    .X(_12231_));
 sky130_fd_sc_hd__a21o_2 _16259_ (.A1(_12230_),
    .A2(_11486_),
    .B1(_12231_),
    .X(_12232_));
 sky130_fd_sc_hd__or3_2 _16260_ (.A(_11679_),
    .B(\decode.regfile.registers_27[24] ),
    .C(_11869_),
    .X(_12233_));
 sky130_fd_sc_hd__o2111a_2 _16261_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[24] ),
    .B1(_11871_),
    .C1(_11681_),
    .D1(_11448_),
    .X(_12234_));
 sky130_fd_sc_hd__a31o_2 _16262_ (.A1(_11396_),
    .A2(_12232_),
    .A3(_12233_),
    .B1(_12234_),
    .X(_12235_));
 sky130_fd_sc_hd__o221a_2 _16263_ (.A1(_11646_),
    .A2(_11834_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[24] ),
    .C1(_12235_),
    .X(_12236_));
 sky130_fd_sc_hd__o221a_2 _16264_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[24] ),
    .B1(_12202_),
    .B2(_12236_),
    .C1(_12132_),
    .X(_00412_));
 sky130_fd_sc_hd__o2111a_2 _16265_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[25] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12237_));
 sky130_fd_sc_hd__or2_2 _16266_ (.A(_11493_),
    .B(\decode.regfile.registers_24[25] ),
    .X(_12238_));
 sky130_fd_sc_hd__a221o_2 _16267_ (.A1(\decode.regfile.registers_14[25] ),
    .A2(_11206_),
    .B1(_11272_),
    .B2(\decode.regfile.registers_15[25] ),
    .C1(_11201_),
    .X(_12239_));
 sky130_fd_sc_hd__a22o_2 _16268_ (.A1(\decode.regfile.registers_13[25] ),
    .A2(_11275_),
    .B1(_11278_),
    .B2(\decode.regfile.registers_12[25] ),
    .X(_12240_));
 sky130_fd_sc_hd__and4b_2 _16269_ (.A_N(\decode.regfile.registers_5[25] ),
    .B(_11117_),
    .C(_11092_),
    .D(_11058_),
    .X(_12241_));
 sky130_fd_sc_hd__nor2_2 _16270_ (.A(\decode.regfile.registers_1[25] ),
    .B(_11300_),
    .Y(_12242_));
 sky130_fd_sc_hd__o21bai_2 _16271_ (.A1(\decode.regfile.registers_0[25] ),
    .A2(_11539_),
    .B1_N(_12242_),
    .Y(_12243_));
 sky130_fd_sc_hd__o2bb2a_2 _16272_ (.A1_N(\decode.regfile.registers_2[25] ),
    .A2_N(_11156_),
    .B1(_11150_),
    .B2(_11120_),
    .X(_12244_));
 sky130_fd_sc_hd__o21ai_2 _16273_ (.A1(_11156_),
    .A2(_12243_),
    .B1(_12244_),
    .Y(_12245_));
 sky130_fd_sc_hd__o32a_2 _16274_ (.A1(_11150_),
    .A2(\decode.regfile.registers_3[25] ),
    .A3(_11121_),
    .B1(_11178_),
    .B2(_11367_),
    .X(_12246_));
 sky130_fd_sc_hd__o211a_2 _16275_ (.A1(\decode.regfile.registers_4[25] ),
    .A2(_11178_),
    .B1(_11143_),
    .C1(_11091_),
    .X(_12247_));
 sky130_fd_sc_hd__a21oi_2 _16276_ (.A1(_12245_),
    .A2(_12246_),
    .B1(_12247_),
    .Y(_12248_));
 sky130_fd_sc_hd__o21ai_2 _16277_ (.A1(_12241_),
    .A2(_12248_),
    .B1(_11135_),
    .Y(_12249_));
 sky130_fd_sc_hd__o32a_2 _16278_ (.A1(\decode.regfile.registers_7[25] ),
    .A2(_11462_),
    .A3(_11297_),
    .B1(\decode.regfile.registers_6[25] ),
    .B2(_11534_),
    .X(_12250_));
 sky130_fd_sc_hd__a221o_2 _16279_ (.A1(\decode.regfile.registers_8[25] ),
    .A2(_11165_),
    .B1(_11547_),
    .B2(\decode.regfile.registers_9[25] ),
    .C1(_11182_),
    .X(_12251_));
 sky130_fd_sc_hd__a31o_2 _16280_ (.A1(_11174_),
    .A2(_12249_),
    .A3(_12250_),
    .B1(_12251_),
    .X(_12252_));
 sky130_fd_sc_hd__o31a_2 _16281_ (.A1(\decode.regfile.registers_10[25] ),
    .A2(_10637_),
    .A3(_11131_),
    .B1(_11315_),
    .X(_12253_));
 sky130_fd_sc_hd__a22oi_2 _16282_ (.A1(\decode.regfile.registers_11[25] ),
    .A2(_11180_),
    .B1(_12252_),
    .B2(_12253_),
    .Y(_12254_));
 sky130_fd_sc_hd__a21oi_2 _16283_ (.A1(_11143_),
    .A2(_11035_),
    .B1(_12254_),
    .Y(_12255_));
 sky130_fd_sc_hd__o32a_2 _16284_ (.A1(_10649_),
    .A2(_10625_),
    .A3(_11052_),
    .B1(_12240_),
    .B2(_12255_),
    .X(_12256_));
 sky130_fd_sc_hd__o22a_2 _16285_ (.A1(\decode.regfile.registers_16[25] ),
    .A2(_11122_),
    .B1(_12239_),
    .B2(_12256_),
    .X(_12257_));
 sky130_fd_sc_hd__mux2_2 _16286_ (.A0(_12257_),
    .A1(\decode.regfile.registers_17[25] ),
    .S(_11356_),
    .X(_12258_));
 sky130_fd_sc_hd__o2111a_2 _16287_ (.A1(\decode.regfile.registers_18[25] ),
    .A2(_10640_),
    .B1(_11112_),
    .C1(_10651_),
    .D1(_10633_),
    .X(_12259_));
 sky130_fd_sc_hd__a21o_2 _16288_ (.A1(_11105_),
    .A2(_12258_),
    .B1(_12259_),
    .X(_12260_));
 sky130_fd_sc_hd__o211a_2 _16289_ (.A1(\decode.regfile.registers_19[25] ),
    .A2(_11354_),
    .B1(_11218_),
    .C1(_12260_),
    .X(_12261_));
 sky130_fd_sc_hd__a211o_2 _16290_ (.A1(\decode.regfile.registers_20[25] ),
    .A2(_11101_),
    .B1(_11221_),
    .C1(_12261_),
    .X(_12262_));
 sky130_fd_sc_hd__o311a_2 _16291_ (.A1(\decode.regfile.registers_21[25] ),
    .A2(_11060_),
    .A3(_11098_),
    .B1(_11227_),
    .C1(_12262_),
    .X(_12263_));
 sky130_fd_sc_hd__a211o_2 _16292_ (.A1(\decode.regfile.registers_22[25] ),
    .A2(_11096_),
    .B1(_11232_),
    .C1(_12263_),
    .X(_12264_));
 sky130_fd_sc_hd__o221a_2 _16293_ (.A1(\decode.regfile.registers_23[25] ),
    .A2(_11262_),
    .B1(_11089_),
    .B2(_11493_),
    .C1(_12264_),
    .X(_12265_));
 sky130_fd_sc_hd__a41o_2 _16294_ (.A1(_11079_),
    .A2(_11244_),
    .A3(_11080_),
    .A4(_12238_),
    .B1(_12265_),
    .X(_12266_));
 sky130_fd_sc_hd__or3_2 _16295_ (.A(_11050_),
    .B(\decode.regfile.registers_25[25] ),
    .C(_11089_),
    .X(_12267_));
 sky130_fd_sc_hd__o2111a_2 _16296_ (.A1(_10958_),
    .A2(\decode.regfile.registers_26[25] ),
    .B1(_11676_),
    .C1(_11338_),
    .D1(_11564_),
    .X(_12268_));
 sky130_fd_sc_hd__a31o_2 _16297_ (.A1(_11260_),
    .A2(_12266_),
    .A3(_12267_),
    .B1(_12268_),
    .X(_12269_));
 sky130_fd_sc_hd__or3_2 _16298_ (.A(_11679_),
    .B(\decode.regfile.registers_27[25] ),
    .C(_11869_),
    .X(_12270_));
 sky130_fd_sc_hd__o2111a_2 _16299_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[25] ),
    .B1(_11871_),
    .C1(_11681_),
    .D1(_11448_),
    .X(_12271_));
 sky130_fd_sc_hd__a31o_2 _16300_ (.A1(_11396_),
    .A2(_12269_),
    .A3(_12270_),
    .B1(_12271_),
    .X(_12272_));
 sky130_fd_sc_hd__o221a_2 _16301_ (.A1(_11646_),
    .A2(_11834_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[25] ),
    .C1(_12272_),
    .X(_12273_));
 sky130_fd_sc_hd__o221a_2 _16302_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[25] ),
    .B1(_12237_),
    .B2(_12273_),
    .C1(_12132_),
    .X(_00413_));
 sky130_fd_sc_hd__o2111a_2 _16303_ (.A1(_11942_),
    .A2(\decode.regfile.registers_30[26] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12274_));
 sky130_fd_sc_hd__and4_2 _16304_ (.A(\decode.regfile.registers_17[26] ),
    .B(_10988_),
    .C(_11113_),
    .D(_11118_),
    .X(_12275_));
 sky130_fd_sc_hd__a31o_2 _16305_ (.A1(\decode.regfile.registers_15[26] ),
    .A2(_11036_),
    .A3(_11205_),
    .B1(_11203_),
    .X(_12276_));
 sky130_fd_sc_hd__a21oi_2 _16306_ (.A1(\decode.regfile.registers_10[26] ),
    .A2(_11184_),
    .B1(_11181_),
    .Y(_12277_));
 sky130_fd_sc_hd__a221oi_2 _16307_ (.A1(\decode.regfile.registers_7[26] ),
    .A2(_11378_),
    .B1(_11170_),
    .B2(\decode.regfile.registers_6[26] ),
    .C1(_11281_),
    .Y(_12278_));
 sky130_fd_sc_hd__and4_2 _16308_ (.A(\decode.regfile.registers_1[26] ),
    .B(_11116_),
    .C(_11056_),
    .D(_11108_),
    .X(_12279_));
 sky130_fd_sc_hd__a211o_2 _16309_ (.A1(_11371_),
    .A2(\decode.regfile.registers_0[26] ),
    .B1(_11156_),
    .C1(_12279_),
    .X(_12280_));
 sky130_fd_sc_hd__o221ai_2 _16310_ (.A1(\decode.regfile.registers_2[26] ),
    .A2(_11369_),
    .B1(_11297_),
    .B2(_11121_),
    .C1(_12280_),
    .Y(_12281_));
 sky130_fd_sc_hd__o2bb2a_2 _16311_ (.A1_N(\decode.regfile.registers_3[26] ),
    .A2_N(_11614_),
    .B1(_11367_),
    .B2(_11178_),
    .X(_12282_));
 sky130_fd_sc_hd__nand2_2 _16312_ (.A(_12281_),
    .B(_12282_),
    .Y(_12283_));
 sky130_fd_sc_hd__a2111o_2 _16313_ (.A1(_11313_),
    .A2(\decode.regfile.registers_4[26] ),
    .B1(_10647_),
    .C1(_10629_),
    .D1(_11462_),
    .X(_12284_));
 sky130_fd_sc_hd__a32o_2 _16314_ (.A1(\decode.regfile.registers_5[26] ),
    .A2(_11192_),
    .A3(_11139_),
    .B1(_12283_),
    .B2(_12284_),
    .X(_12285_));
 sky130_fd_sc_hd__o21ai_2 _16315_ (.A1(_11318_),
    .A2(_11085_),
    .B1(_12285_),
    .Y(_12286_));
 sky130_fd_sc_hd__a2bb2oi_2 _16316_ (.A1_N(\decode.regfile.registers_9[26] ),
    .A2_N(_11365_),
    .B1(_12278_),
    .B2(_12286_),
    .Y(_12287_));
 sky130_fd_sc_hd__o211ai_2 _16317_ (.A1(\decode.regfile.registers_8[26] ),
    .A2(_11285_),
    .B1(_11382_),
    .C1(_12287_),
    .Y(_12288_));
 sky130_fd_sc_hd__a2bb2o_2 _16318_ (.A1_N(\decode.regfile.registers_11[26] ),
    .A2_N(_11364_),
    .B1(_12277_),
    .B2(_12288_),
    .X(_12289_));
 sky130_fd_sc_hd__nand2_2 _16319_ (.A(_11690_),
    .B(_12289_),
    .Y(_12290_));
 sky130_fd_sc_hd__o221a_2 _16320_ (.A1(_11194_),
    .A2(\decode.regfile.registers_12[26] ),
    .B1(\decode.regfile.registers_13[26] ),
    .B2(_11196_),
    .C1(_12074_),
    .X(_12291_));
 sky130_fd_sc_hd__a22o_2 _16321_ (.A1(\decode.regfile.registers_14[26] ),
    .A2(_12018_),
    .B1(_12290_),
    .B2(_12291_),
    .X(_12292_));
 sky130_fd_sc_hd__o31a_2 _16322_ (.A1(_11048_),
    .A2(_11054_),
    .A3(_11318_),
    .B1(_12292_),
    .X(_12293_));
 sky130_fd_sc_hd__o221a_2 _16323_ (.A1(\decode.regfile.registers_16[26] ),
    .A2(_11124_),
    .B1(_12276_),
    .B2(_12293_),
    .C1(_11127_),
    .X(_12294_));
 sky130_fd_sc_hd__o22a_2 _16324_ (.A1(_11059_),
    .A2(_11149_),
    .B1(_12275_),
    .B2(_12294_),
    .X(_12295_));
 sky130_fd_sc_hd__a211o_2 _16325_ (.A1(\decode.regfile.registers_18[26] ),
    .A2(_11455_),
    .B1(_11456_),
    .C1(_12295_),
    .X(_12296_));
 sky130_fd_sc_hd__o41a_2 _16326_ (.A1(\decode.regfile.registers_19[26] ),
    .A2(_11048_),
    .A3(_11215_),
    .A4(_11217_),
    .B1(_11219_),
    .X(_12297_));
 sky130_fd_sc_hd__a221o_2 _16327_ (.A1(\decode.regfile.registers_20[26] ),
    .A2(_11103_),
    .B1(_12296_),
    .B2(_12297_),
    .C1(_11222_),
    .X(_12298_));
 sky130_fd_sc_hd__o311a_2 _16328_ (.A1(\decode.regfile.registers_21[26] ),
    .A2(_11061_),
    .A3(_11099_),
    .B1(_11228_),
    .C1(_12298_),
    .X(_12299_));
 sky130_fd_sc_hd__a21oi_2 _16329_ (.A1(\decode.regfile.registers_22[26] ),
    .A2(_11096_),
    .B1(_12299_),
    .Y(_12300_));
 sky130_fd_sc_hd__a21oi_2 _16330_ (.A1(\decode.regfile.registers_23[26] ),
    .A2(_11232_),
    .B1(_11074_),
    .Y(_12301_));
 sky130_fd_sc_hd__o21ai_2 _16331_ (.A1(_11232_),
    .A2(_12300_),
    .B1(_12301_),
    .Y(_12302_));
 sky130_fd_sc_hd__o22a_2 _16332_ (.A1(\decode.regfile.registers_25[26] ),
    .A2(_11333_),
    .B1(_11336_),
    .B2(\decode.regfile.registers_24[26] ),
    .X(_12303_));
 sky130_fd_sc_hd__o2111a_2 _16333_ (.A1(_10958_),
    .A2(\decode.regfile.registers_26[26] ),
    .B1(_11676_),
    .C1(_11338_),
    .D1(_11564_),
    .X(_12304_));
 sky130_fd_sc_hd__a31o_2 _16334_ (.A1(_11260_),
    .A2(_12302_),
    .A3(_12303_),
    .B1(_12304_),
    .X(_12305_));
 sky130_fd_sc_hd__or3_2 _16335_ (.A(_11679_),
    .B(\decode.regfile.registers_27[26] ),
    .C(_11869_),
    .X(_12306_));
 sky130_fd_sc_hd__o2111a_2 _16336_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[26] ),
    .B1(_11871_),
    .C1(_11681_),
    .D1(_11448_),
    .X(_12307_));
 sky130_fd_sc_hd__a31o_2 _16337_ (.A1(_11396_),
    .A2(_12305_),
    .A3(_12306_),
    .B1(_12307_),
    .X(_12308_));
 sky130_fd_sc_hd__o221a_2 _16338_ (.A1(_11646_),
    .A2(_11834_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[26] ),
    .C1(_12308_),
    .X(_12309_));
 sky130_fd_sc_hd__o221a_2 _16339_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[26] ),
    .B1(_12274_),
    .B2(_12309_),
    .C1(_12132_),
    .X(_00414_));
 sky130_fd_sc_hd__o2111a_2 _16340_ (.A1(_11346_),
    .A2(\decode.regfile.registers_30[27] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12310_));
 sky130_fd_sc_hd__o2111a_2 _16341_ (.A1(_11435_),
    .A2(\decode.regfile.registers_24[27] ),
    .B1(_11244_),
    .C1(_11080_),
    .D1(_10991_),
    .X(_12311_));
 sky130_fd_sc_hd__o2111a_2 _16342_ (.A1(_11263_),
    .A2(\decode.regfile.registers_22[27] ),
    .B1(_11404_),
    .C1(_11264_),
    .D1(_11265_),
    .X(_12312_));
 sky130_fd_sc_hd__nand2_2 _16343_ (.A(\decode.regfile.registers_17[27] ),
    .B(_11356_),
    .Y(_12313_));
 sky130_fd_sc_hd__a31o_2 _16344_ (.A1(\decode.regfile.registers_3[27] ),
    .A2(_11110_),
    .A3(_11141_),
    .B1(_11145_),
    .X(_12314_));
 sky130_fd_sc_hd__inv_2 _16345_ (.A(\decode.regfile.registers_1[27] ),
    .Y(_12315_));
 sky130_fd_sc_hd__nand2_2 _16346_ (.A(_11371_),
    .B(\decode.regfile.registers_0[27] ),
    .Y(_12316_));
 sky130_fd_sc_hd__o221ai_2 _16347_ (.A1(_12315_),
    .A2(_11371_),
    .B1(_10646_),
    .B2(_11298_),
    .C1(_12316_),
    .Y(_12317_));
 sky130_fd_sc_hd__o311a_2 _16348_ (.A1(\decode.regfile.registers_2[27] ),
    .A2(_11190_),
    .A3(_11148_),
    .B1(_11151_),
    .C1(_12317_),
    .X(_12318_));
 sky130_fd_sc_hd__o32a_2 _16349_ (.A1(\decode.regfile.registers_4[27] ),
    .A2(_10636_),
    .A3(_11410_),
    .B1(_12314_),
    .B2(_12318_),
    .X(_12319_));
 sky130_fd_sc_hd__and3_2 _16350_ (.A(\decode.regfile.registers_5[27] ),
    .B(_11192_),
    .C(_11138_),
    .X(_12320_));
 sky130_fd_sc_hd__a21oi_2 _16351_ (.A1(_12319_),
    .A2(_12065_),
    .B1(_12320_),
    .Y(_12321_));
 sky130_fd_sc_hd__a221oi_2 _16352_ (.A1(\decode.regfile.registers_7[27] ),
    .A2(_11465_),
    .B1(_11466_),
    .B2(\decode.regfile.registers_6[27] ),
    .C1(_11166_),
    .Y(_12322_));
 sky130_fd_sc_hd__o21ai_2 _16353_ (.A1(_11289_),
    .A2(_12321_),
    .B1(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__a21o_2 _16354_ (.A1(\decode.regfile.registers_8[27] ),
    .A2(_11045_),
    .B1(_11174_),
    .X(_12324_));
 sky130_fd_sc_hd__a221o_2 _16355_ (.A1(\decode.regfile.registers_9[27] ),
    .A2(_11547_),
    .B1(_12323_),
    .B2(_12324_),
    .C1(_11509_),
    .X(_12325_));
 sky130_fd_sc_hd__o2bb2a_2 _16356_ (.A1_N(_11070_),
    .A2_N(_11470_),
    .B1(\decode.regfile.registers_10[27] ),
    .B2(_11382_),
    .X(_12326_));
 sky130_fd_sc_hd__a221o_2 _16357_ (.A1(\decode.regfile.registers_11[27] ),
    .A2(_11181_),
    .B1(_12325_),
    .B2(_12326_),
    .C1(_11187_),
    .X(_12327_));
 sky130_fd_sc_hd__o221a_2 _16358_ (.A1(_11194_),
    .A2(\decode.regfile.registers_12[27] ),
    .B1(\decode.regfile.registers_13[27] ),
    .B2(_11196_),
    .C1(_11198_),
    .X(_12328_));
 sky130_fd_sc_hd__nand2_2 _16359_ (.A(_12327_),
    .B(_12328_),
    .Y(_12329_));
 sky130_fd_sc_hd__a221oi_2 _16360_ (.A1(\decode.regfile.registers_14[27] ),
    .A2(_11360_),
    .B1(_11274_),
    .B2(\decode.regfile.registers_15[27] ),
    .C1(_11361_),
    .Y(_12330_));
 sky130_fd_sc_hd__nor2_2 _16361_ (.A(\decode.regfile.registers_16[27] ),
    .B(_11123_),
    .Y(_12331_));
 sky130_fd_sc_hd__a211o_2 _16362_ (.A1(_12329_),
    .A2(_12330_),
    .B1(_12331_),
    .C1(_11356_),
    .X(_12332_));
 sky130_fd_sc_hd__o2bb2a_2 _16363_ (.A1_N(_12313_),
    .A2_N(_12332_),
    .B1(_11059_),
    .B2(_11149_),
    .X(_12333_));
 sky130_fd_sc_hd__a211o_2 _16364_ (.A1(\decode.regfile.registers_18[27] ),
    .A2(_11269_),
    .B1(_11271_),
    .C1(_12333_),
    .X(_12334_));
 sky130_fd_sc_hd__o211a_2 _16365_ (.A1(\decode.regfile.registers_19[27] ),
    .A2(_11406_),
    .B1(_11325_),
    .C1(_12334_),
    .X(_12335_));
 sky130_fd_sc_hd__a211o_2 _16366_ (.A1(\decode.regfile.registers_20[27] ),
    .A2(_11102_),
    .B1(_11327_),
    .C1(_12335_),
    .X(_12336_));
 sky130_fd_sc_hd__o311a_2 _16367_ (.A1(\decode.regfile.registers_21[27] ),
    .A2(_11267_),
    .A3(_11098_),
    .B1(_11227_),
    .C1(_12336_),
    .X(_12337_));
 sky130_fd_sc_hd__o221a_2 _16368_ (.A1(\decode.regfile.registers_23[27] ),
    .A2(_11262_),
    .B1(_12312_),
    .B2(_12337_),
    .C1(_11335_),
    .X(_12338_));
 sky130_fd_sc_hd__o32a_2 _16369_ (.A1(_11076_),
    .A2(_11090_),
    .A3(\decode.regfile.registers_25[27] ),
    .B1(_12311_),
    .B2(_12338_),
    .X(_12339_));
 sky130_fd_sc_hd__o2111a_2 _16370_ (.A1(_10959_),
    .A2(\decode.regfile.registers_26[27] ),
    .B1(_11349_),
    .C1(_10980_),
    .D1(_11347_),
    .X(_12340_));
 sky130_fd_sc_hd__a21o_2 _16371_ (.A1(_12339_),
    .A2(_11486_),
    .B1(_12340_),
    .X(_12341_));
 sky130_fd_sc_hd__or3_2 _16372_ (.A(_11076_),
    .B(\decode.regfile.registers_27[27] ),
    .C(_11869_),
    .X(_12342_));
 sky130_fd_sc_hd__o2111a_2 _16373_ (.A1(_11756_),
    .A2(\decode.regfile.registers_28[27] ),
    .B1(_11871_),
    .C1(_11037_),
    .D1(_11448_),
    .X(_12343_));
 sky130_fd_sc_hd__a31o_2 _16374_ (.A1(_11396_),
    .A2(_12341_),
    .A3(_12342_),
    .B1(_12343_),
    .X(_12344_));
 sky130_fd_sc_hd__o221a_2 _16375_ (.A1(_10961_),
    .A2(_11834_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[27] ),
    .C1(_12344_),
    .X(_12345_));
 sky130_fd_sc_hd__o221a_2 _16376_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[27] ),
    .B1(_12310_),
    .B2(_12345_),
    .C1(_12132_),
    .X(_00415_));
 sky130_fd_sc_hd__o2111a_2 _16377_ (.A1(_11346_),
    .A2(\decode.regfile.registers_30[28] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12346_));
 sky130_fd_sc_hd__a31o_2 _16378_ (.A1(\decode.regfile.registers_15[28] ),
    .A2(_11036_),
    .A3(_11205_),
    .B1(_11202_),
    .X(_12347_));
 sky130_fd_sc_hd__a221o_2 _16379_ (.A1(\decode.regfile.registers_13[28] ),
    .A2(_11276_),
    .B1(_11407_),
    .B2(\decode.regfile.registers_12[28] ),
    .C1(_11360_),
    .X(_12348_));
 sky130_fd_sc_hd__a22o_2 _16380_ (.A1(_11071_),
    .A2(_11204_),
    .B1(_11184_),
    .B2(\decode.regfile.registers_10[28] ),
    .X(_12349_));
 sky130_fd_sc_hd__a31o_2 _16381_ (.A1(\decode.regfile.registers_5[28] ),
    .A2(_10636_),
    .A3(_11138_),
    .B1(_11169_),
    .X(_12350_));
 sky130_fd_sc_hd__a31o_2 _16382_ (.A1(\decode.regfile.registers_3[28] ),
    .A2(_11110_),
    .A3(_11141_),
    .B1(_11145_),
    .X(_12351_));
 sky130_fd_sc_hd__and4_2 _16383_ (.A(\decode.regfile.registers_1[28] ),
    .B(_11116_),
    .C(_11137_),
    .D(_11157_),
    .X(_12352_));
 sky130_fd_sc_hd__a21oi_2 _16384_ (.A1(\decode.regfile.registers_0[28] ),
    .A2(_11154_),
    .B1(_12352_),
    .Y(_12353_));
 sky130_fd_sc_hd__nor2_2 _16385_ (.A(\decode.regfile.registers_2[28] ),
    .B(_11296_),
    .Y(_12354_));
 sky130_fd_sc_hd__a211oi_2 _16386_ (.A1(_12353_),
    .A2(_11369_),
    .B1(_11614_),
    .C1(_12354_),
    .Y(_12355_));
 sky130_fd_sc_hd__a2111o_2 _16387_ (.A1(_11042_),
    .A2(\decode.regfile.registers_4[28] ),
    .B1(_11190_),
    .C1(_10628_),
    .D1(_11083_),
    .X(_12356_));
 sky130_fd_sc_hd__o21a_2 _16388_ (.A1(_12351_),
    .A2(_12355_),
    .B1(_12356_),
    .X(_12357_));
 sky130_fd_sc_hd__o32a_2 _16389_ (.A1(\decode.regfile.registers_6[28] ),
    .A2(_10637_),
    .A3(_11136_),
    .B1(_12350_),
    .B2(_12357_),
    .X(_12358_));
 sky130_fd_sc_hd__mux2_2 _16390_ (.A0(_12358_),
    .A1(\decode.regfile.registers_7[28] ),
    .S(_11378_),
    .X(_12359_));
 sky130_fd_sc_hd__o221a_2 _16391_ (.A1(\decode.regfile.registers_8[28] ),
    .A2(_11285_),
    .B1(_11365_),
    .B2(\decode.regfile.registers_9[28] ),
    .C1(_11381_),
    .X(_12360_));
 sky130_fd_sc_hd__o21a_2 _16392_ (.A1(_11134_),
    .A2(_12359_),
    .B1(_12360_),
    .X(_12361_));
 sky130_fd_sc_hd__o221a_2 _16393_ (.A1(_11364_),
    .A2(\decode.regfile.registers_11[28] ),
    .B1(_12349_),
    .B2(_12361_),
    .C1(_11690_),
    .X(_12362_));
 sky130_fd_sc_hd__a211o_2 _16394_ (.A1(\decode.regfile.registers_14[28] ),
    .A2(_11047_),
    .B1(_11053_),
    .C1(_11318_),
    .X(_12363_));
 sky130_fd_sc_hd__o21a_2 _16395_ (.A1(_12348_),
    .A2(_12362_),
    .B1(_12363_),
    .X(_12364_));
 sky130_fd_sc_hd__o22a_2 _16396_ (.A1(\decode.regfile.registers_16[28] ),
    .A2(_11359_),
    .B1(_12347_),
    .B2(_12364_),
    .X(_12365_));
 sky130_fd_sc_hd__a31o_2 _16397_ (.A1(_10988_),
    .A2(_11113_),
    .A3(_11119_),
    .B1(_12365_),
    .X(_12366_));
 sky130_fd_sc_hd__o32a_2 _16398_ (.A1(_11225_),
    .A2(_11125_),
    .A3(_11216_),
    .B1(\decode.regfile.registers_17[28] ),
    .B2(_11128_),
    .X(_12367_));
 sky130_fd_sc_hd__a221o_2 _16399_ (.A1(\decode.regfile.registers_18[28] ),
    .A2(_11269_),
    .B1(_12366_),
    .B2(_12367_),
    .C1(_11456_),
    .X(_12368_));
 sky130_fd_sc_hd__o211a_2 _16400_ (.A1(\decode.regfile.registers_19[28] ),
    .A2(_11453_),
    .B1(_11219_),
    .C1(_12368_),
    .X(_12369_));
 sky130_fd_sc_hd__a211o_2 _16401_ (.A1(\decode.regfile.registers_20[28] ),
    .A2(_11452_),
    .B1(_11223_),
    .C1(_12369_),
    .X(_12370_));
 sky130_fd_sc_hd__o32a_2 _16402_ (.A1(_11263_),
    .A2(_11217_),
    .A3(_11085_),
    .B1(\decode.regfile.registers_21[28] ),
    .B2(_11648_),
    .X(_12371_));
 sky130_fd_sc_hd__a22o_2 _16403_ (.A1(\decode.regfile.registers_22[28] ),
    .A2(_11096_),
    .B1(_12370_),
    .B2(_12371_),
    .X(_12372_));
 sky130_fd_sc_hd__a32o_2 _16404_ (.A1(_10991_),
    .A2(_11065_),
    .A3(_11080_),
    .B1(_11232_),
    .B2(\decode.regfile.registers_23[28] ),
    .X(_12373_));
 sky130_fd_sc_hd__a21o_2 _16405_ (.A1(_11088_),
    .A2(_12372_),
    .B1(_12373_),
    .X(_12374_));
 sky130_fd_sc_hd__o22a_2 _16406_ (.A1(\decode.regfile.registers_25[28] ),
    .A2(_11333_),
    .B1(_11336_),
    .B2(\decode.regfile.registers_24[28] ),
    .X(_12375_));
 sky130_fd_sc_hd__o2111a_2 _16407_ (.A1(_10958_),
    .A2(\decode.regfile.registers_26[28] ),
    .B1(_11676_),
    .C1(_11338_),
    .D1(_10992_),
    .X(_12376_));
 sky130_fd_sc_hd__a31o_2 _16408_ (.A1(_11260_),
    .A2(_12374_),
    .A3(_12375_),
    .B1(_12376_),
    .X(_12377_));
 sky130_fd_sc_hd__or3_2 _16409_ (.A(_11076_),
    .B(\decode.regfile.registers_27[28] ),
    .C(_11869_),
    .X(_12378_));
 sky130_fd_sc_hd__o2111a_2 _16410_ (.A1(_11446_),
    .A2(\decode.regfile.registers_28[28] ),
    .B1(_11871_),
    .C1(_11037_),
    .D1(_11448_),
    .X(_12379_));
 sky130_fd_sc_hd__a31o_2 _16411_ (.A1(_11396_),
    .A2(_12377_),
    .A3(_12378_),
    .B1(_12379_),
    .X(_12380_));
 sky130_fd_sc_hd__o221a_2 _16412_ (.A1(_10961_),
    .A2(_11834_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[28] ),
    .C1(_12380_),
    .X(_12381_));
 sky130_fd_sc_hd__o221a_2 _16413_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[28] ),
    .B1(_12346_),
    .B2(_12381_),
    .C1(_12132_),
    .X(_00416_));
 sky130_fd_sc_hd__o2111a_2 _16414_ (.A1(_11346_),
    .A2(\decode.regfile.registers_30[29] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12382_));
 sky130_fd_sc_hd__o2111a_2 _16415_ (.A1(_11446_),
    .A2(\decode.regfile.registers_26[29] ),
    .B1(_11447_),
    .C1(_11348_),
    .D1(_10993_),
    .X(_12383_));
 sky130_fd_sc_hd__o2111a_2 _16416_ (.A1(_11493_),
    .A2(\decode.regfile.registers_22[29] ),
    .B1(_11450_),
    .C1(_10978_),
    .D1(_10991_),
    .X(_12384_));
 sky130_fd_sc_hd__o221ai_2 _16417_ (.A1(\decode.regfile.registers_9[29] ),
    .A2(_11365_),
    .B1(\decode.regfile.registers_8[29] ),
    .B2(_11285_),
    .C1(_11382_),
    .Y(_12385_));
 sky130_fd_sc_hd__a31o_2 _16418_ (.A1(\decode.regfile.registers_3[29] ),
    .A2(_11110_),
    .A3(_11141_),
    .B1(_11146_),
    .X(_12386_));
 sky130_fd_sc_hd__inv_2 _16419_ (.A(\decode.regfile.registers_1[29] ),
    .Y(_12387_));
 sky130_fd_sc_hd__nand2_2 _16420_ (.A(_11371_),
    .B(\decode.regfile.registers_0[29] ),
    .Y(_12388_));
 sky130_fd_sc_hd__o221ai_2 _16421_ (.A1(_12387_),
    .A2(_11371_),
    .B1(_10646_),
    .B2(_11298_),
    .C1(_12388_),
    .Y(_12389_));
 sky130_fd_sc_hd__o311a_2 _16422_ (.A1(\decode.regfile.registers_2[29] ),
    .A2(_11503_),
    .A3(_11148_),
    .B1(_11152_),
    .C1(_12389_),
    .X(_12390_));
 sky130_fd_sc_hd__a2111o_2 _16423_ (.A1(_11043_),
    .A2(\decode.regfile.registers_4[29] ),
    .B1(_11503_),
    .C1(_10629_),
    .D1(_11083_),
    .X(_12391_));
 sky130_fd_sc_hd__o21a_2 _16424_ (.A1(_12386_),
    .A2(_12390_),
    .B1(_12391_),
    .X(_12392_));
 sky130_fd_sc_hd__a311o_2 _16425_ (.A1(\decode.regfile.registers_5[29] ),
    .A2(_11280_),
    .A3(_11139_),
    .B1(_11466_),
    .C1(_12392_),
    .X(_12393_));
 sky130_fd_sc_hd__a211o_2 _16426_ (.A1(_11044_),
    .A2(\decode.regfile.registers_6[29] ),
    .B1(_11085_),
    .C1(_11318_),
    .X(_12394_));
 sky130_fd_sc_hd__a221oi_2 _16427_ (.A1(\decode.regfile.registers_7[29] ),
    .A2(_11378_),
    .B1(_12393_),
    .B2(_12394_),
    .C1(_11134_),
    .Y(_12395_));
 sky130_fd_sc_hd__a2bb2o_2 _16428_ (.A1_N(_12385_),
    .A2_N(_12395_),
    .B1(_11184_),
    .B2(\decode.regfile.registers_10[29] ),
    .X(_12396_));
 sky130_fd_sc_hd__a31o_2 _16429_ (.A1(\decode.regfile.registers_11[29] ),
    .A2(_11071_),
    .A3(_11204_),
    .B1(_11407_),
    .X(_12397_));
 sky130_fd_sc_hd__a21o_2 _16430_ (.A1(_11364_),
    .A2(_12396_),
    .B1(_12397_),
    .X(_12398_));
 sky130_fd_sc_hd__a2111o_2 _16431_ (.A1(_11047_),
    .A2(\decode.regfile.registers_12[29] ),
    .B1(_10650_),
    .C1(_11053_),
    .D1(_10632_),
    .X(_12399_));
 sky130_fd_sc_hd__a32o_2 _16432_ (.A1(\decode.regfile.registers_13[29] ),
    .A2(_10640_),
    .A3(_11187_),
    .B1(_12398_),
    .B2(_12399_),
    .X(_12400_));
 sky130_fd_sc_hd__a32o_2 _16433_ (.A1(\decode.regfile.registers_15[29] ),
    .A2(_11036_),
    .A3(_11205_),
    .B1(_11208_),
    .B2(\decode.regfile.registers_14[29] ),
    .X(_12401_));
 sky130_fd_sc_hd__a211o_2 _16434_ (.A1(_11199_),
    .A2(_12400_),
    .B1(_12401_),
    .C1(_11203_),
    .X(_12402_));
 sky130_fd_sc_hd__o211a_2 _16435_ (.A1(_11124_),
    .A2(\decode.regfile.registers_16[29] ),
    .B1(_11128_),
    .C1(_12402_),
    .X(_12403_));
 sky130_fd_sc_hd__a41o_2 _16436_ (.A1(\decode.regfile.registers_17[29] ),
    .A2(_10989_),
    .A3(_11114_),
    .A4(_11119_),
    .B1(_12403_),
    .X(_12404_));
 sky130_fd_sc_hd__o2111a_2 _16437_ (.A1(\decode.regfile.registers_18[29] ),
    .A2(_10956_),
    .B1(_11114_),
    .C1(_10989_),
    .D1(_10977_),
    .X(_12405_));
 sky130_fd_sc_hd__a21o_2 _16438_ (.A1(_11106_),
    .A2(_12404_),
    .B1(_12405_),
    .X(_12406_));
 sky130_fd_sc_hd__o41a_2 _16439_ (.A1(\decode.regfile.registers_19[29] ),
    .A2(_11049_),
    .A3(_11215_),
    .A4(_11217_),
    .B1(_11454_),
    .X(_12407_));
 sky130_fd_sc_hd__a221o_2 _16440_ (.A1(\decode.regfile.registers_20[29] ),
    .A2(_11452_),
    .B1(_12406_),
    .B2(_12407_),
    .C1(_11223_),
    .X(_12408_));
 sky130_fd_sc_hd__o311a_2 _16441_ (.A1(\decode.regfile.registers_21[29] ),
    .A2(_11061_),
    .A3(_11100_),
    .B1(_11229_),
    .C1(_12408_),
    .X(_12409_));
 sky130_fd_sc_hd__o22a_2 _16442_ (.A1(\decode.regfile.registers_23[29] ),
    .A2(_11088_),
    .B1(_12384_),
    .B2(_12409_),
    .X(_12410_));
 sky130_fd_sc_hd__o22a_2 _16443_ (.A1(\decode.regfile.registers_25[29] ),
    .A2(_11483_),
    .B1(_11484_),
    .B2(\decode.regfile.registers_24[29] ),
    .X(_12411_));
 sky130_fd_sc_hd__o211a_2 _16444_ (.A1(_11075_),
    .A2(_12410_),
    .B1(_12411_),
    .C1(_11486_),
    .X(_12412_));
 sky130_fd_sc_hd__o32a_2 _16445_ (.A1(_11251_),
    .A2(_11259_),
    .A3(\decode.regfile.registers_27[29] ),
    .B1(_12383_),
    .B2(_12412_),
    .X(_12413_));
 sky130_fd_sc_hd__o221a_2 _16446_ (.A1(_11489_),
    .A2(\decode.regfile.registers_28[29] ),
    .B1(\decode.regfile.registers_29[29] ),
    .B2(_11063_),
    .C1(_11245_),
    .X(_12414_));
 sky130_fd_sc_hd__o21a_2 _16447_ (.A1(_11445_),
    .A2(_12413_),
    .B1(_12414_),
    .X(_12415_));
 sky130_fd_sc_hd__o221a_2 _16448_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[29] ),
    .B1(_12382_),
    .B2(_12415_),
    .C1(_12132_),
    .X(_00417_));
 sky130_fd_sc_hd__o2111a_2 _16449_ (.A1(_11346_),
    .A2(\decode.regfile.registers_30[30] ),
    .B1(_12095_),
    .C1(_12096_),
    .D1(_12097_),
    .X(_12416_));
 sky130_fd_sc_hd__o2111a_2 _16450_ (.A1(_11263_),
    .A2(\decode.regfile.registers_22[30] ),
    .B1(_11404_),
    .C1(_11264_),
    .D1(_11265_),
    .X(_12417_));
 sky130_fd_sc_hd__a221o_2 _16451_ (.A1(\decode.regfile.registers_14[30] ),
    .A2(_11207_),
    .B1(_11273_),
    .B2(\decode.regfile.registers_15[30] ),
    .C1(_11361_),
    .X(_12418_));
 sky130_fd_sc_hd__a31o_2 _16452_ (.A1(\decode.regfile.registers_11[30] ),
    .A2(_11069_),
    .A3(_11167_),
    .B1(_11277_),
    .X(_12419_));
 sky130_fd_sc_hd__a221o_2 _16453_ (.A1(\decode.regfile.registers_7[30] ),
    .A2(_11308_),
    .B1(_11169_),
    .B2(\decode.regfile.registers_6[30] ),
    .C1(_11133_),
    .X(_12420_));
 sky130_fd_sc_hd__or3b_2 _16454_ (.A(_10647_),
    .B(_11097_),
    .C_N(\decode.regfile.registers_5[30] ),
    .X(_12421_));
 sky130_fd_sc_hd__a31o_2 _16455_ (.A1(\decode.regfile.registers_3[30] ),
    .A2(_11110_),
    .A3(_11141_),
    .B1(_11145_),
    .X(_12422_));
 sky130_fd_sc_hd__and4_2 _16456_ (.A(\decode.regfile.registers_1[30] ),
    .B(_11115_),
    .C(_11056_),
    .D(_11108_),
    .X(_12423_));
 sky130_fd_sc_hd__a211o_2 _16457_ (.A1(_11300_),
    .A2(\decode.regfile.registers_0[30] ),
    .B1(_11155_),
    .C1(_12423_),
    .X(_12424_));
 sky130_fd_sc_hd__o311a_2 _16458_ (.A1(\decode.regfile.registers_2[30] ),
    .A2(_11190_),
    .A3(_11148_),
    .B1(_11151_),
    .C1(_12424_),
    .X(_12425_));
 sky130_fd_sc_hd__a2111o_2 _16459_ (.A1(_11043_),
    .A2(\decode.regfile.registers_4[30] ),
    .B1(_11503_),
    .C1(_10629_),
    .D1(_11083_),
    .X(_12426_));
 sky130_fd_sc_hd__o21ai_2 _16460_ (.A1(_12422_),
    .A2(_12425_),
    .B1(_12426_),
    .Y(_12427_));
 sky130_fd_sc_hd__a21oi_2 _16461_ (.A1(_12421_),
    .A2(_12427_),
    .B1(_11289_),
    .Y(_12428_));
 sky130_fd_sc_hd__o221a_2 _16462_ (.A1(\decode.regfile.registers_8[30] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(\decode.regfile.registers_9[30] ),
    .C1(_11131_),
    .X(_12429_));
 sky130_fd_sc_hd__o21a_2 _16463_ (.A1(_12420_),
    .A2(_12428_),
    .B1(_12429_),
    .X(_12430_));
 sky130_fd_sc_hd__a211o_2 _16464_ (.A1(\decode.regfile.registers_10[30] ),
    .A2(_11509_),
    .B1(_12419_),
    .C1(_12430_),
    .X(_12431_));
 sky130_fd_sc_hd__a2111o_2 _16465_ (.A1(_11045_),
    .A2(\decode.regfile.registers_12[30] ),
    .B1(_10649_),
    .C1(_11051_),
    .D1(_10631_),
    .X(_12432_));
 sky130_fd_sc_hd__a32o_2 _16466_ (.A1(\decode.regfile.registers_13[30] ),
    .A2(_10639_),
    .A3(_11186_),
    .B1(_12431_),
    .B2(_12432_),
    .X(_12433_));
 sky130_fd_sc_hd__o31a_2 _16467_ (.A1(_10650_),
    .A2(_10625_),
    .A3(_11053_),
    .B1(_12433_),
    .X(_12434_));
 sky130_fd_sc_hd__o22a_2 _16468_ (.A1(\decode.regfile.registers_16[30] ),
    .A2(_11123_),
    .B1(_12418_),
    .B2(_12434_),
    .X(_12435_));
 sky130_fd_sc_hd__a31o_2 _16469_ (.A1(_10652_),
    .A2(_11112_),
    .A3(_11118_),
    .B1(_12435_),
    .X(_12436_));
 sky130_fd_sc_hd__o32a_2 _16470_ (.A1(_10642_),
    .A2(_11125_),
    .A3(_11104_),
    .B1(\decode.regfile.registers_17[30] ),
    .B2(_11127_),
    .X(_12437_));
 sky130_fd_sc_hd__a221o_2 _16471_ (.A1(\decode.regfile.registers_18[30] ),
    .A2(_11269_),
    .B1(_12436_),
    .B2(_12437_),
    .C1(_11271_),
    .X(_12438_));
 sky130_fd_sc_hd__o211a_2 _16472_ (.A1(\decode.regfile.registers_19[30] ),
    .A2(_11406_),
    .B1(_11325_),
    .C1(_12438_),
    .X(_12439_));
 sky130_fd_sc_hd__a211o_2 _16473_ (.A1(\decode.regfile.registers_20[30] ),
    .A2(_11103_),
    .B1(_11327_),
    .C1(_12439_),
    .X(_12440_));
 sky130_fd_sc_hd__o311a_2 _16474_ (.A1(\decode.regfile.registers_21[30] ),
    .A2(_11267_),
    .A3(_11099_),
    .B1(_11228_),
    .C1(_12440_),
    .X(_12441_));
 sky130_fd_sc_hd__o22a_2 _16475_ (.A1(\decode.regfile.registers_23[30] ),
    .A2(_11087_),
    .B1(_12417_),
    .B2(_12441_),
    .X(_12442_));
 sky130_fd_sc_hd__a31o_2 _16476_ (.A1(_10992_),
    .A2(_11244_),
    .A3(_11261_),
    .B1(_12442_),
    .X(_12443_));
 sky130_fd_sc_hd__o22a_2 _16477_ (.A1(\decode.regfile.registers_25[30] ),
    .A2(_11333_),
    .B1(_11336_),
    .B2(\decode.regfile.registers_24[30] ),
    .X(_12444_));
 sky130_fd_sc_hd__o2111a_2 _16478_ (.A1(_10958_),
    .A2(\decode.regfile.registers_26[30] ),
    .B1(_11676_),
    .C1(_11338_),
    .D1(_10992_),
    .X(_12445_));
 sky130_fd_sc_hd__a31o_2 _16479_ (.A1(_11260_),
    .A2(_12443_),
    .A3(_12444_),
    .B1(_12445_),
    .X(_12446_));
 sky130_fd_sc_hd__or3_2 _16480_ (.A(_11076_),
    .B(\decode.regfile.registers_27[30] ),
    .C(_11869_),
    .X(_12447_));
 sky130_fd_sc_hd__o2111a_2 _16481_ (.A1(_11446_),
    .A2(\decode.regfile.registers_28[30] ),
    .B1(_11871_),
    .C1(_11037_),
    .D1(_11448_),
    .X(_12448_));
 sky130_fd_sc_hd__a31o_2 _16482_ (.A1(_11396_),
    .A2(_12446_),
    .A3(_12447_),
    .B1(_12448_),
    .X(_12449_));
 sky130_fd_sc_hd__o221a_2 _16483_ (.A1(_10961_),
    .A2(_11834_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[30] ),
    .C1(_12449_),
    .X(_12450_));
 sky130_fd_sc_hd__o221a_2 _16484_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[30] ),
    .B1(_12416_),
    .B2(_12450_),
    .C1(_12132_),
    .X(_00418_));
 sky130_fd_sc_hd__o2111a_2 _16485_ (.A1(_11346_),
    .A2(\decode.regfile.registers_30[31] ),
    .B1(_11038_),
    .C1(_10981_),
    .D1(_10994_),
    .X(_12451_));
 sky130_fd_sc_hd__o2111a_2 _16486_ (.A1(_11435_),
    .A2(\decode.regfile.registers_24[31] ),
    .B1(_11065_),
    .C1(_11080_),
    .D1(_10991_),
    .X(_12452_));
 sky130_fd_sc_hd__o2111a_2 _16487_ (.A1(_11263_),
    .A2(\decode.regfile.registers_22[31] ),
    .B1(_11404_),
    .C1(_11264_),
    .D1(_11265_),
    .X(_12453_));
 sky130_fd_sc_hd__a221o_2 _16488_ (.A1(\decode.regfile.registers_14[31] ),
    .A2(_11207_),
    .B1(_11273_),
    .B2(\decode.regfile.registers_15[31] ),
    .C1(_11361_),
    .X(_12454_));
 sky130_fd_sc_hd__a22o_2 _16489_ (.A1(\decode.regfile.registers_13[31] ),
    .A2(_11276_),
    .B1(_11407_),
    .B2(\decode.regfile.registers_12[31] ),
    .X(_12455_));
 sky130_fd_sc_hd__nand2_2 _16490_ (.A(\decode.regfile.registers_1[31] ),
    .B(_11539_),
    .Y(_12456_));
 sky130_fd_sc_hd__nand2_2 _16491_ (.A(_11300_),
    .B(\decode.regfile.registers_0[31] ),
    .Y(_12457_));
 sky130_fd_sc_hd__o211ai_2 _16492_ (.A1(_10646_),
    .A2(_11298_),
    .B1(_12456_),
    .C1(_12457_),
    .Y(_12458_));
 sky130_fd_sc_hd__o221ai_2 _16493_ (.A1(\decode.regfile.registers_2[31] ),
    .A2(_11296_),
    .B1(_11297_),
    .B2(_11121_),
    .C1(_12458_),
    .Y(_12459_));
 sky130_fd_sc_hd__o2bb2a_2 _16494_ (.A1_N(\decode.regfile.registers_3[31] ),
    .A2_N(_11292_),
    .B1(_11293_),
    .B2(_10635_),
    .X(_12460_));
 sky130_fd_sc_hd__nand2_2 _16495_ (.A(_12459_),
    .B(_12460_),
    .Y(_12461_));
 sky130_fd_sc_hd__a2111o_2 _16496_ (.A1(_11042_),
    .A2(\decode.regfile.registers_4[31] ),
    .B1(_11190_),
    .C1(_10628_),
    .D1(_11083_),
    .X(_12462_));
 sky130_fd_sc_hd__a22oi_2 _16497_ (.A1(\decode.regfile.registers_5[31] ),
    .A2(_11291_),
    .B1(_12461_),
    .B2(_12462_),
    .Y(_12463_));
 sky130_fd_sc_hd__a221oi_2 _16498_ (.A1(\decode.regfile.registers_7[31] ),
    .A2(_11308_),
    .B1(_11169_),
    .B2(\decode.regfile.registers_6[31] ),
    .C1(_11133_),
    .Y(_12464_));
 sky130_fd_sc_hd__o21ai_2 _16499_ (.A1(_11289_),
    .A2(_12463_),
    .B1(_12464_),
    .Y(_12465_));
 sky130_fd_sc_hd__o22a_2 _16500_ (.A1(\decode.regfile.registers_8[31] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(\decode.regfile.registers_9[31] ),
    .X(_12466_));
 sky130_fd_sc_hd__and3_2 _16501_ (.A(_11381_),
    .B(_12465_),
    .C(_12466_),
    .X(_12467_));
 sky130_fd_sc_hd__a221o_2 _16502_ (.A1(_11070_),
    .A2(_11470_),
    .B1(_11509_),
    .B2(\decode.regfile.registers_10[31] ),
    .C1(_12467_),
    .X(_12468_));
 sky130_fd_sc_hd__o211a_2 _16503_ (.A1(_11364_),
    .A2(\decode.regfile.registers_11[31] ),
    .B1(_11690_),
    .C1(_12468_),
    .X(_12469_));
 sky130_fd_sc_hd__o32a_2 _16504_ (.A1(_10650_),
    .A2(_10625_),
    .A3(_11053_),
    .B1(_12455_),
    .B2(_12469_),
    .X(_12470_));
 sky130_fd_sc_hd__o22a_2 _16505_ (.A1(\decode.regfile.registers_16[31] ),
    .A2(_11359_),
    .B1(_12454_),
    .B2(_12470_),
    .X(_12471_));
 sky130_fd_sc_hd__o32a_2 _16506_ (.A1(_10640_),
    .A2(_11125_),
    .A3(_11104_),
    .B1(\decode.regfile.registers_17[31] ),
    .B2(_11126_),
    .X(_12472_));
 sky130_fd_sc_hd__o21a_2 _16507_ (.A1(_11357_),
    .A2(_12471_),
    .B1(_12472_),
    .X(_12473_));
 sky130_fd_sc_hd__a211o_2 _16508_ (.A1(\decode.regfile.registers_18[31] ),
    .A2(_11269_),
    .B1(_11271_),
    .C1(_12473_),
    .X(_12474_));
 sky130_fd_sc_hd__o211a_2 _16509_ (.A1(\decode.regfile.registers_19[31] ),
    .A2(_11406_),
    .B1(_11325_),
    .C1(_12474_),
    .X(_12475_));
 sky130_fd_sc_hd__a211o_2 _16510_ (.A1(\decode.regfile.registers_20[31] ),
    .A2(_11102_),
    .B1(_11327_),
    .C1(_12475_),
    .X(_12476_));
 sky130_fd_sc_hd__o311a_2 _16511_ (.A1(\decode.regfile.registers_21[31] ),
    .A2(_11267_),
    .A3(_11098_),
    .B1(_11227_),
    .C1(_12476_),
    .X(_12477_));
 sky130_fd_sc_hd__o221a_2 _16512_ (.A1(\decode.regfile.registers_23[31] ),
    .A2(_11262_),
    .B1(_12453_),
    .B2(_12477_),
    .C1(_11335_),
    .X(_12478_));
 sky130_fd_sc_hd__o32a_2 _16513_ (.A1(_11050_),
    .A2(_11090_),
    .A3(\decode.regfile.registers_25[31] ),
    .B1(_12452_),
    .B2(_12478_),
    .X(_12479_));
 sky130_fd_sc_hd__o2111a_2 _16514_ (.A1(_11436_),
    .A2(\decode.regfile.registers_26[31] ),
    .B1(_11349_),
    .C1(_10980_),
    .D1(_11347_),
    .X(_12480_));
 sky130_fd_sc_hd__a21o_2 _16515_ (.A1(_12479_),
    .A2(_11236_),
    .B1(_12480_),
    .X(_12481_));
 sky130_fd_sc_hd__or3_2 _16516_ (.A(_11076_),
    .B(\decode.regfile.registers_27[31] ),
    .C(_11257_),
    .X(_12482_));
 sky130_fd_sc_hd__o2111a_2 _16517_ (.A1(_11446_),
    .A2(\decode.regfile.registers_28[31] ),
    .B1(_11066_),
    .C1(_11037_),
    .D1(_11448_),
    .X(_12483_));
 sky130_fd_sc_hd__a31o_2 _16518_ (.A1(_11396_),
    .A2(_12481_),
    .A3(_12482_),
    .B1(_12483_),
    .X(_12484_));
 sky130_fd_sc_hd__o221a_2 _16519_ (.A1(_10961_),
    .A2(_11252_),
    .B1(_11944_),
    .B2(\decode.regfile.registers_29[31] ),
    .C1(_12484_),
    .X(_12485_));
 sky130_fd_sc_hd__o221a_2 _16520_ (.A1(_12133_),
    .A2(\decode.regfile.registers_31[31] ),
    .B1(_12451_),
    .B2(_12485_),
    .C1(_11248_),
    .X(_00419_));
 sky130_fd_sc_hd__and4_2 _16521_ (.A(_11027_),
    .B(_11015_),
    .C(_11012_),
    .D(_11011_),
    .X(_12486_));
 sky130_fd_sc_hd__buf_1 _16522_ (.A(_12486_),
    .X(_12487_));
 sky130_fd_sc_hd__nand2_2 _16523_ (.A(_10598_),
    .B(\decode.immGen._imm_T_24[17] ),
    .Y(_12488_));
 sky130_fd_sc_hd__buf_1 _16524_ (.A(_12488_),
    .X(_12489_));
 sky130_fd_sc_hd__buf_1 _16525_ (.A(_12489_),
    .X(_12490_));
 sky130_fd_sc_hd__buf_1 _16526_ (.A(_12490_),
    .X(_12491_));
 sky130_fd_sc_hd__or4b_2 _16527_ (.A(_10939_),
    .B(_12491_),
    .C(_11011_),
    .D_N(_10928_),
    .X(_12492_));
 sky130_fd_sc_hd__buf_1 _16528_ (.A(_12492_),
    .X(_12493_));
 sky130_fd_sc_hd__buf_1 _16529_ (.A(_10926_),
    .X(_12494_));
 sky130_fd_sc_hd__or4_2 _16530_ (.A(_11010_),
    .B(_12494_),
    .C(_12491_),
    .D(_10939_),
    .X(_12495_));
 sky130_fd_sc_hd__buf_1 _16531_ (.A(_12495_),
    .X(_12496_));
 sky130_fd_sc_hd__buf_1 _16532_ (.A(_11016_),
    .X(_12497_));
 sky130_fd_sc_hd__buf_1 _16533_ (.A(_12497_),
    .X(_12498_));
 sky130_fd_sc_hd__buf_1 _16534_ (.A(_12498_),
    .X(_12499_));
 sky130_fd_sc_hd__nand2_2 _16535_ (.A(_12499_),
    .B(_10611_),
    .Y(_12500_));
 sky130_fd_sc_hd__nand2_2 _16536_ (.A(_10934_),
    .B(_10597_),
    .Y(_12501_));
 sky130_fd_sc_hd__buf_1 _16537_ (.A(_12501_),
    .X(_12502_));
 sky130_fd_sc_hd__buf_1 _16538_ (.A(_12502_),
    .X(_12503_));
 sky130_fd_sc_hd__buf_2 _16539_ (.A(_12503_),
    .X(_12504_));
 sky130_fd_sc_hd__buf_1 _16540_ (.A(_12504_),
    .X(_12505_));
 sky130_fd_sc_hd__buf_1 _16541_ (.A(_12505_),
    .X(_12506_));
 sky130_fd_sc_hd__buf_1 _16542_ (.A(_12506_),
    .X(_12507_));
 sky130_fd_sc_hd__buf_1 _16543_ (.A(_10614_),
    .X(_12508_));
 sky130_fd_sc_hd__nand2_2 _16544_ (.A(_10601_),
    .B(_12508_),
    .Y(_12509_));
 sky130_fd_sc_hd__buf_1 _16545_ (.A(_12509_),
    .X(_12510_));
 sky130_fd_sc_hd__buf_1 _16546_ (.A(_12510_),
    .X(_12511_));
 sky130_fd_sc_hd__buf_1 _16547_ (.A(_12511_),
    .X(_12512_));
 sky130_fd_sc_hd__or4_2 _16548_ (.A(_10595_),
    .B(_10606_),
    .C(_11012_),
    .D(_12512_),
    .X(_12513_));
 sky130_fd_sc_hd__or4_2 _16549_ (.A(_10595_),
    .B(_11009_),
    .C(_10925_),
    .D(_12504_),
    .X(_12514_));
 sky130_fd_sc_hd__buf_1 _16550_ (.A(_12514_),
    .X(_12515_));
 sky130_fd_sc_hd__buf_1 _16551_ (.A(_12515_),
    .X(_12516_));
 sky130_fd_sc_hd__o22ai_2 _16552_ (.A1(\decode.regfile.registers_25[0] ),
    .A2(_12513_),
    .B1(_12516_),
    .B2(\decode.regfile.registers_24[0] ),
    .Y(_12517_));
 sky130_fd_sc_hd__or3b_2 _16553_ (.A(_10594_),
    .B(_10604_),
    .C_N(_10924_),
    .X(_12518_));
 sky130_fd_sc_hd__buf_1 _16554_ (.A(_12518_),
    .X(_12519_));
 sky130_fd_sc_hd__buf_1 _16555_ (.A(_12519_),
    .X(_12520_));
 sky130_fd_sc_hd__or4_2 _16556_ (.A(_11015_),
    .B(_10937_),
    .C(\decode.regfile.registers_23[0] ),
    .D(_12520_),
    .X(_12521_));
 sky130_fd_sc_hd__nor2b_2 _16557_ (.A(_10597_),
    .B_N(\decode.immGen._imm_T_24[17] ),
    .Y(_12522_));
 sky130_fd_sc_hd__buf_1 _16558_ (.A(_12522_),
    .X(_12523_));
 sky130_fd_sc_hd__buf_1 _16559_ (.A(_11021_),
    .X(_12524_));
 sky130_fd_sc_hd__buf_1 _16560_ (.A(_12524_),
    .X(_12525_));
 sky130_fd_sc_hd__and4b_2 _16561_ (.A_N(_10925_),
    .B(_12523_),
    .C(_12525_),
    .D(_11009_),
    .X(_12526_));
 sky130_fd_sc_hd__buf_1 _16562_ (.A(_12526_),
    .X(_12527_));
 sky130_fd_sc_hd__buf_1 _16563_ (.A(_12527_),
    .X(_12528_));
 sky130_fd_sc_hd__and2b_2 _16564_ (.A_N(\decode.immGen._imm_T_24[16] ),
    .B(\decode.immGen._imm_T_24[15] ),
    .X(_12529_));
 sky130_fd_sc_hd__buf_1 _16565_ (.A(_12529_),
    .X(_12530_));
 sky130_fd_sc_hd__buf_1 _16566_ (.A(_12530_),
    .X(_12531_));
 sky130_fd_sc_hd__buf_1 _16567_ (.A(_12531_),
    .X(_12532_));
 sky130_fd_sc_hd__buf_1 _16568_ (.A(_12532_),
    .X(_12533_));
 sky130_fd_sc_hd__buf_1 _16569_ (.A(_12533_),
    .X(_12534_));
 sky130_fd_sc_hd__buf_1 _16570_ (.A(_12534_),
    .X(_12535_));
 sky130_fd_sc_hd__and3_2 _16571_ (.A(_12524_),
    .B(_12523_),
    .C(_12535_),
    .X(_12536_));
 sky130_fd_sc_hd__buf_1 _16572_ (.A(_12536_),
    .X(_12537_));
 sky130_fd_sc_hd__buf_1 _16573_ (.A(_12537_),
    .X(_12538_));
 sky130_fd_sc_hd__or2_2 _16574_ (.A(_10608_),
    .B(_12508_),
    .X(_12539_));
 sky130_fd_sc_hd__buf_1 _16575_ (.A(_12539_),
    .X(_12540_));
 sky130_fd_sc_hd__buf_1 _16576_ (.A(_12540_),
    .X(_12541_));
 sky130_fd_sc_hd__buf_1 _16577_ (.A(_12541_),
    .X(_12542_));
 sky130_fd_sc_hd__or4_2 _16578_ (.A(_10594_),
    .B(_10598_),
    .C(_10935_),
    .D(_12542_),
    .X(_12543_));
 sky130_fd_sc_hd__buf_1 _16579_ (.A(_12543_),
    .X(_12544_));
 sky130_fd_sc_hd__buf_1 _16580_ (.A(_12544_),
    .X(_12545_));
 sky130_fd_sc_hd__buf_1 _16581_ (.A(_11024_),
    .X(_12546_));
 sky130_fd_sc_hd__nor2_2 _16582_ (.A(_10607_),
    .B(_10614_),
    .Y(_12547_));
 sky130_fd_sc_hd__buf_1 _16583_ (.A(_12547_),
    .X(_12548_));
 sky130_fd_sc_hd__buf_1 _16584_ (.A(_12548_),
    .X(_12549_));
 sky130_fd_sc_hd__buf_1 _16585_ (.A(_12549_),
    .X(_12550_));
 sky130_fd_sc_hd__buf_1 _16586_ (.A(_12550_),
    .X(_12551_));
 sky130_fd_sc_hd__buf_1 _16587_ (.A(_12551_),
    .X(_12552_));
 sky130_fd_sc_hd__buf_1 _16588_ (.A(_12552_),
    .X(_12553_));
 sky130_fd_sc_hd__buf_1 _16589_ (.A(_12523_),
    .X(_12554_));
 sky130_fd_sc_hd__buf_1 _16590_ (.A(_10611_),
    .X(_12555_));
 sky130_fd_sc_hd__nor2_2 _16591_ (.A(_10597_),
    .B(\decode.immGen._imm_T_24[17] ),
    .Y(_12556_));
 sky130_fd_sc_hd__buf_1 _16592_ (.A(_12556_),
    .X(_12557_));
 sky130_fd_sc_hd__buf_1 _16593_ (.A(_12557_),
    .X(_12558_));
 sky130_fd_sc_hd__buf_1 _16594_ (.A(_12558_),
    .X(_12559_));
 sky130_fd_sc_hd__and4_2 _16595_ (.A(_11020_),
    .B(_12555_),
    .C(_10923_),
    .D(_12559_),
    .X(_12560_));
 sky130_fd_sc_hd__buf_1 _16596_ (.A(_12560_),
    .X(_12561_));
 sky130_fd_sc_hd__buf_1 _16597_ (.A(_12561_),
    .X(_12562_));
 sky130_fd_sc_hd__a32o_2 _16598_ (.A1(_12546_),
    .A2(_12553_),
    .A3(_12554_),
    .B1(_12562_),
    .B2(\decode.regfile.registers_19[0] ),
    .X(_12563_));
 sky130_fd_sc_hd__or4_2 _16599_ (.A(_10598_),
    .B(_10588_),
    .C(_10618_),
    .D(_12500_),
    .X(_12564_));
 sky130_fd_sc_hd__buf_1 _16600_ (.A(_12564_),
    .X(_12565_));
 sky130_fd_sc_hd__buf_1 _16601_ (.A(_12565_),
    .X(_12566_));
 sky130_fd_sc_hd__buf_1 _16602_ (.A(_12559_),
    .X(_12567_));
 sky130_fd_sc_hd__buf_1 _16603_ (.A(_12567_),
    .X(_12568_));
 sky130_fd_sc_hd__buf_1 _16604_ (.A(_12568_),
    .X(_12569_));
 sky130_fd_sc_hd__and4b_2 _16605_ (.A_N(_10923_),
    .B(_12559_),
    .C(_11020_),
    .D(_12555_),
    .X(_12570_));
 sky130_fd_sc_hd__buf_1 _16606_ (.A(_12570_),
    .X(_12571_));
 sky130_fd_sc_hd__buf_1 _16607_ (.A(_12571_),
    .X(_12572_));
 sky130_fd_sc_hd__a41o_2 _16608_ (.A1(\decode.regfile.registers_17[0] ),
    .A2(_12525_),
    .A3(_12569_),
    .A4(_12535_),
    .B1(_12572_),
    .X(_12573_));
 sky130_fd_sc_hd__or4_2 _16609_ (.A(_10594_),
    .B(_10598_),
    .C(_10588_),
    .D(_12540_),
    .X(_12574_));
 sky130_fd_sc_hd__buf_1 _16610_ (.A(_12574_),
    .X(_12575_));
 sky130_fd_sc_hd__buf_1 _16611_ (.A(_12575_),
    .X(_12576_));
 sky130_fd_sc_hd__or4_2 _16612_ (.A(_10594_),
    .B(_10598_),
    .C(_10588_),
    .D(_12511_),
    .X(_12577_));
 sky130_fd_sc_hd__buf_1 _16613_ (.A(_12577_),
    .X(_12578_));
 sky130_fd_sc_hd__buf_1 _16614_ (.A(_12578_),
    .X(_12579_));
 sky130_fd_sc_hd__buf_1 _16615_ (.A(_12579_),
    .X(_12580_));
 sky130_fd_sc_hd__and3_2 _16616_ (.A(_10593_),
    .B(_10598_),
    .C(\decode.immGen._imm_T_24[17] ),
    .X(_12581_));
 sky130_fd_sc_hd__buf_1 _16617_ (.A(_12581_),
    .X(_12582_));
 sky130_fd_sc_hd__buf_1 _16618_ (.A(_12582_),
    .X(_12583_));
 sky130_fd_sc_hd__and3_2 _16619_ (.A(_10611_),
    .B(_10618_),
    .C(_12583_),
    .X(_12584_));
 sky130_fd_sc_hd__buf_1 _16620_ (.A(_12584_),
    .X(_12585_));
 sky130_fd_sc_hd__buf_1 _16621_ (.A(_12534_),
    .X(_12586_));
 sky130_fd_sc_hd__buf_1 _16622_ (.A(_12582_),
    .X(_12587_));
 sky130_fd_sc_hd__buf_1 _16623_ (.A(_12587_),
    .X(_12588_));
 sky130_fd_sc_hd__buf_1 _16624_ (.A(_12588_),
    .X(_12589_));
 sky130_fd_sc_hd__or4_2 _16625_ (.A(_12497_),
    .B(_10610_),
    .C(_10617_),
    .D(_12488_),
    .X(_12590_));
 sky130_fd_sc_hd__buf_1 _16626_ (.A(_12590_),
    .X(_12591_));
 sky130_fd_sc_hd__nor2_2 _16627_ (.A(\decode.immGen._imm_T_24[17] ),
    .B(_10605_),
    .Y(_12592_));
 sky130_fd_sc_hd__and4_2 _16628_ (.A(_10609_),
    .B(_10616_),
    .C(_12592_),
    .D(_10593_),
    .X(_12593_));
 sky130_fd_sc_hd__buf_1 _16629_ (.A(_12593_),
    .X(_12594_));
 sky130_fd_sc_hd__buf_1 _16630_ (.A(_12594_),
    .X(_12595_));
 sky130_fd_sc_hd__a22o_2 _16631_ (.A1(\decode.regfile.registers_11[0] ),
    .A2(_12595_),
    .B1(_12583_),
    .B2(_12551_),
    .X(_12596_));
 sky130_fd_sc_hd__nor2_2 _16632_ (.A(\decode.immGen._imm_T_24[19] ),
    .B(\decode.immGen._imm_T_24[15] ),
    .Y(_12597_));
 sky130_fd_sc_hd__and3_2 _16633_ (.A(_10609_),
    .B(_12592_),
    .C(_12597_),
    .X(_12598_));
 sky130_fd_sc_hd__buf_1 _16634_ (.A(_12598_),
    .X(_12599_));
 sky130_fd_sc_hd__buf_1 _16635_ (.A(_12599_),
    .X(_12600_));
 sky130_fd_sc_hd__or4_2 _16636_ (.A(_11016_),
    .B(_10605_),
    .C(\decode.immGen._imm_T_24[17] ),
    .D(_12509_),
    .X(_12601_));
 sky130_fd_sc_hd__buf_1 _16637_ (.A(_12601_),
    .X(_12602_));
 sky130_fd_sc_hd__buf_1 _16638_ (.A(_12602_),
    .X(_12603_));
 sky130_fd_sc_hd__buf_1 _16639_ (.A(_12592_),
    .X(_12604_));
 sky130_fd_sc_hd__and3_2 _16640_ (.A(_12592_),
    .B(_12531_),
    .C(_10592_),
    .X(_12605_));
 sky130_fd_sc_hd__buf_1 _16641_ (.A(_12605_),
    .X(_12606_));
 sky130_fd_sc_hd__buf_1 _16642_ (.A(_12606_),
    .X(_12607_));
 sky130_fd_sc_hd__a41o_2 _16643_ (.A1(\decode.regfile.registers_8[0] ),
    .A2(_10594_),
    .A3(_12550_),
    .A4(_12604_),
    .B1(_12607_),
    .X(_12608_));
 sky130_fd_sc_hd__and4_2 _16644_ (.A(_10607_),
    .B(_10614_),
    .C(_12522_),
    .D(_10591_),
    .X(_12609_));
 sky130_fd_sc_hd__buf_1 _16645_ (.A(_12609_),
    .X(_12610_));
 sky130_fd_sc_hd__buf_1 _16646_ (.A(_12610_),
    .X(_12611_));
 sky130_fd_sc_hd__buf_1 _16647_ (.A(_12611_),
    .X(_12612_));
 sky130_fd_sc_hd__or3_2 _16648_ (.A(\decode.immGen._imm_T_24[19] ),
    .B(_10597_),
    .C(_10934_),
    .X(_12613_));
 sky130_fd_sc_hd__buf_1 _16649_ (.A(_12613_),
    .X(_12614_));
 sky130_fd_sc_hd__buf_1 _16650_ (.A(_12614_),
    .X(_12615_));
 sky130_fd_sc_hd__buf_1 _16651_ (.A(_10591_),
    .X(_12616_));
 sky130_fd_sc_hd__and3_2 _16652_ (.A(_12522_),
    .B(_12616_),
    .C(_12547_),
    .X(_12617_));
 sky130_fd_sc_hd__buf_1 _16653_ (.A(_12617_),
    .X(_12618_));
 sky130_fd_sc_hd__and3_2 _16654_ (.A(_12522_),
    .B(_12530_),
    .C(_12616_),
    .X(_12619_));
 sky130_fd_sc_hd__buf_1 _16655_ (.A(_12619_),
    .X(_12620_));
 sky130_fd_sc_hd__and3_2 _16656_ (.A(_10607_),
    .B(_12522_),
    .C(_12597_),
    .X(_12621_));
 sky130_fd_sc_hd__buf_1 _16657_ (.A(_12621_),
    .X(_12622_));
 sky130_fd_sc_hd__buf_1 _16658_ (.A(_12622_),
    .X(_12623_));
 sky130_fd_sc_hd__a221o_2 _16659_ (.A1(\decode.regfile.registers_4[0] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[0] ),
    .C1(_12623_),
    .X(_12624_));
 sky130_fd_sc_hd__buf_1 _16660_ (.A(_12613_),
    .X(_12625_));
 sky130_fd_sc_hd__buf_1 _16661_ (.A(_12625_),
    .X(_12626_));
 sky130_fd_sc_hd__nand4_2 _16662_ (.A(_10607_),
    .B(_10614_),
    .C(_12557_),
    .D(_10591_),
    .Y(_12627_));
 sky130_fd_sc_hd__buf_1 _16663_ (.A(_12627_),
    .X(_12628_));
 sky130_fd_sc_hd__buf_1 _16664_ (.A(_12628_),
    .X(_12629_));
 sky130_fd_sc_hd__nand4_2 _16665_ (.A(_12556_),
    .B(_10601_),
    .C(_10591_),
    .D(_10614_),
    .Y(_12630_));
 sky130_fd_sc_hd__buf_1 _16666_ (.A(_12630_),
    .X(_12631_));
 sky130_fd_sc_hd__mux2_2 _16667_ (.A0(\decode.regfile.registers_1[0] ),
    .A1(\decode.regfile.registers_0[0] ),
    .S(_12631_),
    .X(_12632_));
 sky130_fd_sc_hd__nand4_2 _16668_ (.A(_12597_),
    .B(_10934_),
    .C(_10605_),
    .D(_10607_),
    .Y(_12633_));
 sky130_fd_sc_hd__buf_1 _16669_ (.A(_12633_),
    .X(_12634_));
 sky130_fd_sc_hd__nor3_2 _16670_ (.A(_11016_),
    .B(_10597_),
    .C(\decode.immGen._imm_T_24[17] ),
    .Y(_12635_));
 sky130_fd_sc_hd__buf_1 _16671_ (.A(_12635_),
    .X(_12636_));
 sky130_fd_sc_hd__nand2_2 _16672_ (.A(\decode.immGen._imm_T_24[16] ),
    .B(_10614_),
    .Y(_12637_));
 sky130_fd_sc_hd__nor4_2 _16673_ (.A(_11016_),
    .B(_10597_),
    .C(\decode.immGen._imm_T_24[17] ),
    .D(_12637_),
    .Y(_12638_));
 sky130_fd_sc_hd__buf_1 _16674_ (.A(_12638_),
    .X(_12639_));
 sky130_fd_sc_hd__a31o_2 _16675_ (.A1(\decode.regfile.registers_2[0] ),
    .A2(_10608_),
    .A3(_12636_),
    .B1(_12639_),
    .X(_12640_));
 sky130_fd_sc_hd__a21o_2 _16676_ (.A1(_12632_),
    .A2(_12634_),
    .B1(_12640_),
    .X(_12641_));
 sky130_fd_sc_hd__o221a_2 _16677_ (.A1(_10610_),
    .A2(_12626_),
    .B1(_12629_),
    .B2(\decode.regfile.registers_3[0] ),
    .C1(_12641_),
    .X(_12642_));
 sky130_fd_sc_hd__o32a_2 _16678_ (.A1(\decode.regfile.registers_6[0] ),
    .A2(_10603_),
    .A3(_12615_),
    .B1(_12624_),
    .B2(_12642_),
    .X(_12643_));
 sky130_fd_sc_hd__or4_2 _16679_ (.A(_11016_),
    .B(_10597_),
    .C(_10935_),
    .D(_12637_),
    .X(_12644_));
 sky130_fd_sc_hd__buf_1 _16680_ (.A(_12644_),
    .X(_12645_));
 sky130_fd_sc_hd__o32a_2 _16681_ (.A1(_12497_),
    .A2(_12539_),
    .A3(_12503_),
    .B1(\decode.regfile.registers_7[0] ),
    .B2(_12645_),
    .X(_12646_));
 sky130_fd_sc_hd__o21a_2 _16682_ (.A1(_12612_),
    .A2(_12643_),
    .B1(_12646_),
    .X(_12647_));
 sky130_fd_sc_hd__o22a_2 _16683_ (.A1(\decode.regfile.registers_9[0] ),
    .A2(_12603_),
    .B1(_12608_),
    .B2(_12647_),
    .X(_12648_));
 sky130_fd_sc_hd__buf_1 _16684_ (.A(_12637_),
    .X(_12649_));
 sky130_fd_sc_hd__buf_1 _16685_ (.A(_12649_),
    .X(_12650_));
 sky130_fd_sc_hd__or4_2 _16686_ (.A(_11016_),
    .B(_10602_),
    .C(_12508_),
    .D(_12501_),
    .X(_12651_));
 sky130_fd_sc_hd__buf_1 _16687_ (.A(_12651_),
    .X(_12652_));
 sky130_fd_sc_hd__buf_1 _16688_ (.A(_12652_),
    .X(_12653_));
 sky130_fd_sc_hd__buf_1 _16689_ (.A(_12653_),
    .X(_12654_));
 sky130_fd_sc_hd__o32a_2 _16690_ (.A1(_11019_),
    .A2(_12504_),
    .A3(_12650_),
    .B1(\decode.regfile.registers_10[0] ),
    .B2(_12654_),
    .X(_12655_));
 sky130_fd_sc_hd__o21a_2 _16691_ (.A1(_12600_),
    .A2(_12648_),
    .B1(_12655_),
    .X(_12656_));
 sky130_fd_sc_hd__or4_2 _16692_ (.A(_12497_),
    .B(_10606_),
    .C(_10935_),
    .D(_12510_),
    .X(_12657_));
 sky130_fd_sc_hd__buf_1 _16693_ (.A(_12657_),
    .X(_12658_));
 sky130_fd_sc_hd__buf_1 _16694_ (.A(_12658_),
    .X(_12659_));
 sky130_fd_sc_hd__o221a_2 _16695_ (.A1(\decode.regfile.registers_12[0] ),
    .A2(_12591_),
    .B1(_12596_),
    .B2(_12656_),
    .C1(_12659_),
    .X(_12660_));
 sky130_fd_sc_hd__and4_2 _16696_ (.A(_10598_),
    .B(_10588_),
    .C(_10610_),
    .D(_12597_),
    .X(_12661_));
 sky130_fd_sc_hd__buf_1 _16697_ (.A(_12661_),
    .X(_12662_));
 sky130_fd_sc_hd__buf_1 _16698_ (.A(_12662_),
    .X(_12663_));
 sky130_fd_sc_hd__buf_1 _16699_ (.A(_12663_),
    .X(_12664_));
 sky130_fd_sc_hd__a311o_2 _16700_ (.A1(\decode.regfile.registers_13[0] ),
    .A2(_12586_),
    .A3(_12589_),
    .B1(_12660_),
    .C1(_12664_),
    .X(_12665_));
 sky130_fd_sc_hd__buf_1 _16701_ (.A(_12650_),
    .X(_12666_));
 sky130_fd_sc_hd__buf_1 _16702_ (.A(_12666_),
    .X(_12667_));
 sky130_fd_sc_hd__or4_2 _16703_ (.A(_11018_),
    .B(_10617_),
    .C(_12488_),
    .D(_10603_),
    .X(_12668_));
 sky130_fd_sc_hd__buf_1 _16704_ (.A(_12668_),
    .X(_12669_));
 sky130_fd_sc_hd__buf_1 _16705_ (.A(_12669_),
    .X(_12670_));
 sky130_fd_sc_hd__o32a_2 _16706_ (.A1(_11021_),
    .A2(_12491_),
    .A3(_12667_),
    .B1(\decode.regfile.registers_14[0] ),
    .B2(_12670_),
    .X(_12671_));
 sky130_fd_sc_hd__and3_2 _16707_ (.A(_11019_),
    .B(_12550_),
    .C(_12559_),
    .X(_12672_));
 sky130_fd_sc_hd__buf_1 _16708_ (.A(_12672_),
    .X(_12673_));
 sky130_fd_sc_hd__buf_1 _16709_ (.A(_12673_),
    .X(_12674_));
 sky130_fd_sc_hd__a221o_2 _16710_ (.A1(\decode.regfile.registers_15[0] ),
    .A2(_12585_),
    .B1(_12665_),
    .B2(_12671_),
    .C1(_12674_),
    .X(_12675_));
 sky130_fd_sc_hd__o211a_2 _16711_ (.A1(_12576_),
    .A2(\decode.regfile.registers_16[0] ),
    .B1(_12580_),
    .C1(_12675_),
    .X(_12676_));
 sky130_fd_sc_hd__or4_2 _16712_ (.A(_10598_),
    .B(_10588_),
    .C(_12666_),
    .D(_10594_),
    .X(_12677_));
 sky130_fd_sc_hd__buf_1 _16713_ (.A(_12677_),
    .X(_12678_));
 sky130_fd_sc_hd__buf_1 _16714_ (.A(_12678_),
    .X(_12679_));
 sky130_fd_sc_hd__o221a_2 _16715_ (.A1(\decode.regfile.registers_18[0] ),
    .A2(_12566_),
    .B1(_12573_),
    .B2(_12676_),
    .C1(_12679_),
    .X(_12680_));
 sky130_fd_sc_hd__or4_2 _16716_ (.A(_10595_),
    .B(_10599_),
    .C(_10935_),
    .D(_12512_),
    .X(_12681_));
 sky130_fd_sc_hd__buf_1 _16717_ (.A(_12681_),
    .X(_12682_));
 sky130_fd_sc_hd__o221a_2 _16718_ (.A1(\decode.regfile.registers_20[0] ),
    .A2(_12545_),
    .B1(_12563_),
    .B2(_12680_),
    .C1(_12682_),
    .X(_12683_));
 sky130_fd_sc_hd__a21oi_2 _16719_ (.A1(\decode.regfile.registers_21[0] ),
    .A2(_12538_),
    .B1(_12683_),
    .Y(_12684_));
 sky130_fd_sc_hd__and4_2 _16720_ (.A(_12525_),
    .B(_11009_),
    .C(_10925_),
    .D(_12523_),
    .X(_12685_));
 sky130_fd_sc_hd__buf_1 _16721_ (.A(_12685_),
    .X(_12686_));
 sky130_fd_sc_hd__buf_1 _16722_ (.A(_12686_),
    .X(_12687_));
 sky130_fd_sc_hd__a21oi_2 _16723_ (.A1(\decode.regfile.registers_22[0] ),
    .A2(_12528_),
    .B1(_12687_),
    .Y(_12688_));
 sky130_fd_sc_hd__o21ai_2 _16724_ (.A1(_12528_),
    .A2(_12684_),
    .B1(_12688_),
    .Y(_12689_));
 sky130_fd_sc_hd__buf_1 _16725_ (.A(_12604_),
    .X(_12690_));
 sky130_fd_sc_hd__and3_2 _16726_ (.A(_11025_),
    .B(_12690_),
    .C(_10604_),
    .X(_12691_));
 sky130_fd_sc_hd__a21oi_2 _16727_ (.A1(_12521_),
    .A2(_12689_),
    .B1(_12691_),
    .Y(_12692_));
 sky130_fd_sc_hd__o22ai_2 _16728_ (.A1(_12500_),
    .A2(_12507_),
    .B1(_12517_),
    .B2(_12692_),
    .Y(_12693_));
 sky130_fd_sc_hd__or4_2 _16729_ (.A(_11012_),
    .B(_10926_),
    .C(_12500_),
    .D(_10606_),
    .X(_12694_));
 sky130_fd_sc_hd__buf_1 _16730_ (.A(_12694_),
    .X(_12695_));
 sky130_fd_sc_hd__o32a_2 _16731_ (.A1(\decode.regfile.registers_27[0] ),
    .A2(_12507_),
    .A3(_12520_),
    .B1(_12695_),
    .B2(\decode.regfile.registers_26[0] ),
    .X(_12696_));
 sky130_fd_sc_hd__and4_2 _16732_ (.A(_10933_),
    .B(_11012_),
    .C(_11015_),
    .D(_11026_),
    .X(_12697_));
 sky130_fd_sc_hd__buf_1 _16733_ (.A(_12697_),
    .X(_12698_));
 sky130_fd_sc_hd__a21o_2 _16734_ (.A1(_12693_),
    .A2(_12696_),
    .B1(_12698_),
    .X(_12699_));
 sky130_fd_sc_hd__o221a_2 _16735_ (.A1(\decode.regfile.registers_29[0] ),
    .A2(_12493_),
    .B1(_12496_),
    .B2(\decode.regfile.registers_28[0] ),
    .C1(_12699_),
    .X(_12700_));
 sky130_fd_sc_hd__buf_1 _16736_ (.A(_10928_),
    .X(_12701_));
 sky130_fd_sc_hd__or4_2 _16737_ (.A(_12701_),
    .B(_12500_),
    .C(_10606_),
    .D(_10937_),
    .X(_12702_));
 sky130_fd_sc_hd__o32a_2 _16738_ (.A1(\decode.regfile.registers_31[0] ),
    .A2(_12491_),
    .A3(_12520_),
    .B1(\decode.regfile.registers_30[0] ),
    .B2(_12702_),
    .X(_12703_));
 sky130_fd_sc_hd__o41a_2 _16739_ (.A1(_11027_),
    .A2(_11015_),
    .A3(_11012_),
    .A4(_12542_),
    .B1(_10973_),
    .X(_12704_));
 sky130_fd_sc_hd__buf_1 _16740_ (.A(_12704_),
    .X(_12705_));
 sky130_fd_sc_hd__o211a_2 _16741_ (.A1(_12487_),
    .A2(_12700_),
    .B1(_12703_),
    .C1(_12705_),
    .X(_00420_));
 sky130_fd_sc_hd__buf_1 _16742_ (.A(_12667_),
    .X(_12706_));
 sky130_fd_sc_hd__or4_2 _16743_ (.A(_10940_),
    .B(_10606_),
    .C(_10937_),
    .D(_12706_),
    .X(_12707_));
 sky130_fd_sc_hd__buf_1 _16744_ (.A(_12707_),
    .X(_12708_));
 sky130_fd_sc_hd__buf_1 _16745_ (.A(_12708_),
    .X(_12709_));
 sky130_fd_sc_hd__o21a_2 _16746_ (.A1(_10931_),
    .A2(\decode.regfile.registers_30[1] ),
    .B1(_12487_),
    .X(_12710_));
 sky130_fd_sc_hd__o21a_2 _16747_ (.A1(_10930_),
    .A2(\decode.regfile.registers_28[1] ),
    .B1(_12698_),
    .X(_12711_));
 sky130_fd_sc_hd__buf_1 _16748_ (.A(_10926_),
    .X(_12712_));
 sky130_fd_sc_hd__o2111a_2 _16749_ (.A1(_12712_),
    .A2(\decode.regfile.registers_24[1] ),
    .B1(_10604_),
    .C1(_12690_),
    .D1(_11025_),
    .X(_12713_));
 sky130_fd_sc_hd__or4_2 _16750_ (.A(_11013_),
    .B(_10935_),
    .C(_12667_),
    .D(_10595_),
    .X(_12714_));
 sky130_fd_sc_hd__o2111a_2 _16751_ (.A1(_10926_),
    .A2(\decode.regfile.registers_22[1] ),
    .B1(_12554_),
    .C1(_11009_),
    .D1(_12546_),
    .X(_12715_));
 sky130_fd_sc_hd__buf_1 _16752_ (.A(_12681_),
    .X(_12716_));
 sky130_fd_sc_hd__a41o_2 _16753_ (.A1(\decode.regfile.registers_20[1] ),
    .A2(_12525_),
    .A3(_12552_),
    .A4(_12523_),
    .B1(_12536_),
    .X(_12717_));
 sky130_fd_sc_hd__o2111a_2 _16754_ (.A1(\decode.regfile.registers_18[1] ),
    .A2(_10924_),
    .B1(_12568_),
    .C1(_12524_),
    .D1(_11008_),
    .X(_12718_));
 sky130_fd_sc_hd__buf_1 _16755_ (.A(_12578_),
    .X(_12719_));
 sky130_fd_sc_hd__a41o_2 _16756_ (.A1(\decode.regfile.registers_15[1] ),
    .A2(_10611_),
    .A3(_10618_),
    .A4(_12588_),
    .B1(_12672_),
    .X(_12720_));
 sky130_fd_sc_hd__or3_2 _16757_ (.A(_11017_),
    .B(_10606_),
    .C(_10935_),
    .X(_12721_));
 sky130_fd_sc_hd__buf_1 _16758_ (.A(_12721_),
    .X(_12722_));
 sky130_fd_sc_hd__buf_1 _16759_ (.A(_12722_),
    .X(_12723_));
 sky130_fd_sc_hd__buf_1 _16760_ (.A(_12594_),
    .X(_12724_));
 sky130_fd_sc_hd__or4_2 _16761_ (.A(_11016_),
    .B(_10608_),
    .C(_12508_),
    .D(_12502_),
    .X(_12725_));
 sky130_fd_sc_hd__buf_1 _16762_ (.A(_12725_),
    .X(_12726_));
 sky130_fd_sc_hd__a22o_2 _16763_ (.A1(\decode.regfile.registers_4[1] ),
    .A2(_12617_),
    .B1(_12619_),
    .B2(\decode.regfile.registers_5[1] ),
    .X(_12727_));
 sky130_fd_sc_hd__and3_2 _16764_ (.A(_12557_),
    .B(_10591_),
    .C(_10607_),
    .X(_12728_));
 sky130_fd_sc_hd__buf_1 _16765_ (.A(_12728_),
    .X(_12729_));
 sky130_fd_sc_hd__mux2_2 _16766_ (.A0(\decode.regfile.registers_1[1] ),
    .A1(\decode.regfile.registers_0[1] ),
    .S(_12630_),
    .X(_12730_));
 sky130_fd_sc_hd__or4_2 _16767_ (.A(\decode.immGen._imm_T_24[19] ),
    .B(_10597_),
    .C(_10607_),
    .D(_10934_),
    .X(_12731_));
 sky130_fd_sc_hd__buf_1 _16768_ (.A(_12731_),
    .X(_12732_));
 sky130_fd_sc_hd__o221a_2 _16769_ (.A1(\decode.regfile.registers_2[1] ),
    .A2(_12633_),
    .B1(_12627_),
    .B2(\decode.regfile.registers_3[1] ),
    .C1(_12732_),
    .X(_12733_));
 sky130_fd_sc_hd__o21a_2 _16770_ (.A1(_12729_),
    .A2(_12730_),
    .B1(_12733_),
    .X(_12734_));
 sky130_fd_sc_hd__or4_2 _16771_ (.A(_11016_),
    .B(_10597_),
    .C(_10935_),
    .D(_10602_),
    .X(_12735_));
 sky130_fd_sc_hd__o21ai_2 _16772_ (.A1(_12727_),
    .A2(_12734_),
    .B1(_12735_),
    .Y(_12736_));
 sky130_fd_sc_hd__buf_1 _16773_ (.A(_12621_),
    .X(_12737_));
 sky130_fd_sc_hd__a22oi_2 _16774_ (.A1(\decode.regfile.registers_7[1] ),
    .A2(_12610_),
    .B1(_12737_),
    .B2(\decode.regfile.registers_6[1] ),
    .Y(_12738_));
 sky130_fd_sc_hd__nand2_2 _16775_ (.A(_12736_),
    .B(_12738_),
    .Y(_12739_));
 sky130_fd_sc_hd__a41o_2 _16776_ (.A1(\decode.regfile.registers_8[1] ),
    .A2(_10593_),
    .A3(_12549_),
    .A4(_12592_),
    .B1(_12605_),
    .X(_12740_));
 sky130_fd_sc_hd__a21o_2 _16777_ (.A1(_12726_),
    .A2(_12739_),
    .B1(_12740_),
    .X(_12741_));
 sky130_fd_sc_hd__o41a_2 _16778_ (.A1(\decode.regfile.registers_9[1] ),
    .A2(_12497_),
    .A3(_12503_),
    .A4(_12510_),
    .B1(_12652_),
    .X(_12742_));
 sky130_fd_sc_hd__a22oi_2 _16779_ (.A1(\decode.regfile.registers_10[1] ),
    .A2(_12599_),
    .B1(_12741_),
    .B2(_12742_),
    .Y(_12743_));
 sky130_fd_sc_hd__or4b_2 _16780_ (.A(_12497_),
    .B(_12503_),
    .C(_12637_),
    .D_N(\decode.regfile.registers_11[1] ),
    .X(_12744_));
 sky130_fd_sc_hd__buf_1 _16781_ (.A(_12590_),
    .X(_12745_));
 sky130_fd_sc_hd__o211ai_2 _16782_ (.A1(_12724_),
    .A2(_12743_),
    .B1(_12744_),
    .C1(_12745_),
    .Y(_12746_));
 sky130_fd_sc_hd__or4_2 _16783_ (.A(\decode.regfile.registers_12[1] ),
    .B(_12489_),
    .C(_12498_),
    .D(_12540_),
    .X(_12747_));
 sky130_fd_sc_hd__a31o_2 _16784_ (.A1(\decode.regfile.registers_13[1] ),
    .A2(_12533_),
    .A3(_12582_),
    .B1(_12662_),
    .X(_12748_));
 sky130_fd_sc_hd__a31o_2 _16785_ (.A1(_12658_),
    .A2(_12746_),
    .A3(_12747_),
    .B1(_12748_),
    .X(_12749_));
 sky130_fd_sc_hd__o221a_2 _16786_ (.A1(_12650_),
    .A2(_12723_),
    .B1(_12669_),
    .B2(\decode.regfile.registers_14[1] ),
    .C1(_12749_),
    .X(_12750_));
 sky130_fd_sc_hd__o22a_2 _16787_ (.A1(\decode.regfile.registers_16[1] ),
    .A2(_12575_),
    .B1(_12720_),
    .B2(_12750_),
    .X(_12751_));
 sky130_fd_sc_hd__a31o_2 _16788_ (.A1(_11022_),
    .A2(_12567_),
    .A3(_12586_),
    .B1(_12751_),
    .X(_12752_));
 sky130_fd_sc_hd__o211a_2 _16789_ (.A1(\decode.regfile.registers_17[1] ),
    .A2(_12719_),
    .B1(_12565_),
    .C1(_12752_),
    .X(_12753_));
 sky130_fd_sc_hd__o221a_2 _16790_ (.A1(\decode.regfile.registers_19[1] ),
    .A2(_12678_),
    .B1(_12718_),
    .B2(_12753_),
    .C1(_12544_),
    .X(_12754_));
 sky130_fd_sc_hd__or4_2 _16791_ (.A(_10599_),
    .B(_10924_),
    .C(_12500_),
    .D(_10935_),
    .X(_12755_));
 sky130_fd_sc_hd__o221a_2 _16792_ (.A1(\decode.regfile.registers_21[1] ),
    .A2(_12716_),
    .B1(_12717_),
    .B2(_12754_),
    .C1(_12755_),
    .X(_12756_));
 sky130_fd_sc_hd__o221a_2 _16793_ (.A1(\decode.regfile.registers_23[1] ),
    .A2(_12714_),
    .B1(_12715_),
    .B2(_12756_),
    .C1(_12514_),
    .X(_12757_));
 sky130_fd_sc_hd__o221a_2 _16794_ (.A1(_12513_),
    .A2(\decode.regfile.registers_25[1] ),
    .B1(_12713_),
    .B2(_12757_),
    .C1(_12694_),
    .X(_12758_));
 sky130_fd_sc_hd__buf_1 _16795_ (.A(_12690_),
    .X(_12759_));
 sky130_fd_sc_hd__o2111a_2 _16796_ (.A1(_12494_),
    .A2(\decode.regfile.registers_26[1] ),
    .B1(_12759_),
    .C1(_11010_),
    .D1(_11026_),
    .X(_12760_));
 sky130_fd_sc_hd__or2_2 _16797_ (.A(_12758_),
    .B(_12760_),
    .X(_12761_));
 sky130_fd_sc_hd__o311a_2 _16798_ (.A1(\decode.regfile.registers_27[1] ),
    .A2(_12507_),
    .A3(_12520_),
    .B1(_12495_),
    .C1(_12761_),
    .X(_12762_));
 sky130_fd_sc_hd__o221a_2 _16799_ (.A1(_12492_),
    .A2(\decode.regfile.registers_29[1] ),
    .B1(_12711_),
    .B2(_12762_),
    .C1(_12702_),
    .X(_12763_));
 sky130_fd_sc_hd__o221a_2 _16800_ (.A1(\decode.regfile.registers_31[1] ),
    .A2(_12709_),
    .B1(_12710_),
    .B2(_12763_),
    .C1(_12705_),
    .X(_00421_));
 sky130_fd_sc_hd__o21a_2 _16801_ (.A1(_10931_),
    .A2(\decode.regfile.registers_30[2] ),
    .B1(_12487_),
    .X(_12764_));
 sky130_fd_sc_hd__buf_1 _16802_ (.A(_10930_),
    .X(_12765_));
 sky130_fd_sc_hd__or4_2 _16803_ (.A(_10939_),
    .B(_10606_),
    .C(_10937_),
    .D(_10933_),
    .X(_12766_));
 sky130_fd_sc_hd__buf_1 _16804_ (.A(_12766_),
    .X(_12767_));
 sky130_fd_sc_hd__buf_1 _16805_ (.A(_12767_),
    .X(_12768_));
 sky130_fd_sc_hd__o21ai_2 _16806_ (.A1(\decode.regfile.registers_23[2] ),
    .A2(_12714_),
    .B1(_12515_),
    .Y(_12769_));
 sky130_fd_sc_hd__and3_2 _16807_ (.A(_12524_),
    .B(_12551_),
    .C(_12523_),
    .X(_12770_));
 sky130_fd_sc_hd__buf_1 _16808_ (.A(_12770_),
    .X(_12771_));
 sky130_fd_sc_hd__buf_1 _16809_ (.A(_12722_),
    .X(_12772_));
 sky130_fd_sc_hd__buf_1 _16810_ (.A(_12772_),
    .X(_12773_));
 sky130_fd_sc_hd__and3_2 _16811_ (.A(_12582_),
    .B(_10603_),
    .C(_10617_),
    .X(_12774_));
 sky130_fd_sc_hd__buf_1 _16812_ (.A(_12774_),
    .X(_12775_));
 sky130_fd_sc_hd__buf_1 _16813_ (.A(_10593_),
    .X(_12776_));
 sky130_fd_sc_hd__a41o_2 _16814_ (.A1(\decode.regfile.registers_8[2] ),
    .A2(_12776_),
    .A3(_12550_),
    .A4(_12604_),
    .B1(_12607_),
    .X(_12777_));
 sky130_fd_sc_hd__buf_1 _16815_ (.A(_12630_),
    .X(_12778_));
 sky130_fd_sc_hd__a31o_2 _16816_ (.A1(_12531_),
    .A2(_10592_),
    .A3(_12558_),
    .B1(\decode.regfile.registers_0[2] ),
    .X(_12779_));
 sky130_fd_sc_hd__o211ai_2 _16817_ (.A1(\decode.regfile.registers_1[2] ),
    .A2(_12778_),
    .B1(_12634_),
    .C1(_12779_),
    .Y(_12780_));
 sky130_fd_sc_hd__o21ai_2 _16818_ (.A1(\decode.regfile.registers_2[2] ),
    .A2(_10616_),
    .B1(_12729_),
    .Y(_12781_));
 sky130_fd_sc_hd__o21ai_2 _16819_ (.A1(\decode.regfile.registers_3[2] ),
    .A2(_12629_),
    .B1(_12732_),
    .Y(_12782_));
 sky130_fd_sc_hd__a21oi_2 _16820_ (.A1(_12780_),
    .A2(_12781_),
    .B1(_12782_),
    .Y(_12783_));
 sky130_fd_sc_hd__a221o_2 _16821_ (.A1(\decode.regfile.registers_4[2] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[2] ),
    .C1(_12737_),
    .X(_12784_));
 sky130_fd_sc_hd__o32a_2 _16822_ (.A1(\decode.regfile.registers_6[2] ),
    .A2(_10602_),
    .A3(_12615_),
    .B1(_12783_),
    .B2(_12784_),
    .X(_12785_));
 sky130_fd_sc_hd__o32a_2 _16823_ (.A1(_12497_),
    .A2(_12539_),
    .A3(_12503_),
    .B1(\decode.regfile.registers_7[2] ),
    .B2(_12645_),
    .X(_12786_));
 sky130_fd_sc_hd__o21a_2 _16824_ (.A1(_12612_),
    .A2(_12785_),
    .B1(_12786_),
    .X(_12787_));
 sky130_fd_sc_hd__o22ai_2 _16825_ (.A1(\decode.regfile.registers_9[2] ),
    .A2(_12603_),
    .B1(_12777_),
    .B2(_12787_),
    .Y(_12788_));
 sky130_fd_sc_hd__nand2_2 _16826_ (.A(_12654_),
    .B(_12788_),
    .Y(_12789_));
 sky130_fd_sc_hd__buf_1 _16827_ (.A(_12652_),
    .X(_12790_));
 sky130_fd_sc_hd__or4_2 _16828_ (.A(_11017_),
    .B(_10588_),
    .C(_12637_),
    .D(_10605_),
    .X(_12791_));
 sky130_fd_sc_hd__buf_1 _16829_ (.A(_12791_),
    .X(_12792_));
 sky130_fd_sc_hd__o21a_2 _16830_ (.A1(\decode.regfile.registers_10[2] ),
    .A2(_12790_),
    .B1(_12792_),
    .X(_12793_));
 sky130_fd_sc_hd__and4_2 _16831_ (.A(_10598_),
    .B(_10588_),
    .C(_12549_),
    .D(_12776_),
    .X(_12794_));
 sky130_fd_sc_hd__a221o_2 _16832_ (.A1(\decode.regfile.registers_11[2] ),
    .A2(_12595_),
    .B1(_12789_),
    .B2(_12793_),
    .C1(_12794_),
    .X(_12795_));
 sky130_fd_sc_hd__o32a_2 _16833_ (.A1(_11020_),
    .A2(_12490_),
    .A3(_12512_),
    .B1(\decode.regfile.registers_12[2] ),
    .B2(_12591_),
    .X(_12796_));
 sky130_fd_sc_hd__a221o_2 _16834_ (.A1(\decode.regfile.registers_13[2] ),
    .A2(_12775_),
    .B1(_12795_),
    .B2(_12796_),
    .C1(_12664_),
    .X(_12797_));
 sky130_fd_sc_hd__o221a_2 _16835_ (.A1(_12667_),
    .A2(_12773_),
    .B1(_12670_),
    .B2(\decode.regfile.registers_14[2] ),
    .C1(_12797_),
    .X(_12798_));
 sky130_fd_sc_hd__a211o_2 _16836_ (.A1(\decode.regfile.registers_15[2] ),
    .A2(_12585_),
    .B1(_12674_),
    .C1(_12798_),
    .X(_12799_));
 sky130_fd_sc_hd__o21ai_2 _16837_ (.A1(\decode.regfile.registers_16[2] ),
    .A2(_12576_),
    .B1(_12799_),
    .Y(_12800_));
 sky130_fd_sc_hd__o21ai_2 _16838_ (.A1(\decode.regfile.registers_17[2] ),
    .A2(_12580_),
    .B1(_12566_),
    .Y(_12801_));
 sky130_fd_sc_hd__a21oi_2 _16839_ (.A1(_12580_),
    .A2(_12800_),
    .B1(_12801_),
    .Y(_12802_));
 sky130_fd_sc_hd__a211o_2 _16840_ (.A1(\decode.regfile.registers_18[2] ),
    .A2(_12572_),
    .B1(_12562_),
    .C1(_12802_),
    .X(_12803_));
 sky130_fd_sc_hd__o41a_2 _16841_ (.A1(\decode.regfile.registers_19[2] ),
    .A2(_11013_),
    .A3(_11012_),
    .A4(_12519_),
    .B1(_12545_),
    .X(_12804_));
 sky130_fd_sc_hd__a221o_2 _16842_ (.A1(\decode.regfile.registers_20[2] ),
    .A2(_12771_),
    .B1(_12803_),
    .B2(_12804_),
    .C1(_12538_),
    .X(_12805_));
 sky130_fd_sc_hd__buf_1 _16843_ (.A(_12755_),
    .X(_12806_));
 sky130_fd_sc_hd__o21a_2 _16844_ (.A1(\decode.regfile.registers_21[2] ),
    .A2(_12682_),
    .B1(_12806_),
    .X(_12807_));
 sky130_fd_sc_hd__a221oi_2 _16845_ (.A1(\decode.regfile.registers_22[2] ),
    .A2(_12528_),
    .B1(_12805_),
    .B2(_12807_),
    .C1(_12687_),
    .Y(_12808_));
 sky130_fd_sc_hd__o21ai_2 _16846_ (.A1(_12494_),
    .A2(\decode.regfile.registers_24[2] ),
    .B1(_12691_),
    .Y(_12809_));
 sky130_fd_sc_hd__o21ai_2 _16847_ (.A1(_12769_),
    .A2(_12808_),
    .B1(_12809_),
    .Y(_12810_));
 sky130_fd_sc_hd__buf_1 _16848_ (.A(_12512_),
    .X(_12811_));
 sky130_fd_sc_hd__buf_1 _16849_ (.A(_12811_),
    .X(_12812_));
 sky130_fd_sc_hd__or4_2 _16850_ (.A(_10939_),
    .B(\decode.regfile.registers_25[2] ),
    .C(_12506_),
    .D(_12812_),
    .X(_12813_));
 sky130_fd_sc_hd__buf_1 _16851_ (.A(_12759_),
    .X(_12814_));
 sky130_fd_sc_hd__o2111a_2 _16852_ (.A1(_10928_),
    .A2(\decode.regfile.registers_26[2] ),
    .B1(_12814_),
    .C1(_11011_),
    .D1(_11027_),
    .X(_12815_));
 sky130_fd_sc_hd__a31o_2 _16853_ (.A1(_12695_),
    .A2(_12810_),
    .A3(_12813_),
    .B1(_12815_),
    .X(_12816_));
 sky130_fd_sc_hd__or4_2 _16854_ (.A(_10940_),
    .B(_12706_),
    .C(\decode.regfile.registers_27[2] ),
    .D(_12507_),
    .X(_12817_));
 sky130_fd_sc_hd__o21a_2 _16855_ (.A1(_12701_),
    .A2(\decode.regfile.registers_28[2] ),
    .B1(_12698_),
    .X(_12818_));
 sky130_fd_sc_hd__a31o_2 _16856_ (.A1(_12496_),
    .A2(_12816_),
    .A3(_12817_),
    .B1(_12818_),
    .X(_12819_));
 sky130_fd_sc_hd__o221a_2 _16857_ (.A1(_12765_),
    .A2(_12768_),
    .B1(_12493_),
    .B2(\decode.regfile.registers_29[2] ),
    .C1(_12819_),
    .X(_12820_));
 sky130_fd_sc_hd__o221a_2 _16858_ (.A1(\decode.regfile.registers_31[2] ),
    .A2(_12709_),
    .B1(_12764_),
    .B2(_12820_),
    .C1(_12705_),
    .X(_00422_));
 sky130_fd_sc_hd__o21a_2 _16859_ (.A1(_10931_),
    .A2(\decode.regfile.registers_30[3] ),
    .B1(_12487_),
    .X(_12821_));
 sky130_fd_sc_hd__buf_1 _16860_ (.A(_12681_),
    .X(_12822_));
 sky130_fd_sc_hd__buf_1 _16861_ (.A(_12523_),
    .X(_12823_));
 sky130_fd_sc_hd__buf_1 _16862_ (.A(_12536_),
    .X(_12824_));
 sky130_fd_sc_hd__a41o_2 _16863_ (.A1(\decode.regfile.registers_20[3] ),
    .A2(_11024_),
    .A3(_12553_),
    .A4(_12823_),
    .B1(_12824_),
    .X(_12825_));
 sky130_fd_sc_hd__buf_1 _16864_ (.A(_12564_),
    .X(_12826_));
 sky130_fd_sc_hd__a41o_2 _16865_ (.A1(\decode.regfile.registers_17[3] ),
    .A2(_11022_),
    .A3(_12567_),
    .A4(_12586_),
    .B1(_12570_),
    .X(_12827_));
 sky130_fd_sc_hd__a31o_2 _16866_ (.A1(\decode.regfile.registers_13[3] ),
    .A2(_12533_),
    .A3(_12587_),
    .B1(_12662_),
    .X(_12828_));
 sky130_fd_sc_hd__nand4_2 _16867_ (.A(_10591_),
    .B(_10605_),
    .C(_10934_),
    .D(_10607_),
    .Y(_12829_));
 sky130_fd_sc_hd__buf_1 _16868_ (.A(_12829_),
    .X(_12830_));
 sky130_fd_sc_hd__mux2_2 _16869_ (.A0(\decode.regfile.registers_1[3] ),
    .A1(\decode.regfile.registers_0[3] ),
    .S(_12631_),
    .X(_12831_));
 sky130_fd_sc_hd__nand2_2 _16870_ (.A(_12830_),
    .B(_12831_),
    .Y(_12832_));
 sky130_fd_sc_hd__and4_2 _16871_ (.A(_12597_),
    .B(_10934_),
    .C(_10605_),
    .D(_10607_),
    .X(_12833_));
 sky130_fd_sc_hd__buf_1 _16872_ (.A(_12833_),
    .X(_12834_));
 sky130_fd_sc_hd__buf_1 _16873_ (.A(_12834_),
    .X(_12835_));
 sky130_fd_sc_hd__buf_1 _16874_ (.A(_12638_),
    .X(_12836_));
 sky130_fd_sc_hd__and3_2 _16875_ (.A(_12522_),
    .B(_10601_),
    .C(_10591_),
    .X(_12837_));
 sky130_fd_sc_hd__buf_1 _16876_ (.A(_12837_),
    .X(_12838_));
 sky130_fd_sc_hd__a221oi_2 _16877_ (.A1(\decode.regfile.registers_2[3] ),
    .A2(_12835_),
    .B1(_12836_),
    .B2(\decode.regfile.registers_3[3] ),
    .C1(_12838_),
    .Y(_12839_));
 sky130_fd_sc_hd__a221o_2 _16878_ (.A1(\decode.regfile.registers_4[3] ),
    .A2(_12548_),
    .B1(_12531_),
    .B2(\decode.regfile.registers_5[3] ),
    .C1(_12625_),
    .X(_12840_));
 sky130_fd_sc_hd__a21bo_2 _16879_ (.A1(_12832_),
    .A2(_12839_),
    .B1_N(_12840_),
    .X(_12841_));
 sky130_fd_sc_hd__and3_2 _16880_ (.A(_12592_),
    .B(_12616_),
    .C(_12547_),
    .X(_12842_));
 sky130_fd_sc_hd__buf_1 _16881_ (.A(_12842_),
    .X(_12843_));
 sky130_fd_sc_hd__a221oi_2 _16882_ (.A1(\decode.regfile.registers_7[3] ),
    .A2(_12610_),
    .B1(_12737_),
    .B2(\decode.regfile.registers_6[3] ),
    .C1(_12843_),
    .Y(_12844_));
 sky130_fd_sc_hd__nand2_2 _16883_ (.A(_12841_),
    .B(_12844_),
    .Y(_12845_));
 sky130_fd_sc_hd__o32a_2 _16884_ (.A1(_11017_),
    .A2(_12502_),
    .A3(_12509_),
    .B1(\decode.regfile.registers_8[3] ),
    .B2(_12725_),
    .X(_12846_));
 sky130_fd_sc_hd__a22oi_2 _16885_ (.A1(\decode.regfile.registers_9[3] ),
    .A2(_12606_),
    .B1(_12845_),
    .B2(_12846_),
    .Y(_12847_));
 sky130_fd_sc_hd__o21ai_2 _16886_ (.A1(\decode.regfile.registers_10[3] ),
    .A2(_12652_),
    .B1(_12791_),
    .Y(_12848_));
 sky130_fd_sc_hd__a21oi_2 _16887_ (.A1(_12847_),
    .A2(_12653_),
    .B1(_12848_),
    .Y(_12849_));
 sky130_fd_sc_hd__a221o_2 _16888_ (.A1(\decode.regfile.registers_11[3] ),
    .A2(_12594_),
    .B1(_12582_),
    .B2(_12550_),
    .C1(_12849_),
    .X(_12850_));
 sky130_fd_sc_hd__o311a_2 _16889_ (.A1(\decode.regfile.registers_12[3] ),
    .A2(_12541_),
    .A3(_12722_),
    .B1(_12658_),
    .C1(_12850_),
    .X(_12851_));
 sky130_fd_sc_hd__or4_2 _16890_ (.A(_11019_),
    .B(_10606_),
    .C(_10935_),
    .D(_12649_),
    .X(_12852_));
 sky130_fd_sc_hd__o221a_2 _16891_ (.A1(\decode.regfile.registers_14[3] ),
    .A2(_12669_),
    .B1(_12828_),
    .B2(_12851_),
    .C1(_12852_),
    .X(_12853_));
 sky130_fd_sc_hd__a211o_2 _16892_ (.A1(\decode.regfile.registers_15[3] ),
    .A2(_12584_),
    .B1(_12673_),
    .C1(_12853_),
    .X(_12854_));
 sky130_fd_sc_hd__o211a_2 _16893_ (.A1(\decode.regfile.registers_16[3] ),
    .A2(_12576_),
    .B1(_12579_),
    .C1(_12854_),
    .X(_12855_));
 sky130_fd_sc_hd__o22a_2 _16894_ (.A1(\decode.regfile.registers_18[3] ),
    .A2(_12826_),
    .B1(_12827_),
    .B2(_12855_),
    .X(_12856_));
 sky130_fd_sc_hd__or4_2 _16895_ (.A(\decode.regfile.registers_19[3] ),
    .B(_10599_),
    .C(_10589_),
    .D(_12518_),
    .X(_12857_));
 sky130_fd_sc_hd__o211a_2 _16896_ (.A1(_12562_),
    .A2(_12856_),
    .B1(_12857_),
    .C1(_12545_),
    .X(_12858_));
 sky130_fd_sc_hd__o221a_2 _16897_ (.A1(\decode.regfile.registers_21[3] ),
    .A2(_12822_),
    .B1(_12825_),
    .B2(_12858_),
    .C1(_12806_),
    .X(_12859_));
 sky130_fd_sc_hd__a211o_2 _16898_ (.A1(\decode.regfile.registers_22[3] ),
    .A2(_12528_),
    .B1(_12859_),
    .C1(_12687_),
    .X(_12860_));
 sky130_fd_sc_hd__or4_2 _16899_ (.A(_11015_),
    .B(_10937_),
    .C(\decode.regfile.registers_23[3] ),
    .D(_12520_),
    .X(_12861_));
 sky130_fd_sc_hd__buf_1 _16900_ (.A(_12546_),
    .X(_12862_));
 sky130_fd_sc_hd__o2111a_2 _16901_ (.A1(_10927_),
    .A2(\decode.regfile.registers_24[3] ),
    .B1(_10933_),
    .C1(_12759_),
    .D1(_12862_),
    .X(_12863_));
 sky130_fd_sc_hd__a31o_2 _16902_ (.A1(_12516_),
    .A2(_12860_),
    .A3(_12861_),
    .B1(_12863_),
    .X(_12864_));
 sky130_fd_sc_hd__or4_2 _16903_ (.A(_10939_),
    .B(\decode.regfile.registers_25[3] ),
    .C(_12506_),
    .D(_12812_),
    .X(_12865_));
 sky130_fd_sc_hd__o2111a_2 _16904_ (.A1(_10928_),
    .A2(\decode.regfile.registers_26[3] ),
    .B1(_12814_),
    .C1(_11011_),
    .D1(_11027_),
    .X(_12866_));
 sky130_fd_sc_hd__a31o_2 _16905_ (.A1(_12695_),
    .A2(_12864_),
    .A3(_12865_),
    .B1(_12866_),
    .X(_12867_));
 sky130_fd_sc_hd__or4_2 _16906_ (.A(_10940_),
    .B(_12706_),
    .C(\decode.regfile.registers_27[3] ),
    .D(_12507_),
    .X(_12868_));
 sky130_fd_sc_hd__o21a_2 _16907_ (.A1(_12701_),
    .A2(\decode.regfile.registers_28[3] ),
    .B1(_12698_),
    .X(_12869_));
 sky130_fd_sc_hd__a31o_2 _16908_ (.A1(_12496_),
    .A2(_12867_),
    .A3(_12868_),
    .B1(_12869_),
    .X(_12870_));
 sky130_fd_sc_hd__o221a_2 _16909_ (.A1(_12765_),
    .A2(_12768_),
    .B1(_12493_),
    .B2(\decode.regfile.registers_29[3] ),
    .C1(_12870_),
    .X(_12871_));
 sky130_fd_sc_hd__o221a_2 _16910_ (.A1(\decode.regfile.registers_31[3] ),
    .A2(_12709_),
    .B1(_12821_),
    .B2(_12871_),
    .C1(_12705_),
    .X(_00423_));
 sky130_fd_sc_hd__buf_1 _16911_ (.A(_12707_),
    .X(_12872_));
 sky130_fd_sc_hd__o21a_2 _16912_ (.A1(_10931_),
    .A2(\decode.regfile.registers_30[4] ),
    .B1(_12487_),
    .X(_12873_));
 sky130_fd_sc_hd__buf_1 _16913_ (.A(_12852_),
    .X(_12874_));
 sky130_fd_sc_hd__o211a_2 _16914_ (.A1(\decode.regfile.registers_14[4] ),
    .A2(_10924_),
    .B1(_12589_),
    .C1(_10612_),
    .X(_12875_));
 sky130_fd_sc_hd__buf_1 _16915_ (.A(_12583_),
    .X(_12876_));
 sky130_fd_sc_hd__a22o_2 _16916_ (.A1(\decode.regfile.registers_11[4] ),
    .A2(_12595_),
    .B1(_12876_),
    .B2(_12551_),
    .X(_12877_));
 sky130_fd_sc_hd__buf_1 _16917_ (.A(_12791_),
    .X(_12878_));
 sky130_fd_sc_hd__or3_2 _16918_ (.A(_10602_),
    .B(_12508_),
    .C(_12613_),
    .X(_12879_));
 sky130_fd_sc_hd__buf_1 _16919_ (.A(_12879_),
    .X(_12880_));
 sky130_fd_sc_hd__a221oi_2 _16920_ (.A1(\decode.regfile.registers_4[4] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[4] ),
    .C1(_12623_),
    .Y(_12881_));
 sky130_fd_sc_hd__buf_1 _16921_ (.A(_12508_),
    .X(_12882_));
 sky130_fd_sc_hd__a31o_2 _16922_ (.A1(_12531_),
    .A2(_10592_),
    .A3(_12558_),
    .B1(\decode.regfile.registers_0[4] ),
    .X(_12883_));
 sky130_fd_sc_hd__o221a_2 _16923_ (.A1(\decode.regfile.registers_1[4] ),
    .A2(_12778_),
    .B1(_12830_),
    .B2(_12882_),
    .C1(_12883_),
    .X(_12884_));
 sky130_fd_sc_hd__a211o_2 _16924_ (.A1(\decode.regfile.registers_2[4] ),
    .A2(_12835_),
    .B1(_12836_),
    .C1(_12884_),
    .X(_12885_));
 sky130_fd_sc_hd__o221ai_2 _16925_ (.A1(_10610_),
    .A2(_12615_),
    .B1(_12629_),
    .B2(\decode.regfile.registers_3[4] ),
    .C1(_12885_),
    .Y(_12886_));
 sky130_fd_sc_hd__a2bb2o_2 _16926_ (.A1_N(\decode.regfile.registers_6[4] ),
    .A2_N(_12880_),
    .B1(_12881_),
    .B2(_12886_),
    .X(_12887_));
 sky130_fd_sc_hd__buf_1 _16927_ (.A(_12843_),
    .X(_12888_));
 sky130_fd_sc_hd__buf_1 _16928_ (.A(_12888_),
    .X(_12889_));
 sky130_fd_sc_hd__a21oi_2 _16929_ (.A1(\decode.regfile.registers_7[4] ),
    .A2(_12612_),
    .B1(_12889_),
    .Y(_12890_));
 sky130_fd_sc_hd__o21ai_2 _16930_ (.A1(_12612_),
    .A2(_12887_),
    .B1(_12890_),
    .Y(_12891_));
 sky130_fd_sc_hd__buf_1 _16931_ (.A(_12726_),
    .X(_12892_));
 sky130_fd_sc_hd__o32a_2 _16932_ (.A1(_11019_),
    .A2(_12504_),
    .A3(_12511_),
    .B1(\decode.regfile.registers_8[4] ),
    .B2(_12892_),
    .X(_12893_));
 sky130_fd_sc_hd__a221o_2 _16933_ (.A1(\decode.regfile.registers_9[4] ),
    .A2(_12607_),
    .B1(_12891_),
    .B2(_12893_),
    .C1(_12600_),
    .X(_12894_));
 sky130_fd_sc_hd__o211a_2 _16934_ (.A1(\decode.regfile.registers_10[4] ),
    .A2(_12654_),
    .B1(_12878_),
    .C1(_12894_),
    .X(_12895_));
 sky130_fd_sc_hd__o22ai_2 _16935_ (.A1(\decode.regfile.registers_12[4] ),
    .A2(_12591_),
    .B1(_12877_),
    .B2(_12895_),
    .Y(_12896_));
 sky130_fd_sc_hd__o21ai_2 _16936_ (.A1(\decode.regfile.registers_13[4] ),
    .A2(_12659_),
    .B1(_12670_),
    .Y(_12897_));
 sky130_fd_sc_hd__a21oi_2 _16937_ (.A1(_12659_),
    .A2(_12896_),
    .B1(_12897_),
    .Y(_12898_));
 sky130_fd_sc_hd__o22ai_2 _16938_ (.A1(\decode.regfile.registers_15[4] ),
    .A2(_12874_),
    .B1(_12875_),
    .B2(_12898_),
    .Y(_12899_));
 sky130_fd_sc_hd__and3_2 _16939_ (.A(_11020_),
    .B(_12559_),
    .C(_12534_),
    .X(_12900_));
 sky130_fd_sc_hd__buf_1 _16940_ (.A(_12900_),
    .X(_12901_));
 sky130_fd_sc_hd__a21oi_2 _16941_ (.A1(\decode.regfile.registers_16[4] ),
    .A2(_12674_),
    .B1(_12901_),
    .Y(_12902_));
 sky130_fd_sc_hd__o21ai_2 _16942_ (.A1(_12674_),
    .A2(_12899_),
    .B1(_12902_),
    .Y(_12903_));
 sky130_fd_sc_hd__o21a_2 _16943_ (.A1(\decode.regfile.registers_17[4] ),
    .A2(_12719_),
    .B1(_12826_),
    .X(_12904_));
 sky130_fd_sc_hd__a221o_2 _16944_ (.A1(\decode.regfile.registers_18[4] ),
    .A2(_12572_),
    .B1(_12903_),
    .B2(_12904_),
    .C1(_12562_),
    .X(_12905_));
 sky130_fd_sc_hd__buf_1 _16945_ (.A(_12543_),
    .X(_12906_));
 sky130_fd_sc_hd__o41a_2 _16946_ (.A1(\decode.regfile.registers_19[4] ),
    .A2(_11013_),
    .A3(_11012_),
    .A4(_12519_),
    .B1(_12906_),
    .X(_12907_));
 sky130_fd_sc_hd__a221o_2 _16947_ (.A1(\decode.regfile.registers_20[4] ),
    .A2(_12771_),
    .B1(_12905_),
    .B2(_12907_),
    .C1(_12538_),
    .X(_12908_));
 sky130_fd_sc_hd__buf_1 _16948_ (.A(_12755_),
    .X(_12909_));
 sky130_fd_sc_hd__o21a_2 _16949_ (.A1(\decode.regfile.registers_21[4] ),
    .A2(_12682_),
    .B1(_12909_),
    .X(_12910_));
 sky130_fd_sc_hd__a221o_2 _16950_ (.A1(\decode.regfile.registers_22[4] ),
    .A2(_12527_),
    .B1(_12908_),
    .B2(_12910_),
    .C1(_12686_),
    .X(_12911_));
 sky130_fd_sc_hd__or4_2 _16951_ (.A(_11015_),
    .B(_10937_),
    .C(\decode.regfile.registers_23[4] ),
    .D(_12520_),
    .X(_12912_));
 sky130_fd_sc_hd__o2111a_2 _16952_ (.A1(_10927_),
    .A2(\decode.regfile.registers_24[4] ),
    .B1(_10933_),
    .C1(_12759_),
    .D1(_12862_),
    .X(_12913_));
 sky130_fd_sc_hd__a31o_2 _16953_ (.A1(_12516_),
    .A2(_12911_),
    .A3(_12912_),
    .B1(_12913_),
    .X(_12914_));
 sky130_fd_sc_hd__buf_1 _16954_ (.A(_10595_),
    .X(_12915_));
 sky130_fd_sc_hd__or4_2 _16955_ (.A(_12915_),
    .B(\decode.regfile.registers_25[4] ),
    .C(_12506_),
    .D(_12812_),
    .X(_12916_));
 sky130_fd_sc_hd__o2111a_2 _16956_ (.A1(_10928_),
    .A2(\decode.regfile.registers_26[4] ),
    .B1(_12814_),
    .C1(_11011_),
    .D1(_11027_),
    .X(_12917_));
 sky130_fd_sc_hd__a31o_2 _16957_ (.A1(_12695_),
    .A2(_12914_),
    .A3(_12916_),
    .B1(_12917_),
    .X(_12918_));
 sky130_fd_sc_hd__or4_2 _16958_ (.A(_10940_),
    .B(_12706_),
    .C(\decode.regfile.registers_27[4] ),
    .D(_12507_),
    .X(_12919_));
 sky130_fd_sc_hd__o21a_2 _16959_ (.A1(_12701_),
    .A2(\decode.regfile.registers_28[4] ),
    .B1(_12698_),
    .X(_12920_));
 sky130_fd_sc_hd__a31o_2 _16960_ (.A1(_12496_),
    .A2(_12918_),
    .A3(_12919_),
    .B1(_12920_),
    .X(_12921_));
 sky130_fd_sc_hd__o221a_2 _16961_ (.A1(_12765_),
    .A2(_12768_),
    .B1(_12493_),
    .B2(\decode.regfile.registers_29[4] ),
    .C1(_12921_),
    .X(_12922_));
 sky130_fd_sc_hd__o221a_2 _16962_ (.A1(_12872_),
    .A2(\decode.regfile.registers_31[4] ),
    .B1(_12873_),
    .B2(_12922_),
    .C1(_12705_),
    .X(_00424_));
 sky130_fd_sc_hd__o21a_2 _16963_ (.A1(_10931_),
    .A2(\decode.regfile.registers_30[5] ),
    .B1(_12487_),
    .X(_12923_));
 sky130_fd_sc_hd__a41o_2 _16964_ (.A1(\decode.regfile.registers_20[5] ),
    .A2(_11024_),
    .A3(_12553_),
    .A4(_12823_),
    .B1(_12824_),
    .X(_12924_));
 sky130_fd_sc_hd__o2111a_2 _16965_ (.A1(\decode.regfile.registers_18[5] ),
    .A2(_10925_),
    .B1(_12569_),
    .C1(_11023_),
    .D1(_11008_),
    .X(_12925_));
 sky130_fd_sc_hd__a41o_2 _16966_ (.A1(\decode.regfile.registers_15[5] ),
    .A2(_12555_),
    .A3(_10923_),
    .A4(_12876_),
    .B1(_12672_),
    .X(_12926_));
 sky130_fd_sc_hd__buf_1 _16967_ (.A(_12533_),
    .X(_12927_));
 sky130_fd_sc_hd__a31o_2 _16968_ (.A1(\decode.regfile.registers_13[5] ),
    .A2(_12927_),
    .A3(_12587_),
    .B1(_12663_),
    .X(_12928_));
 sky130_fd_sc_hd__a22o_2 _16969_ (.A1(\decode.regfile.registers_11[5] ),
    .A2(_12594_),
    .B1(_12582_),
    .B2(_12550_),
    .X(_12929_));
 sky130_fd_sc_hd__a41o_2 _16970_ (.A1(\decode.regfile.registers_9[5] ),
    .A2(_12776_),
    .A3(_12604_),
    .A4(_12532_),
    .B1(_12598_),
    .X(_12930_));
 sky130_fd_sc_hd__or4b_2 _16971_ (.A(_11017_),
    .B(_12539_),
    .C(_12502_),
    .D_N(\decode.regfile.registers_8[5] ),
    .X(_12931_));
 sky130_fd_sc_hd__buf_1 _16972_ (.A(_12630_),
    .X(_12932_));
 sky130_fd_sc_hd__buf_1 _16973_ (.A(_12829_),
    .X(_12933_));
 sky130_fd_sc_hd__buf_1 _16974_ (.A(_12530_),
    .X(_12934_));
 sky130_fd_sc_hd__a31o_2 _16975_ (.A1(_12934_),
    .A2(_12616_),
    .A3(_12557_),
    .B1(\decode.regfile.registers_0[5] ),
    .X(_12935_));
 sky130_fd_sc_hd__o221ai_2 _16976_ (.A1(\decode.regfile.registers_1[5] ),
    .A2(_12932_),
    .B1(_12933_),
    .B2(_10615_),
    .C1(_12935_),
    .Y(_12936_));
 sky130_fd_sc_hd__o21ai_2 _16977_ (.A1(\decode.regfile.registers_2[5] ),
    .A2(_10615_),
    .B1(_12729_),
    .Y(_12937_));
 sky130_fd_sc_hd__o21ai_2 _16978_ (.A1(\decode.regfile.registers_3[5] ),
    .A2(_12628_),
    .B1(_12732_),
    .Y(_12938_));
 sky130_fd_sc_hd__a21oi_2 _16979_ (.A1(_12936_),
    .A2(_12937_),
    .B1(_12938_),
    .Y(_12939_));
 sky130_fd_sc_hd__a221o_2 _16980_ (.A1(\decode.regfile.registers_4[5] ),
    .A2(_12617_),
    .B1(_12619_),
    .B2(\decode.regfile.registers_5[5] ),
    .C1(_12622_),
    .X(_12940_));
 sky130_fd_sc_hd__o32a_2 _16981_ (.A1(\decode.regfile.registers_6[5] ),
    .A2(_10602_),
    .A3(_12614_),
    .B1(_12939_),
    .B2(_12940_),
    .X(_12941_));
 sky130_fd_sc_hd__o32a_2 _16982_ (.A1(_11017_),
    .A2(_12539_),
    .A3(_12502_),
    .B1(\decode.regfile.registers_7[5] ),
    .B2(_12644_),
    .X(_12942_));
 sky130_fd_sc_hd__o21ai_2 _16983_ (.A1(_12611_),
    .A2(_12941_),
    .B1(_12942_),
    .Y(_12943_));
 sky130_fd_sc_hd__a21oi_2 _16984_ (.A1(_12931_),
    .A2(_12943_),
    .B1(_12607_),
    .Y(_12944_));
 sky130_fd_sc_hd__o221a_2 _16985_ (.A1(\decode.regfile.registers_10[5] ),
    .A2(_12653_),
    .B1(_12930_),
    .B2(_12944_),
    .C1(_12792_),
    .X(_12945_));
 sky130_fd_sc_hd__o221a_2 _16986_ (.A1(\decode.regfile.registers_12[5] ),
    .A2(_12745_),
    .B1(_12929_),
    .B2(_12945_),
    .C1(_12658_),
    .X(_12946_));
 sky130_fd_sc_hd__or4_2 _16987_ (.A(\decode.regfile.registers_14[5] ),
    .B(_10603_),
    .C(_10618_),
    .D(_12722_),
    .X(_12947_));
 sky130_fd_sc_hd__o211a_2 _16988_ (.A1(_12928_),
    .A2(_12946_),
    .B1(_12852_),
    .C1(_12947_),
    .X(_12948_));
 sky130_fd_sc_hd__o22a_2 _16989_ (.A1(\decode.regfile.registers_16[5] ),
    .A2(_12575_),
    .B1(_12926_),
    .B2(_12948_),
    .X(_12949_));
 sky130_fd_sc_hd__a31o_2 _16990_ (.A1(_11022_),
    .A2(_12568_),
    .A3(_12535_),
    .B1(_12949_),
    .X(_12950_));
 sky130_fd_sc_hd__o211a_2 _16991_ (.A1(\decode.regfile.registers_17[5] ),
    .A2(_12580_),
    .B1(_12826_),
    .C1(_12950_),
    .X(_12951_));
 sky130_fd_sc_hd__o221a_2 _16992_ (.A1(\decode.regfile.registers_19[5] ),
    .A2(_12679_),
    .B1(_12925_),
    .B2(_12951_),
    .C1(_12545_),
    .X(_12952_));
 sky130_fd_sc_hd__o221a_2 _16993_ (.A1(\decode.regfile.registers_21[5] ),
    .A2(_12822_),
    .B1(_12924_),
    .B2(_12952_),
    .C1(_12806_),
    .X(_12953_));
 sky130_fd_sc_hd__a211o_2 _16994_ (.A1(\decode.regfile.registers_22[5] ),
    .A2(_12528_),
    .B1(_12953_),
    .C1(_12687_),
    .X(_12954_));
 sky130_fd_sc_hd__or4_2 _16995_ (.A(_11015_),
    .B(_10937_),
    .C(\decode.regfile.registers_23[5] ),
    .D(_12520_),
    .X(_12955_));
 sky130_fd_sc_hd__o2111a_2 _16996_ (.A1(_10927_),
    .A2(\decode.regfile.registers_24[5] ),
    .B1(_10933_),
    .C1(_12759_),
    .D1(_12862_),
    .X(_12956_));
 sky130_fd_sc_hd__a31o_2 _16997_ (.A1(_12516_),
    .A2(_12954_),
    .A3(_12955_),
    .B1(_12956_),
    .X(_12957_));
 sky130_fd_sc_hd__or4_2 _16998_ (.A(_12915_),
    .B(\decode.regfile.registers_25[5] ),
    .C(_12506_),
    .D(_12812_),
    .X(_12958_));
 sky130_fd_sc_hd__o2111a_2 _16999_ (.A1(_10928_),
    .A2(\decode.regfile.registers_26[5] ),
    .B1(_12814_),
    .C1(_11011_),
    .D1(_11027_),
    .X(_12959_));
 sky130_fd_sc_hd__a31o_2 _17000_ (.A1(_12695_),
    .A2(_12957_),
    .A3(_12958_),
    .B1(_12959_),
    .X(_12960_));
 sky130_fd_sc_hd__or4_2 _17001_ (.A(_10940_),
    .B(_12706_),
    .C(\decode.regfile.registers_27[5] ),
    .D(_12507_),
    .X(_12961_));
 sky130_fd_sc_hd__o21a_2 _17002_ (.A1(_12701_),
    .A2(\decode.regfile.registers_28[5] ),
    .B1(_12698_),
    .X(_12962_));
 sky130_fd_sc_hd__a31o_2 _17003_ (.A1(_12496_),
    .A2(_12960_),
    .A3(_12961_),
    .B1(_12962_),
    .X(_12963_));
 sky130_fd_sc_hd__o221a_2 _17004_ (.A1(_12765_),
    .A2(_12768_),
    .B1(_12493_),
    .B2(\decode.regfile.registers_29[5] ),
    .C1(_12963_),
    .X(_12964_));
 sky130_fd_sc_hd__o221a_2 _17005_ (.A1(_12708_),
    .A2(\decode.regfile.registers_31[5] ),
    .B1(_12923_),
    .B2(_12964_),
    .C1(_12705_),
    .X(_00425_));
 sky130_fd_sc_hd__buf_1 _17006_ (.A(_12492_),
    .X(_12965_));
 sky130_fd_sc_hd__o21a_2 _17007_ (.A1(_10930_),
    .A2(\decode.regfile.registers_28[6] ),
    .B1(_12698_),
    .X(_12966_));
 sky130_fd_sc_hd__buf_1 _17008_ (.A(_12495_),
    .X(_12967_));
 sky130_fd_sc_hd__buf_1 _17009_ (.A(_12694_),
    .X(_12968_));
 sky130_fd_sc_hd__a221oi_2 _17010_ (.A1(\decode.regfile.registers_2[6] ),
    .A2(_12835_),
    .B1(_12836_),
    .B2(\decode.regfile.registers_3[6] ),
    .C1(_12838_),
    .Y(_12969_));
 sky130_fd_sc_hd__a31o_2 _17011_ (.A1(_12532_),
    .A2(_10593_),
    .A3(_12559_),
    .B1(\decode.regfile.registers_0[6] ),
    .X(_12970_));
 sky130_fd_sc_hd__o211ai_2 _17012_ (.A1(\decode.regfile.registers_1[6] ),
    .A2(_12778_),
    .B1(_12830_),
    .C1(_12970_),
    .Y(_12971_));
 sky130_fd_sc_hd__a221oi_2 _17013_ (.A1(\decode.regfile.registers_4[6] ),
    .A2(_12549_),
    .B1(_12532_),
    .B2(\decode.regfile.registers_5[6] ),
    .C1(_12615_),
    .Y(_12972_));
 sky130_fd_sc_hd__a21oi_2 _17014_ (.A1(_12969_),
    .A2(_12971_),
    .B1(_12972_),
    .Y(_12973_));
 sky130_fd_sc_hd__a221oi_2 _17015_ (.A1(\decode.regfile.registers_7[6] ),
    .A2(_12612_),
    .B1(_12623_),
    .B2(\decode.regfile.registers_6[6] ),
    .C1(_12973_),
    .Y(_12974_));
 sky130_fd_sc_hd__a21oi_2 _17016_ (.A1(\decode.regfile.registers_8[6] ),
    .A2(_12889_),
    .B1(_12607_),
    .Y(_12975_));
 sky130_fd_sc_hd__o21ai_2 _17017_ (.A1(_12889_),
    .A2(_12974_),
    .B1(_12975_),
    .Y(_12976_));
 sky130_fd_sc_hd__buf_1 _17018_ (.A(_12502_),
    .X(_12977_));
 sky130_fd_sc_hd__o41a_2 _17019_ (.A1(\decode.regfile.registers_9[6] ),
    .A2(_11018_),
    .A3(_12977_),
    .A4(_12510_),
    .B1(_12653_),
    .X(_12978_));
 sky130_fd_sc_hd__a221o_2 _17020_ (.A1(\decode.regfile.registers_10[6] ),
    .A2(_12600_),
    .B1(_12976_),
    .B2(_12978_),
    .C1(_12724_),
    .X(_12979_));
 sky130_fd_sc_hd__o32a_2 _17021_ (.A1(_12499_),
    .A2(_12541_),
    .A3(_12490_),
    .B1(\decode.regfile.registers_11[6] ),
    .B2(_12878_),
    .X(_12980_));
 sky130_fd_sc_hd__a32o_2 _17022_ (.A1(\decode.regfile.registers_12[6] ),
    .A2(_12551_),
    .A3(_12588_),
    .B1(_12979_),
    .B2(_12980_),
    .X(_12981_));
 sky130_fd_sc_hd__and3_2 _17023_ (.A(\decode.regfile.registers_13[6] ),
    .B(_12927_),
    .C(_12588_),
    .X(_12982_));
 sky130_fd_sc_hd__a211o_2 _17024_ (.A1(_12659_),
    .A2(_12981_),
    .B1(_12982_),
    .C1(_12664_),
    .X(_12983_));
 sky130_fd_sc_hd__buf_1 _17025_ (.A(_12669_),
    .X(_12984_));
 sky130_fd_sc_hd__o32a_2 _17026_ (.A1(_11020_),
    .A2(_12491_),
    .A3(_12666_),
    .B1(\decode.regfile.registers_14[6] ),
    .B2(_12984_),
    .X(_12985_));
 sky130_fd_sc_hd__a22oi_2 _17027_ (.A1(\decode.regfile.registers_15[6] ),
    .A2(_12585_),
    .B1(_12983_),
    .B2(_12985_),
    .Y(_12986_));
 sky130_fd_sc_hd__a21oi_2 _17028_ (.A1(\decode.regfile.registers_16[6] ),
    .A2(_12673_),
    .B1(_12901_),
    .Y(_12987_));
 sky130_fd_sc_hd__o21ai_2 _17029_ (.A1(_12674_),
    .A2(_12986_),
    .B1(_12987_),
    .Y(_12988_));
 sky130_fd_sc_hd__o211a_2 _17030_ (.A1(\decode.regfile.registers_17[6] ),
    .A2(_12580_),
    .B1(_12826_),
    .C1(_12988_),
    .X(_12989_));
 sky130_fd_sc_hd__a211o_2 _17031_ (.A1(\decode.regfile.registers_18[6] ),
    .A2(_12572_),
    .B1(_12561_),
    .C1(_12989_),
    .X(_12990_));
 sky130_fd_sc_hd__o41a_2 _17032_ (.A1(\decode.regfile.registers_19[6] ),
    .A2(_10599_),
    .A3(_10589_),
    .A4(_12518_),
    .B1(_12544_),
    .X(_12991_));
 sky130_fd_sc_hd__a221o_2 _17033_ (.A1(\decode.regfile.registers_20[6] ),
    .A2(_12771_),
    .B1(_12990_),
    .B2(_12991_),
    .C1(_12538_),
    .X(_12992_));
 sky130_fd_sc_hd__o21a_2 _17034_ (.A1(\decode.regfile.registers_21[6] ),
    .A2(_12822_),
    .B1(_12909_),
    .X(_12993_));
 sky130_fd_sc_hd__a221o_2 _17035_ (.A1(\decode.regfile.registers_22[6] ),
    .A2(_12527_),
    .B1(_12992_),
    .B2(_12993_),
    .C1(_12686_),
    .X(_12994_));
 sky130_fd_sc_hd__buf_1 _17036_ (.A(_12519_),
    .X(_12995_));
 sky130_fd_sc_hd__or4_2 _17037_ (.A(_11014_),
    .B(_10936_),
    .C(\decode.regfile.registers_23[6] ),
    .D(_12995_),
    .X(_12996_));
 sky130_fd_sc_hd__buf_1 _17038_ (.A(_10604_),
    .X(_12997_));
 sky130_fd_sc_hd__buf_1 _17039_ (.A(_12690_),
    .X(_12998_));
 sky130_fd_sc_hd__o2111a_2 _17040_ (.A1(_12712_),
    .A2(\decode.regfile.registers_24[6] ),
    .B1(_12997_),
    .C1(_12998_),
    .D1(_11025_),
    .X(_12999_));
 sky130_fd_sc_hd__a31o_2 _17041_ (.A1(_12515_),
    .A2(_12994_),
    .A3(_12996_),
    .B1(_12999_),
    .X(_13000_));
 sky130_fd_sc_hd__or4_2 _17042_ (.A(_10938_),
    .B(\decode.regfile.registers_25[6] ),
    .C(_12505_),
    .D(_12811_),
    .X(_13001_));
 sky130_fd_sc_hd__buf_1 _17043_ (.A(_12759_),
    .X(_13002_));
 sky130_fd_sc_hd__o2111a_2 _17044_ (.A1(_12494_),
    .A2(\decode.regfile.registers_26[6] ),
    .B1(_13002_),
    .C1(_11010_),
    .D1(_11026_),
    .X(_13003_));
 sky130_fd_sc_hd__a31o_2 _17045_ (.A1(_12968_),
    .A2(_13000_),
    .A3(_13001_),
    .B1(_13003_),
    .X(_13004_));
 sky130_fd_sc_hd__o311a_2 _17046_ (.A1(\decode.regfile.registers_27[6] ),
    .A2(_12507_),
    .A3(_12520_),
    .B1(_12967_),
    .C1(_13004_),
    .X(_13005_));
 sky130_fd_sc_hd__o221a_2 _17047_ (.A1(\decode.regfile.registers_29[6] ),
    .A2(_12965_),
    .B1(_12966_),
    .B2(_13005_),
    .C1(_12702_),
    .X(_13006_));
 sky130_fd_sc_hd__o21a_2 _17048_ (.A1(_10931_),
    .A2(\decode.regfile.registers_30[6] ),
    .B1(_12487_),
    .X(_13007_));
 sky130_fd_sc_hd__or4_2 _17049_ (.A(\decode.regfile.registers_31[6] ),
    .B(_12491_),
    .C(_12706_),
    .D(_10940_),
    .X(_13008_));
 sky130_fd_sc_hd__o211a_2 _17050_ (.A1(_13006_),
    .A2(_13007_),
    .B1(_12704_),
    .C1(_13008_),
    .X(_00426_));
 sky130_fd_sc_hd__o21a_2 _17051_ (.A1(_10931_),
    .A2(\decode.regfile.registers_30[7] ),
    .B1(_12487_),
    .X(_13009_));
 sky130_fd_sc_hd__a32o_2 _17052_ (.A1(_11023_),
    .A2(_12552_),
    .A3(_12523_),
    .B1(_12561_),
    .B2(\decode.regfile.registers_19[7] ),
    .X(_13010_));
 sky130_fd_sc_hd__buf_1 _17053_ (.A(_12575_),
    .X(_13011_));
 sky130_fd_sc_hd__a2bb2o_2 _17054_ (.A1_N(\decode.regfile.registers_12[7] ),
    .A2_N(_12745_),
    .B1(_12587_),
    .B2(_12533_),
    .X(_13012_));
 sky130_fd_sc_hd__a31o_2 _17055_ (.A1(\decode.regfile.registers_2[7] ),
    .A2(_10608_),
    .A3(_12635_),
    .B1(_12638_),
    .X(_13013_));
 sky130_fd_sc_hd__a31o_2 _17056_ (.A1(_12530_),
    .A2(_12616_),
    .A3(_12557_),
    .B1(\decode.regfile.registers_0[7] ),
    .X(_13014_));
 sky130_fd_sc_hd__o221a_2 _17057_ (.A1(\decode.regfile.registers_1[7] ),
    .A2(_12631_),
    .B1(_12933_),
    .B2(_12508_),
    .C1(_13014_),
    .X(_13015_));
 sky130_fd_sc_hd__o22a_2 _17058_ (.A1(\decode.regfile.registers_3[7] ),
    .A2(_12628_),
    .B1(_13013_),
    .B2(_13015_),
    .X(_13016_));
 sky130_fd_sc_hd__a221o_2 _17059_ (.A1(\decode.regfile.registers_4[7] ),
    .A2(_12617_),
    .B1(_12619_),
    .B2(\decode.regfile.registers_5[7] ),
    .C1(_12622_),
    .X(_13017_));
 sky130_fd_sc_hd__a21o_2 _17060_ (.A1(_13016_),
    .A2(_12732_),
    .B1(_13017_),
    .X(_13018_));
 sky130_fd_sc_hd__o31a_2 _17061_ (.A1(\decode.regfile.registers_6[7] ),
    .A2(_10602_),
    .A3(_12626_),
    .B1(_12645_),
    .X(_13019_));
 sky130_fd_sc_hd__and3_2 _17062_ (.A(_12522_),
    .B(_12616_),
    .C(_10608_),
    .X(_13020_));
 sky130_fd_sc_hd__and3_2 _17063_ (.A(\decode.regfile.registers_7[7] ),
    .B(_10616_),
    .C(_13020_),
    .X(_13021_));
 sky130_fd_sc_hd__a211o_2 _17064_ (.A1(_13018_),
    .A2(_13019_),
    .B1(_13021_),
    .C1(_12889_),
    .X(_13022_));
 sky130_fd_sc_hd__o211ai_2 _17065_ (.A1(\decode.regfile.registers_8[7] ),
    .A2(_12892_),
    .B1(_12603_),
    .C1(_13022_),
    .Y(_13023_));
 sky130_fd_sc_hd__a21oi_2 _17066_ (.A1(\decode.regfile.registers_9[7] ),
    .A2(_12607_),
    .B1(_12599_),
    .Y(_13024_));
 sky130_fd_sc_hd__o21ai_2 _17067_ (.A1(\decode.regfile.registers_10[7] ),
    .A2(_12790_),
    .B1(_12792_),
    .Y(_13025_));
 sky130_fd_sc_hd__a21oi_2 _17068_ (.A1(_13023_),
    .A2(_13024_),
    .B1(_13025_),
    .Y(_13026_));
 sky130_fd_sc_hd__a221oi_2 _17069_ (.A1(\decode.regfile.registers_11[7] ),
    .A2(_12595_),
    .B1(_12587_),
    .B2(_12551_),
    .C1(_13026_),
    .Y(_13027_));
 sky130_fd_sc_hd__a21oi_2 _17070_ (.A1(\decode.regfile.registers_13[7] ),
    .A2(_12775_),
    .B1(_12663_),
    .Y(_13028_));
 sky130_fd_sc_hd__o21ai_2 _17071_ (.A1(_13012_),
    .A2(_13027_),
    .B1(_13028_),
    .Y(_13029_));
 sky130_fd_sc_hd__o221ai_2 _17072_ (.A1(_12666_),
    .A2(_12723_),
    .B1(_12984_),
    .B2(\decode.regfile.registers_14[7] ),
    .C1(_13029_),
    .Y(_13030_));
 sky130_fd_sc_hd__buf_1 _17073_ (.A(_12672_),
    .X(_13031_));
 sky130_fd_sc_hd__a21oi_2 _17074_ (.A1(\decode.regfile.registers_15[7] ),
    .A2(_12584_),
    .B1(_13031_),
    .Y(_13032_));
 sky130_fd_sc_hd__nand2_2 _17075_ (.A(_13030_),
    .B(_13032_),
    .Y(_13033_));
 sky130_fd_sc_hd__o211a_2 _17076_ (.A1(\decode.regfile.registers_16[7] ),
    .A2(_13011_),
    .B1(_12578_),
    .C1(_13033_),
    .X(_13034_));
 sky130_fd_sc_hd__a211o_2 _17077_ (.A1(\decode.regfile.registers_17[7] ),
    .A2(_12901_),
    .B1(_12571_),
    .C1(_13034_),
    .X(_13035_));
 sky130_fd_sc_hd__o211a_2 _17078_ (.A1(\decode.regfile.registers_18[7] ),
    .A2(_12566_),
    .B1(_12678_),
    .C1(_13035_),
    .X(_13036_));
 sky130_fd_sc_hd__o22a_2 _17079_ (.A1(\decode.regfile.registers_20[7] ),
    .A2(_12545_),
    .B1(_13010_),
    .B2(_13036_),
    .X(_13037_));
 sky130_fd_sc_hd__a31o_2 _17080_ (.A1(_12546_),
    .A2(_12554_),
    .A3(_12535_),
    .B1(_13037_),
    .X(_13038_));
 sky130_fd_sc_hd__o21a_2 _17081_ (.A1(\decode.regfile.registers_21[7] ),
    .A2(_12682_),
    .B1(_12909_),
    .X(_13039_));
 sky130_fd_sc_hd__a221o_2 _17082_ (.A1(\decode.regfile.registers_22[7] ),
    .A2(_12527_),
    .B1(_13038_),
    .B2(_13039_),
    .C1(_12686_),
    .X(_13040_));
 sky130_fd_sc_hd__buf_1 _17083_ (.A(_12519_),
    .X(_13041_));
 sky130_fd_sc_hd__or4_2 _17084_ (.A(_11015_),
    .B(_10937_),
    .C(\decode.regfile.registers_23[7] ),
    .D(_13041_),
    .X(_13042_));
 sky130_fd_sc_hd__o2111a_2 _17085_ (.A1(_10927_),
    .A2(\decode.regfile.registers_24[7] ),
    .B1(_10933_),
    .C1(_12759_),
    .D1(_12862_),
    .X(_13043_));
 sky130_fd_sc_hd__a31o_2 _17086_ (.A1(_12516_),
    .A2(_13040_),
    .A3(_13042_),
    .B1(_13043_),
    .X(_13044_));
 sky130_fd_sc_hd__buf_1 _17087_ (.A(_12505_),
    .X(_13045_));
 sky130_fd_sc_hd__or4_2 _17088_ (.A(_12915_),
    .B(\decode.regfile.registers_25[7] ),
    .C(_13045_),
    .D(_12812_),
    .X(_13046_));
 sky130_fd_sc_hd__buf_1 _17089_ (.A(_11010_),
    .X(_13047_));
 sky130_fd_sc_hd__o2111a_2 _17090_ (.A1(_10928_),
    .A2(\decode.regfile.registers_26[7] ),
    .B1(_12814_),
    .C1(_13047_),
    .D1(_11027_),
    .X(_13048_));
 sky130_fd_sc_hd__a31o_2 _17091_ (.A1(_12695_),
    .A2(_13044_),
    .A3(_13046_),
    .B1(_13048_),
    .X(_13049_));
 sky130_fd_sc_hd__buf_1 _17092_ (.A(_12506_),
    .X(_13050_));
 sky130_fd_sc_hd__or4_2 _17093_ (.A(_10940_),
    .B(_12706_),
    .C(\decode.regfile.registers_27[7] ),
    .D(_13050_),
    .X(_13051_));
 sky130_fd_sc_hd__o21a_2 _17094_ (.A1(_12701_),
    .A2(\decode.regfile.registers_28[7] ),
    .B1(_12698_),
    .X(_13052_));
 sky130_fd_sc_hd__a31o_2 _17095_ (.A1(_12496_),
    .A2(_13049_),
    .A3(_13051_),
    .B1(_13052_),
    .X(_13053_));
 sky130_fd_sc_hd__o221a_2 _17096_ (.A1(_12765_),
    .A2(_12768_),
    .B1(_12493_),
    .B2(\decode.regfile.registers_29[7] ),
    .C1(_13053_),
    .X(_13054_));
 sky130_fd_sc_hd__o221a_2 _17097_ (.A1(\decode.regfile.registers_31[7] ),
    .A2(_12709_),
    .B1(_13009_),
    .B2(_13054_),
    .C1(_12705_),
    .X(_00427_));
 sky130_fd_sc_hd__buf_1 _17098_ (.A(_10930_),
    .X(_13055_));
 sky130_fd_sc_hd__o21a_2 _17099_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[8] ),
    .B1(_12487_),
    .X(_13056_));
 sky130_fd_sc_hd__a221o_2 _17100_ (.A1(\decode.regfile.registers_7[8] ),
    .A2(_12610_),
    .B1(_12737_),
    .B2(\decode.regfile.registers_6[8] ),
    .C1(_12843_),
    .X(_13057_));
 sky130_fd_sc_hd__and3_2 _17101_ (.A(\decode.regfile.registers_1[8] ),
    .B(_12636_),
    .C(_12531_),
    .X(_13058_));
 sky130_fd_sc_hd__a2bb2o_2 _17102_ (.A1_N(_12882_),
    .A2_N(_12933_),
    .B1(_12932_),
    .B2(\decode.regfile.registers_0[8] ),
    .X(_13059_));
 sky130_fd_sc_hd__o221ai_2 _17103_ (.A1(\decode.regfile.registers_2[8] ),
    .A2(_12634_),
    .B1(_13058_),
    .B2(_13059_),
    .C1(_12629_),
    .Y(_13060_));
 sky130_fd_sc_hd__o2bb2a_2 _17104_ (.A1_N(\decode.regfile.registers_3[8] ),
    .A2_N(_12836_),
    .B1(_10609_),
    .B2(_12614_),
    .X(_13061_));
 sky130_fd_sc_hd__a221oi_2 _17105_ (.A1(\decode.regfile.registers_4[8] ),
    .A2(_12549_),
    .B1(_12532_),
    .B2(\decode.regfile.registers_5[8] ),
    .C1(_12626_),
    .Y(_13062_));
 sky130_fd_sc_hd__a21oi_2 _17106_ (.A1(_13060_),
    .A2(_13061_),
    .B1(_13062_),
    .Y(_13063_));
 sky130_fd_sc_hd__o221a_2 _17107_ (.A1(\decode.regfile.registers_8[8] ),
    .A2(_12726_),
    .B1(_13057_),
    .B2(_13063_),
    .C1(_12602_),
    .X(_13064_));
 sky130_fd_sc_hd__a41o_2 _17108_ (.A1(\decode.regfile.registers_9[8] ),
    .A2(_10594_),
    .A3(_12690_),
    .A4(_12533_),
    .B1(_13064_),
    .X(_13065_));
 sky130_fd_sc_hd__o2111a_2 _17109_ (.A1(\decode.regfile.registers_10[8] ),
    .A2(_10617_),
    .B1(_10594_),
    .C1(_10611_),
    .D1(_12690_),
    .X(_13066_));
 sky130_fd_sc_hd__a21o_2 _17110_ (.A1(_12654_),
    .A2(_13065_),
    .B1(_13066_),
    .X(_13067_));
 sky130_fd_sc_hd__o32a_2 _17111_ (.A1(_12499_),
    .A2(_12541_),
    .A3(_12490_),
    .B1(\decode.regfile.registers_11[8] ),
    .B2(_12878_),
    .X(_13068_));
 sky130_fd_sc_hd__a221o_2 _17112_ (.A1(\decode.regfile.registers_12[8] ),
    .A2(_12794_),
    .B1(_13067_),
    .B2(_13068_),
    .C1(_12775_),
    .X(_13069_));
 sky130_fd_sc_hd__o31a_2 _17113_ (.A1(\decode.regfile.registers_13[8] ),
    .A2(_12512_),
    .A3(_12723_),
    .B1(_12984_),
    .X(_13070_));
 sky130_fd_sc_hd__a221o_2 _17114_ (.A1(\decode.regfile.registers_14[8] ),
    .A2(_12664_),
    .B1(_13069_),
    .B2(_13070_),
    .C1(_12585_),
    .X(_13071_));
 sky130_fd_sc_hd__o31a_2 _17115_ (.A1(\decode.regfile.registers_15[8] ),
    .A2(_12667_),
    .A3(_12773_),
    .B1(_13011_),
    .X(_13072_));
 sky130_fd_sc_hd__a32o_2 _17116_ (.A1(_11021_),
    .A2(_12567_),
    .A3(_12586_),
    .B1(_12673_),
    .B2(\decode.regfile.registers_16[8] ),
    .X(_13073_));
 sky130_fd_sc_hd__a21o_2 _17117_ (.A1(_13071_),
    .A2(_13072_),
    .B1(_13073_),
    .X(_13074_));
 sky130_fd_sc_hd__o211a_2 _17118_ (.A1(\decode.regfile.registers_17[8] ),
    .A2(_12580_),
    .B1(_12826_),
    .C1(_13074_),
    .X(_13075_));
 sky130_fd_sc_hd__a211o_2 _17119_ (.A1(\decode.regfile.registers_18[8] ),
    .A2(_12572_),
    .B1(_12562_),
    .C1(_13075_),
    .X(_13076_));
 sky130_fd_sc_hd__o41a_2 _17120_ (.A1(\decode.regfile.registers_19[8] ),
    .A2(_11013_),
    .A3(_10589_),
    .A4(_12519_),
    .B1(_12544_),
    .X(_13077_));
 sky130_fd_sc_hd__a221o_2 _17121_ (.A1(\decode.regfile.registers_20[8] ),
    .A2(_12771_),
    .B1(_13076_),
    .B2(_13077_),
    .C1(_12538_),
    .X(_13078_));
 sky130_fd_sc_hd__o21a_2 _17122_ (.A1(\decode.regfile.registers_21[8] ),
    .A2(_12682_),
    .B1(_12909_),
    .X(_13079_));
 sky130_fd_sc_hd__a221o_2 _17123_ (.A1(\decode.regfile.registers_22[8] ),
    .A2(_12527_),
    .B1(_13078_),
    .B2(_13079_),
    .C1(_12686_),
    .X(_13080_));
 sky130_fd_sc_hd__buf_1 _17124_ (.A(_11013_),
    .X(_13081_));
 sky130_fd_sc_hd__or4_2 _17125_ (.A(_13081_),
    .B(_10937_),
    .C(\decode.regfile.registers_23[8] ),
    .D(_13041_),
    .X(_13082_));
 sky130_fd_sc_hd__buf_1 _17126_ (.A(_12690_),
    .X(_13083_));
 sky130_fd_sc_hd__o2111a_2 _17127_ (.A1(_10927_),
    .A2(\decode.regfile.registers_24[8] ),
    .B1(_10933_),
    .C1(_13083_),
    .D1(_12862_),
    .X(_13084_));
 sky130_fd_sc_hd__a31o_2 _17128_ (.A1(_12516_),
    .A2(_13080_),
    .A3(_13082_),
    .B1(_13084_),
    .X(_13085_));
 sky130_fd_sc_hd__or4_2 _17129_ (.A(_12915_),
    .B(\decode.regfile.registers_25[8] ),
    .C(_13045_),
    .D(_12812_),
    .X(_13086_));
 sky130_fd_sc_hd__buf_1 _17130_ (.A(_12494_),
    .X(_13087_));
 sky130_fd_sc_hd__buf_1 _17131_ (.A(_11026_),
    .X(_13088_));
 sky130_fd_sc_hd__o2111a_2 _17132_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[8] ),
    .B1(_12814_),
    .C1(_13047_),
    .D1(_13088_),
    .X(_13089_));
 sky130_fd_sc_hd__a31o_2 _17133_ (.A1(_12695_),
    .A2(_13085_),
    .A3(_13086_),
    .B1(_13089_),
    .X(_13090_));
 sky130_fd_sc_hd__buf_1 _17134_ (.A(_10939_),
    .X(_13091_));
 sky130_fd_sc_hd__or4_2 _17135_ (.A(_13091_),
    .B(_12706_),
    .C(\decode.regfile.registers_27[8] ),
    .D(_13050_),
    .X(_13092_));
 sky130_fd_sc_hd__buf_1 _17136_ (.A(_12697_),
    .X(_13093_));
 sky130_fd_sc_hd__o21a_2 _17137_ (.A1(_12701_),
    .A2(\decode.regfile.registers_28[8] ),
    .B1(_13093_),
    .X(_13094_));
 sky130_fd_sc_hd__a31o_2 _17138_ (.A1(_12496_),
    .A2(_13090_),
    .A3(_13092_),
    .B1(_13094_),
    .X(_13095_));
 sky130_fd_sc_hd__o221a_2 _17139_ (.A1(_12765_),
    .A2(_12768_),
    .B1(_12493_),
    .B2(\decode.regfile.registers_29[8] ),
    .C1(_13095_),
    .X(_13096_));
 sky130_fd_sc_hd__o221a_2 _17140_ (.A1(_12708_),
    .A2(\decode.regfile.registers_31[8] ),
    .B1(_13056_),
    .B2(_13096_),
    .C1(_12705_),
    .X(_00428_));
 sky130_fd_sc_hd__buf_1 _17141_ (.A(_12486_),
    .X(_13097_));
 sky130_fd_sc_hd__o21a_2 _17142_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[9] ),
    .B1(_13097_),
    .X(_13098_));
 sky130_fd_sc_hd__buf_1 _17143_ (.A(_10930_),
    .X(_13099_));
 sky130_fd_sc_hd__buf_1 _17144_ (.A(_12527_),
    .X(_13100_));
 sky130_fd_sc_hd__a41o_2 _17145_ (.A1(\decode.regfile.registers_15[9] ),
    .A2(_10612_),
    .A3(_10924_),
    .A4(_12589_),
    .B1(_12673_),
    .X(_13101_));
 sky130_fd_sc_hd__a31o_2 _17146_ (.A1(\decode.regfile.registers_2[9] ),
    .A2(_10608_),
    .A3(_12636_),
    .B1(_12639_),
    .X(_13102_));
 sky130_fd_sc_hd__a31o_2 _17147_ (.A1(_12934_),
    .A2(_12616_),
    .A3(_12557_),
    .B1(\decode.regfile.registers_0[9] ),
    .X(_13103_));
 sky130_fd_sc_hd__o221a_2 _17148_ (.A1(\decode.regfile.registers_1[9] ),
    .A2(_12932_),
    .B1(_12933_),
    .B2(_10615_),
    .C1(_13103_),
    .X(_13104_));
 sky130_fd_sc_hd__o22a_2 _17149_ (.A1(\decode.regfile.registers_3[9] ),
    .A2(_12628_),
    .B1(_13102_),
    .B2(_13104_),
    .X(_13105_));
 sky130_fd_sc_hd__a221o_2 _17150_ (.A1(\decode.regfile.registers_4[9] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[9] ),
    .C1(_12622_),
    .X(_13106_));
 sky130_fd_sc_hd__a21o_2 _17151_ (.A1(_13105_),
    .A2(_12732_),
    .B1(_13106_),
    .X(_13107_));
 sky130_fd_sc_hd__o31a_2 _17152_ (.A1(\decode.regfile.registers_6[9] ),
    .A2(_10602_),
    .A3(_12626_),
    .B1(_12645_),
    .X(_13108_));
 sky130_fd_sc_hd__a31o_2 _17153_ (.A1(\decode.regfile.registers_7[9] ),
    .A2(_10617_),
    .A3(_13020_),
    .B1(_12888_),
    .X(_13109_));
 sky130_fd_sc_hd__a21o_2 _17154_ (.A1(_13107_),
    .A2(_13108_),
    .B1(_13109_),
    .X(_13110_));
 sky130_fd_sc_hd__o211ai_2 _17155_ (.A1(\decode.regfile.registers_8[9] ),
    .A2(_12892_),
    .B1(_12603_),
    .C1(_13110_),
    .Y(_13111_));
 sky130_fd_sc_hd__or4b_2 _17156_ (.A(_11018_),
    .B(_12977_),
    .C(_12510_),
    .D_N(\decode.regfile.registers_9[9] ),
    .X(_13112_));
 sky130_fd_sc_hd__o21ai_2 _17157_ (.A1(\decode.regfile.registers_10[9] ),
    .A2(_12790_),
    .B1(_12792_),
    .Y(_13113_));
 sky130_fd_sc_hd__a31o_2 _17158_ (.A1(_12654_),
    .A2(_13111_),
    .A3(_13112_),
    .B1(_13113_),
    .X(_13114_));
 sky130_fd_sc_hd__o2bb2a_2 _17159_ (.A1_N(\decode.regfile.registers_11[9] ),
    .A2_N(_12724_),
    .B1(_12722_),
    .B2(_12540_),
    .X(_13115_));
 sky130_fd_sc_hd__nand2_2 _17160_ (.A(_13114_),
    .B(_13115_),
    .Y(_13116_));
 sky130_fd_sc_hd__o32a_2 _17161_ (.A1(_12499_),
    .A2(_12490_),
    .A3(_12511_),
    .B1(\decode.regfile.registers_12[9] ),
    .B2(_12745_),
    .X(_13117_));
 sky130_fd_sc_hd__a221o_2 _17162_ (.A1(\decode.regfile.registers_13[9] ),
    .A2(_12775_),
    .B1(_13116_),
    .B2(_13117_),
    .C1(_12664_),
    .X(_13118_));
 sky130_fd_sc_hd__o221a_2 _17163_ (.A1(_12667_),
    .A2(_12773_),
    .B1(_12670_),
    .B2(\decode.regfile.registers_14[9] ),
    .C1(_13118_),
    .X(_13119_));
 sky130_fd_sc_hd__o22a_2 _17164_ (.A1(\decode.regfile.registers_16[9] ),
    .A2(_12576_),
    .B1(_13101_),
    .B2(_13119_),
    .X(_13120_));
 sky130_fd_sc_hd__a31o_2 _17165_ (.A1(_11023_),
    .A2(_12569_),
    .A3(_12535_),
    .B1(_13120_),
    .X(_13121_));
 sky130_fd_sc_hd__o21a_2 _17166_ (.A1(\decode.regfile.registers_17[9] ),
    .A2(_12580_),
    .B1(_12826_),
    .X(_13122_));
 sky130_fd_sc_hd__a221o_2 _17167_ (.A1(\decode.regfile.registers_18[9] ),
    .A2(_12572_),
    .B1(_13121_),
    .B2(_13122_),
    .C1(_12562_),
    .X(_13123_));
 sky130_fd_sc_hd__o41a_2 _17168_ (.A1(\decode.regfile.registers_19[9] ),
    .A2(_11013_),
    .A3(_11012_),
    .A4(_12519_),
    .B1(_12545_),
    .X(_13124_));
 sky130_fd_sc_hd__a221o_2 _17169_ (.A1(\decode.regfile.registers_20[9] ),
    .A2(_12771_),
    .B1(_13123_),
    .B2(_13124_),
    .C1(_12538_),
    .X(_13125_));
 sky130_fd_sc_hd__o21a_2 _17170_ (.A1(\decode.regfile.registers_21[9] ),
    .A2(_12682_),
    .B1(_12806_),
    .X(_13126_));
 sky130_fd_sc_hd__a221o_2 _17171_ (.A1(\decode.regfile.registers_22[9] ),
    .A2(_13100_),
    .B1(_13125_),
    .B2(_13126_),
    .C1(_12687_),
    .X(_13127_));
 sky130_fd_sc_hd__o32a_2 _17172_ (.A1(_10938_),
    .A2(_12542_),
    .A3(_12505_),
    .B1(\decode.regfile.registers_23[9] ),
    .B2(_12714_),
    .X(_13128_));
 sky130_fd_sc_hd__o2111a_2 _17173_ (.A1(_10927_),
    .A2(\decode.regfile.registers_24[9] ),
    .B1(_10933_),
    .C1(_12759_),
    .D1(_11026_),
    .X(_13129_));
 sky130_fd_sc_hd__a21o_2 _17174_ (.A1(_13127_),
    .A2(_13128_),
    .B1(_13129_),
    .X(_13130_));
 sky130_fd_sc_hd__or4_2 _17175_ (.A(_12915_),
    .B(\decode.regfile.registers_25[9] ),
    .C(_13045_),
    .D(_12812_),
    .X(_13131_));
 sky130_fd_sc_hd__o2111a_2 _17176_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[9] ),
    .B1(_12814_),
    .C1(_13047_),
    .D1(_13088_),
    .X(_13132_));
 sky130_fd_sc_hd__a31o_2 _17177_ (.A1(_12695_),
    .A2(_13130_),
    .A3(_13131_),
    .B1(_13132_),
    .X(_13133_));
 sky130_fd_sc_hd__or4_2 _17178_ (.A(_13091_),
    .B(_12706_),
    .C(\decode.regfile.registers_27[9] ),
    .D(_13050_),
    .X(_13134_));
 sky130_fd_sc_hd__o21a_2 _17179_ (.A1(_12701_),
    .A2(\decode.regfile.registers_28[9] ),
    .B1(_13093_),
    .X(_13135_));
 sky130_fd_sc_hd__a31o_2 _17180_ (.A1(_12496_),
    .A2(_13133_),
    .A3(_13134_),
    .B1(_13135_),
    .X(_13136_));
 sky130_fd_sc_hd__o221a_2 _17181_ (.A1(_13099_),
    .A2(_12768_),
    .B1(_12493_),
    .B2(\decode.regfile.registers_29[9] ),
    .C1(_13136_),
    .X(_13137_));
 sky130_fd_sc_hd__o221a_2 _17182_ (.A1(\decode.regfile.registers_31[9] ),
    .A2(_12709_),
    .B1(_13098_),
    .B2(_13137_),
    .C1(_12705_),
    .X(_00429_));
 sky130_fd_sc_hd__o21a_2 _17183_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[10] ),
    .B1(_13097_),
    .X(_13138_));
 sky130_fd_sc_hd__a41o_2 _17184_ (.A1(\decode.regfile.registers_20[10] ),
    .A2(_11024_),
    .A3(_12553_),
    .A4(_12554_),
    .B1(_12537_),
    .X(_13139_));
 sky130_fd_sc_hd__a41o_2 _17185_ (.A1(\decode.regfile.registers_15[10] ),
    .A2(_10611_),
    .A3(_10618_),
    .A4(_12583_),
    .B1(_12672_),
    .X(_13140_));
 sky130_fd_sc_hd__a22o_2 _17186_ (.A1(\decode.regfile.registers_7[10] ),
    .A2(_12610_),
    .B1(_12622_),
    .B2(\decode.regfile.registers_6[10] ),
    .X(_13141_));
 sky130_fd_sc_hd__a221oi_2 _17187_ (.A1(\decode.regfile.registers_2[10] ),
    .A2(_12835_),
    .B1(_12836_),
    .B2(\decode.regfile.registers_3[10] ),
    .C1(_12838_),
    .Y(_13142_));
 sky130_fd_sc_hd__a31o_2 _17188_ (.A1(_12934_),
    .A2(_10592_),
    .A3(_12558_),
    .B1(\decode.regfile.registers_0[10] ),
    .X(_13143_));
 sky130_fd_sc_hd__o211ai_2 _17189_ (.A1(\decode.regfile.registers_1[10] ),
    .A2(_12778_),
    .B1(_12830_),
    .C1(_13143_),
    .Y(_13144_));
 sky130_fd_sc_hd__buf_1 _17190_ (.A(_12934_),
    .X(_13145_));
 sky130_fd_sc_hd__a221oi_2 _17191_ (.A1(\decode.regfile.registers_4[10] ),
    .A2(_12548_),
    .B1(_13145_),
    .B2(\decode.regfile.registers_5[10] ),
    .C1(_12614_),
    .Y(_13146_));
 sky130_fd_sc_hd__a21oi_2 _17192_ (.A1(_13142_),
    .A2(_13144_),
    .B1(_13146_),
    .Y(_13147_));
 sky130_fd_sc_hd__o21ai_2 _17193_ (.A1(_13141_),
    .A2(_13147_),
    .B1(_12726_),
    .Y(_13148_));
 sky130_fd_sc_hd__a21oi_2 _17194_ (.A1(\decode.regfile.registers_8[10] ),
    .A2(_12888_),
    .B1(_12606_),
    .Y(_13149_));
 sky130_fd_sc_hd__nand2_2 _17195_ (.A(_13148_),
    .B(_13149_),
    .Y(_13150_));
 sky130_fd_sc_hd__o41a_2 _17196_ (.A1(\decode.regfile.registers_9[10] ),
    .A2(_11017_),
    .A3(_12503_),
    .A4(_12509_),
    .B1(_12652_),
    .X(_13151_));
 sky130_fd_sc_hd__a22oi_2 _17197_ (.A1(\decode.regfile.registers_10[10] ),
    .A2(_12598_),
    .B1(_13150_),
    .B2(_13151_),
    .Y(_13152_));
 sky130_fd_sc_hd__or4b_2 _17198_ (.A(_12497_),
    .B(_12503_),
    .C(_12637_),
    .D_N(\decode.regfile.registers_11[10] ),
    .X(_13153_));
 sky130_fd_sc_hd__o211ai_2 _17199_ (.A1(_12594_),
    .A2(_13152_),
    .B1(_13153_),
    .C1(_12590_),
    .Y(_13154_));
 sky130_fd_sc_hd__or4_2 _17200_ (.A(\decode.regfile.registers_12[10] ),
    .B(_12489_),
    .C(_11018_),
    .D(_12540_),
    .X(_13155_));
 sky130_fd_sc_hd__a31o_2 _17201_ (.A1(\decode.regfile.registers_13[10] ),
    .A2(_12533_),
    .A3(_12582_),
    .B1(_12662_),
    .X(_13156_));
 sky130_fd_sc_hd__a31o_2 _17202_ (.A1(_12658_),
    .A2(_13154_),
    .A3(_13155_),
    .B1(_13156_),
    .X(_13157_));
 sky130_fd_sc_hd__o221a_2 _17203_ (.A1(_12650_),
    .A2(_12772_),
    .B1(_12669_),
    .B2(\decode.regfile.registers_14[10] ),
    .C1(_13157_),
    .X(_13158_));
 sky130_fd_sc_hd__o22a_2 _17204_ (.A1(\decode.regfile.registers_16[10] ),
    .A2(_12575_),
    .B1(_13140_),
    .B2(_13158_),
    .X(_13159_));
 sky130_fd_sc_hd__a31o_2 _17205_ (.A1(_11021_),
    .A2(_12567_),
    .A3(_12586_),
    .B1(_13159_),
    .X(_13160_));
 sky130_fd_sc_hd__o211a_2 _17206_ (.A1(\decode.regfile.registers_17[10] ),
    .A2(_12579_),
    .B1(_12565_),
    .C1(_13160_),
    .X(_13161_));
 sky130_fd_sc_hd__a211o_2 _17207_ (.A1(\decode.regfile.registers_18[10] ),
    .A2(_12571_),
    .B1(_12561_),
    .C1(_13161_),
    .X(_13162_));
 sky130_fd_sc_hd__o211a_2 _17208_ (.A1(\decode.regfile.registers_19[10] ),
    .A2(_12679_),
    .B1(_12545_),
    .C1(_13162_),
    .X(_13163_));
 sky130_fd_sc_hd__buf_1 _17209_ (.A(_12755_),
    .X(_13164_));
 sky130_fd_sc_hd__or2_2 _17210_ (.A(\decode.regfile.registers_21[10] ),
    .B(_12681_),
    .X(_13165_));
 sky130_fd_sc_hd__o211a_2 _17211_ (.A1(_13139_),
    .A2(_13163_),
    .B1(_13164_),
    .C1(_13165_),
    .X(_13166_));
 sky130_fd_sc_hd__a211o_2 _17212_ (.A1(\decode.regfile.registers_22[10] ),
    .A2(_12528_),
    .B1(_13166_),
    .C1(_12687_),
    .X(_13167_));
 sky130_fd_sc_hd__buf_1 _17213_ (.A(_10936_),
    .X(_13168_));
 sky130_fd_sc_hd__or4_2 _17214_ (.A(_13081_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[10] ),
    .D(_13041_),
    .X(_13169_));
 sky130_fd_sc_hd__buf_1 _17215_ (.A(_10604_),
    .X(_13170_));
 sky130_fd_sc_hd__o2111a_2 _17216_ (.A1(_10927_),
    .A2(\decode.regfile.registers_24[10] ),
    .B1(_13170_),
    .C1(_13083_),
    .D1(_12862_),
    .X(_13171_));
 sky130_fd_sc_hd__a31o_2 _17217_ (.A1(_12516_),
    .A2(_13167_),
    .A3(_13169_),
    .B1(_13171_),
    .X(_13172_));
 sky130_fd_sc_hd__or4_2 _17218_ (.A(_12915_),
    .B(\decode.regfile.registers_25[10] ),
    .C(_13045_),
    .D(_12812_),
    .X(_13173_));
 sky130_fd_sc_hd__o2111a_2 _17219_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[10] ),
    .B1(_12814_),
    .C1(_13047_),
    .D1(_13088_),
    .X(_13174_));
 sky130_fd_sc_hd__a31o_2 _17220_ (.A1(_12695_),
    .A2(_13172_),
    .A3(_13173_),
    .B1(_13174_),
    .X(_13175_));
 sky130_fd_sc_hd__buf_1 _17221_ (.A(_12667_),
    .X(_13176_));
 sky130_fd_sc_hd__or4_2 _17222_ (.A(_13091_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[10] ),
    .D(_13050_),
    .X(_13177_));
 sky130_fd_sc_hd__o21a_2 _17223_ (.A1(_12701_),
    .A2(\decode.regfile.registers_28[10] ),
    .B1(_13093_),
    .X(_13178_));
 sky130_fd_sc_hd__a31o_2 _17224_ (.A1(_12496_),
    .A2(_13175_),
    .A3(_13177_),
    .B1(_13178_),
    .X(_13179_));
 sky130_fd_sc_hd__o221a_2 _17225_ (.A1(_13099_),
    .A2(_12768_),
    .B1(_12493_),
    .B2(\decode.regfile.registers_29[10] ),
    .C1(_13179_),
    .X(_13180_));
 sky130_fd_sc_hd__o221a_2 _17226_ (.A1(\decode.regfile.registers_31[10] ),
    .A2(_12709_),
    .B1(_13138_),
    .B2(_13180_),
    .C1(_12705_),
    .X(_00430_));
 sky130_fd_sc_hd__o21a_2 _17227_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[11] ),
    .B1(_13097_),
    .X(_13181_));
 sky130_fd_sc_hd__buf_1 _17228_ (.A(_12492_),
    .X(_13182_));
 sky130_fd_sc_hd__buf_1 _17229_ (.A(_12694_),
    .X(_13183_));
 sky130_fd_sc_hd__a41o_2 _17230_ (.A1(\decode.regfile.registers_20[11] ),
    .A2(_11024_),
    .A3(_12553_),
    .A4(_12823_),
    .B1(_12824_),
    .X(_13184_));
 sky130_fd_sc_hd__o2111a_2 _17231_ (.A1(\decode.regfile.registers_18[11] ),
    .A2(_10925_),
    .B1(_12569_),
    .C1(_11023_),
    .D1(_11008_),
    .X(_13185_));
 sky130_fd_sc_hd__a32o_2 _17232_ (.A1(_11022_),
    .A2(_12567_),
    .A3(_12586_),
    .B1(_12673_),
    .B2(\decode.regfile.registers_16[11] ),
    .X(_13186_));
 sky130_fd_sc_hd__o211a_2 _17233_ (.A1(\decode.regfile.registers_14[11] ),
    .A2(_10619_),
    .B1(_12589_),
    .C1(_10612_),
    .X(_13187_));
 sky130_fd_sc_hd__and3_2 _17234_ (.A(\decode.regfile.registers_13[11] ),
    .B(_12927_),
    .C(_12583_),
    .X(_13188_));
 sky130_fd_sc_hd__a22o_2 _17235_ (.A1(\decode.regfile.registers_11[11] ),
    .A2(_12724_),
    .B1(_12587_),
    .B2(_12550_),
    .X(_13189_));
 sky130_fd_sc_hd__o21ai_2 _17236_ (.A1(\decode.regfile.registers_9[11] ),
    .A2(_12602_),
    .B1(_12653_),
    .Y(_13190_));
 sky130_fd_sc_hd__a31o_2 _17237_ (.A1(_12934_),
    .A2(_10592_),
    .A3(_12558_),
    .B1(\decode.regfile.registers_0[11] ),
    .X(_13191_));
 sky130_fd_sc_hd__o211a_2 _17238_ (.A1(\decode.regfile.registers_1[11] ),
    .A2(_12778_),
    .B1(_12830_),
    .C1(_13191_),
    .X(_13192_));
 sky130_fd_sc_hd__a221o_2 _17239_ (.A1(\decode.regfile.registers_2[11] ),
    .A2(_12835_),
    .B1(_12836_),
    .B2(\decode.regfile.registers_3[11] ),
    .C1(_12838_),
    .X(_13193_));
 sky130_fd_sc_hd__a221o_2 _17240_ (.A1(\decode.regfile.registers_4[11] ),
    .A2(_12548_),
    .B1(_13145_),
    .B2(\decode.regfile.registers_5[11] ),
    .C1(_12614_),
    .X(_13194_));
 sky130_fd_sc_hd__o21ai_2 _17241_ (.A1(_13192_),
    .A2(_13193_),
    .B1(_13194_),
    .Y(_13195_));
 sky130_fd_sc_hd__a22oi_2 _17242_ (.A1(\decode.regfile.registers_7[11] ),
    .A2(_12611_),
    .B1(_12623_),
    .B2(\decode.regfile.registers_6[11] ),
    .Y(_13196_));
 sky130_fd_sc_hd__a21oi_2 _17243_ (.A1(_13195_),
    .A2(_13196_),
    .B1(_12888_),
    .Y(_13197_));
 sky130_fd_sc_hd__a211oi_2 _17244_ (.A1(\decode.regfile.registers_8[11] ),
    .A2(_12889_),
    .B1(_12606_),
    .C1(_13197_),
    .Y(_13198_));
 sky130_fd_sc_hd__a2bb2o_2 _17245_ (.A1_N(_13190_),
    .A2_N(_13198_),
    .B1(_12599_),
    .B2(\decode.regfile.registers_10[11] ),
    .X(_13199_));
 sky130_fd_sc_hd__o31a_2 _17246_ (.A1(_12499_),
    .A2(_12504_),
    .A3(_12650_),
    .B1(_13199_),
    .X(_13200_));
 sky130_fd_sc_hd__o221a_2 _17247_ (.A1(\decode.regfile.registers_12[11] ),
    .A2(_12591_),
    .B1(_13189_),
    .B2(_13200_),
    .C1(_12659_),
    .X(_13201_));
 sky130_fd_sc_hd__o32a_2 _17248_ (.A1(_10604_),
    .A2(_10619_),
    .A3(_12773_),
    .B1(_13188_),
    .B2(_13201_),
    .X(_13202_));
 sky130_fd_sc_hd__o221a_2 _17249_ (.A1(\decode.regfile.registers_15[11] ),
    .A2(_12874_),
    .B1(_13187_),
    .B2(_13202_),
    .C1(_12576_),
    .X(_13203_));
 sky130_fd_sc_hd__o221a_2 _17250_ (.A1(\decode.regfile.registers_17[11] ),
    .A2(_12719_),
    .B1(_13186_),
    .B2(_13203_),
    .C1(_12826_),
    .X(_13204_));
 sky130_fd_sc_hd__o221a_2 _17251_ (.A1(\decode.regfile.registers_19[11] ),
    .A2(_12678_),
    .B1(_13185_),
    .B2(_13204_),
    .C1(_12906_),
    .X(_13205_));
 sky130_fd_sc_hd__o221a_2 _17252_ (.A1(\decode.regfile.registers_21[11] ),
    .A2(_12822_),
    .B1(_13184_),
    .B2(_13205_),
    .C1(_12806_),
    .X(_13206_));
 sky130_fd_sc_hd__a211o_2 _17253_ (.A1(\decode.regfile.registers_22[11] ),
    .A2(_12528_),
    .B1(_13206_),
    .C1(_12687_),
    .X(_13207_));
 sky130_fd_sc_hd__or4_2 _17254_ (.A(_13081_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[11] ),
    .D(_13041_),
    .X(_13208_));
 sky130_fd_sc_hd__o2111a_2 _17255_ (.A1(_10927_),
    .A2(\decode.regfile.registers_24[11] ),
    .B1(_13170_),
    .C1(_13083_),
    .D1(_12862_),
    .X(_13209_));
 sky130_fd_sc_hd__a31o_2 _17256_ (.A1(_12516_),
    .A2(_13207_),
    .A3(_13208_),
    .B1(_13209_),
    .X(_13210_));
 sky130_fd_sc_hd__or4_2 _17257_ (.A(_12915_),
    .B(\decode.regfile.registers_25[11] ),
    .C(_13045_),
    .D(_12812_),
    .X(_13211_));
 sky130_fd_sc_hd__o2111a_2 _17258_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[11] ),
    .B1(_12814_),
    .C1(_13047_),
    .D1(_13088_),
    .X(_13212_));
 sky130_fd_sc_hd__a31o_2 _17259_ (.A1(_13183_),
    .A2(_13210_),
    .A3(_13211_),
    .B1(_13212_),
    .X(_13213_));
 sky130_fd_sc_hd__or4_2 _17260_ (.A(_13091_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[11] ),
    .D(_13050_),
    .X(_13214_));
 sky130_fd_sc_hd__buf_1 _17261_ (.A(_10928_),
    .X(_13215_));
 sky130_fd_sc_hd__o21a_2 _17262_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[11] ),
    .B1(_13093_),
    .X(_13216_));
 sky130_fd_sc_hd__a31o_2 _17263_ (.A1(_12496_),
    .A2(_13213_),
    .A3(_13214_),
    .B1(_13216_),
    .X(_13217_));
 sky130_fd_sc_hd__o221a_2 _17264_ (.A1(_13099_),
    .A2(_12768_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[11] ),
    .C1(_13217_),
    .X(_13218_));
 sky130_fd_sc_hd__buf_1 _17265_ (.A(_12704_),
    .X(_13219_));
 sky130_fd_sc_hd__o221a_2 _17266_ (.A1(_12708_),
    .A2(\decode.regfile.registers_31[11] ),
    .B1(_13181_),
    .B2(_13218_),
    .C1(_13219_),
    .X(_00431_));
 sky130_fd_sc_hd__o21a_2 _17267_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[12] ),
    .B1(_13097_),
    .X(_13220_));
 sky130_fd_sc_hd__buf_1 _17268_ (.A(_12495_),
    .X(_13221_));
 sky130_fd_sc_hd__a41o_2 _17269_ (.A1(\decode.regfile.registers_20[12] ),
    .A2(_11024_),
    .A3(_12553_),
    .A4(_12823_),
    .B1(_12824_),
    .X(_13222_));
 sky130_fd_sc_hd__and4b_2 _17270_ (.A_N(_10923_),
    .B(_12876_),
    .C(\decode.regfile.registers_14[12] ),
    .D(_12555_),
    .X(_13223_));
 sky130_fd_sc_hd__a31o_2 _17271_ (.A1(\decode.regfile.registers_12[12] ),
    .A2(_12551_),
    .A3(_12583_),
    .B1(_12775_),
    .X(_13224_));
 sky130_fd_sc_hd__o21ai_2 _17272_ (.A1(\decode.regfile.registers_9[12] ),
    .A2(_12603_),
    .B1(_12790_),
    .Y(_13225_));
 sky130_fd_sc_hd__a221o_2 _17273_ (.A1(\decode.regfile.registers_4[12] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[12] ),
    .C1(_12737_),
    .X(_13226_));
 sky130_fd_sc_hd__a31o_2 _17274_ (.A1(_12530_),
    .A2(_12616_),
    .A3(_12557_),
    .B1(\decode.regfile.registers_0[12] ),
    .X(_13227_));
 sky130_fd_sc_hd__o211a_2 _17275_ (.A1(\decode.regfile.registers_1[12] ),
    .A2(_12631_),
    .B1(_12633_),
    .C1(_13227_),
    .X(_13228_));
 sky130_fd_sc_hd__a211o_2 _17276_ (.A1(\decode.regfile.registers_2[12] ),
    .A2(_12835_),
    .B1(_12836_),
    .C1(_13228_),
    .X(_13229_));
 sky130_fd_sc_hd__o221a_2 _17277_ (.A1(_10610_),
    .A2(_12626_),
    .B1(_12629_),
    .B2(\decode.regfile.registers_3[12] ),
    .C1(_13229_),
    .X(_13230_));
 sky130_fd_sc_hd__o22ai_2 _17278_ (.A1(\decode.regfile.registers_6[12] ),
    .A2(_12735_),
    .B1(_13226_),
    .B2(_13230_),
    .Y(_13231_));
 sky130_fd_sc_hd__o21ai_2 _17279_ (.A1(_12649_),
    .A2(_12615_),
    .B1(_13231_),
    .Y(_13232_));
 sky130_fd_sc_hd__o32a_2 _17280_ (.A1(_12497_),
    .A2(_12539_),
    .A3(_12503_),
    .B1(\decode.regfile.registers_7[12] ),
    .B2(_12645_),
    .X(_13233_));
 sky130_fd_sc_hd__a41o_2 _17281_ (.A1(\decode.regfile.registers_8[12] ),
    .A2(_12776_),
    .A3(_12549_),
    .A4(_12604_),
    .B1(_12606_),
    .X(_13234_));
 sky130_fd_sc_hd__a21oi_2 _17282_ (.A1(_13232_),
    .A2(_13233_),
    .B1(_13234_),
    .Y(_13235_));
 sky130_fd_sc_hd__a21oi_2 _17283_ (.A1(\decode.regfile.registers_10[12] ),
    .A2(_12600_),
    .B1(_12724_),
    .Y(_13236_));
 sky130_fd_sc_hd__o21ai_2 _17284_ (.A1(_13225_),
    .A2(_13235_),
    .B1(_13236_),
    .Y(_13237_));
 sky130_fd_sc_hd__o221a_2 _17285_ (.A1(\decode.regfile.registers_11[12] ),
    .A2(_12878_),
    .B1(_12772_),
    .B2(_12541_),
    .C1(_13237_),
    .X(_13238_));
 sky130_fd_sc_hd__o221a_2 _17286_ (.A1(\decode.regfile.registers_13[12] ),
    .A2(_12659_),
    .B1(_13224_),
    .B2(_13238_),
    .C1(_12984_),
    .X(_13239_));
 sky130_fd_sc_hd__o31a_2 _17287_ (.A1(\decode.regfile.registers_15[12] ),
    .A2(_12666_),
    .A3(_12723_),
    .B1(_12575_),
    .X(_13240_));
 sky130_fd_sc_hd__o31a_2 _17288_ (.A1(_12585_),
    .A2(_13223_),
    .A3(_13239_),
    .B1(_13240_),
    .X(_13241_));
 sky130_fd_sc_hd__a211o_2 _17289_ (.A1(\decode.regfile.registers_16[12] ),
    .A2(_12674_),
    .B1(_12901_),
    .C1(_13241_),
    .X(_13242_));
 sky130_fd_sc_hd__o21a_2 _17290_ (.A1(\decode.regfile.registers_17[12] ),
    .A2(_12719_),
    .B1(_12565_),
    .X(_13243_));
 sky130_fd_sc_hd__o2111a_2 _17291_ (.A1(\decode.regfile.registers_18[12] ),
    .A2(_10924_),
    .B1(_12568_),
    .C1(_12524_),
    .D1(_11008_),
    .X(_13244_));
 sky130_fd_sc_hd__a21o_2 _17292_ (.A1(_13242_),
    .A2(_13243_),
    .B1(_13244_),
    .X(_13245_));
 sky130_fd_sc_hd__o211a_2 _17293_ (.A1(\decode.regfile.registers_19[12] ),
    .A2(_12679_),
    .B1(_12906_),
    .C1(_13245_),
    .X(_13246_));
 sky130_fd_sc_hd__o221a_2 _17294_ (.A1(\decode.regfile.registers_21[12] ),
    .A2(_12716_),
    .B1(_13222_),
    .B2(_13246_),
    .C1(_12806_),
    .X(_13247_));
 sky130_fd_sc_hd__a211o_2 _17295_ (.A1(\decode.regfile.registers_22[12] ),
    .A2(_12528_),
    .B1(_13247_),
    .C1(_12687_),
    .X(_13248_));
 sky130_fd_sc_hd__or4_2 _17296_ (.A(_13081_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[12] ),
    .D(_13041_),
    .X(_13249_));
 sky130_fd_sc_hd__buf_1 _17297_ (.A(_10926_),
    .X(_13250_));
 sky130_fd_sc_hd__o2111a_2 _17298_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[12] ),
    .B1(_13170_),
    .C1(_13083_),
    .D1(_12862_),
    .X(_13251_));
 sky130_fd_sc_hd__a31o_2 _17299_ (.A1(_12516_),
    .A2(_13248_),
    .A3(_13249_),
    .B1(_13251_),
    .X(_13252_));
 sky130_fd_sc_hd__or4_2 _17300_ (.A(_12915_),
    .B(\decode.regfile.registers_25[12] ),
    .C(_13045_),
    .D(_12812_),
    .X(_13253_));
 sky130_fd_sc_hd__buf_1 _17301_ (.A(_12759_),
    .X(_13254_));
 sky130_fd_sc_hd__o2111a_2 _17302_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[12] ),
    .B1(_13254_),
    .C1(_13047_),
    .D1(_13088_),
    .X(_13255_));
 sky130_fd_sc_hd__a31o_2 _17303_ (.A1(_13183_),
    .A2(_13252_),
    .A3(_13253_),
    .B1(_13255_),
    .X(_13256_));
 sky130_fd_sc_hd__or4_2 _17304_ (.A(_13091_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[12] ),
    .D(_13050_),
    .X(_13257_));
 sky130_fd_sc_hd__o21a_2 _17305_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[12] ),
    .B1(_13093_),
    .X(_13258_));
 sky130_fd_sc_hd__a31o_2 _17306_ (.A1(_13221_),
    .A2(_13256_),
    .A3(_13257_),
    .B1(_13258_),
    .X(_13259_));
 sky130_fd_sc_hd__o221a_2 _17307_ (.A1(_13099_),
    .A2(_12768_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[12] ),
    .C1(_13259_),
    .X(_13260_));
 sky130_fd_sc_hd__o221a_2 _17308_ (.A1(\decode.regfile.registers_31[12] ),
    .A2(_12709_),
    .B1(_13220_),
    .B2(_13260_),
    .C1(_13219_),
    .X(_00432_));
 sky130_fd_sc_hd__o21a_2 _17309_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[13] ),
    .B1(_13097_),
    .X(_13261_));
 sky130_fd_sc_hd__buf_1 _17310_ (.A(_12767_),
    .X(_13262_));
 sky130_fd_sc_hd__a41o_2 _17311_ (.A1(\decode.regfile.registers_20[13] ),
    .A2(_11024_),
    .A3(_12553_),
    .A4(_12823_),
    .B1(_12537_),
    .X(_13263_));
 sky130_fd_sc_hd__a21o_2 _17312_ (.A1(\decode.regfile.registers_18[13] ),
    .A2(_12571_),
    .B1(_12561_),
    .X(_13264_));
 sky130_fd_sc_hd__and4_2 _17313_ (.A(\decode.regfile.registers_17[13] ),
    .B(_11022_),
    .C(_12567_),
    .D(_12586_),
    .X(_13265_));
 sky130_fd_sc_hd__nor2_2 _17314_ (.A(\decode.regfile.registers_11[13] ),
    .B(_12878_),
    .Y(_13266_));
 sky130_fd_sc_hd__a221oi_2 _17315_ (.A1(\decode.regfile.registers_7[13] ),
    .A2(_12611_),
    .B1(_12623_),
    .B2(\decode.regfile.registers_6[13] ),
    .C1(_12888_),
    .Y(_13267_));
 sky130_fd_sc_hd__a31o_2 _17316_ (.A1(\decode.regfile.registers_3[13] ),
    .A2(_10616_),
    .A3(_12729_),
    .B1(_12838_),
    .X(_13268_));
 sky130_fd_sc_hd__and2b_2 _17317_ (.A_N(_12882_),
    .B(\decode.regfile.registers_2[13] ),
    .X(_13269_));
 sky130_fd_sc_hd__mux2_2 _17318_ (.A0(\decode.regfile.registers_1[13] ),
    .A1(\decode.regfile.registers_0[13] ),
    .S(_12778_),
    .X(_13270_));
 sky130_fd_sc_hd__o22a_2 _17319_ (.A1(_12830_),
    .A2(_13269_),
    .B1(_12835_),
    .B2(_13270_),
    .X(_13271_));
 sky130_fd_sc_hd__a221o_2 _17320_ (.A1(\decode.regfile.registers_4[13] ),
    .A2(_12549_),
    .B1(_12532_),
    .B2(\decode.regfile.registers_5[13] ),
    .C1(_12626_),
    .X(_13272_));
 sky130_fd_sc_hd__o21ai_2 _17321_ (.A1(_13268_),
    .A2(_13271_),
    .B1(_13272_),
    .Y(_13273_));
 sky130_fd_sc_hd__o2bb2ai_2 _17322_ (.A1_N(_13267_),
    .A2_N(_13273_),
    .B1(_12892_),
    .B2(\decode.regfile.registers_8[13] ),
    .Y(_13274_));
 sky130_fd_sc_hd__nand2_2 _17323_ (.A(_12603_),
    .B(_13274_),
    .Y(_13275_));
 sky130_fd_sc_hd__o41a_2 _17324_ (.A1(\decode.regfile.registers_9[13] ),
    .A2(_11018_),
    .A3(_12977_),
    .A4(_12510_),
    .B1(_12653_),
    .X(_13276_));
 sky130_fd_sc_hd__a221oi_2 _17325_ (.A1(\decode.regfile.registers_10[13] ),
    .A2(_12600_),
    .B1(_13275_),
    .B2(_13276_),
    .C1(_12724_),
    .Y(_13277_));
 sky130_fd_sc_hd__o21ai_2 _17326_ (.A1(_13266_),
    .A2(_13277_),
    .B1(_12591_),
    .Y(_13278_));
 sky130_fd_sc_hd__o32a_2 _17327_ (.A1(_12499_),
    .A2(_12490_),
    .A3(_12511_),
    .B1(\decode.regfile.registers_12[13] ),
    .B2(_12745_),
    .X(_13279_));
 sky130_fd_sc_hd__a221o_2 _17328_ (.A1(\decode.regfile.registers_13[13] ),
    .A2(_12775_),
    .B1(_13278_),
    .B2(_13279_),
    .C1(_12663_),
    .X(_13280_));
 sky130_fd_sc_hd__or4_2 _17329_ (.A(\decode.regfile.registers_14[13] ),
    .B(_10604_),
    .C(_10618_),
    .D(_12772_),
    .X(_13281_));
 sky130_fd_sc_hd__a41o_2 _17330_ (.A1(\decode.regfile.registers_15[13] ),
    .A2(_12555_),
    .A3(_10923_),
    .A4(_12876_),
    .B1(_13031_),
    .X(_13282_));
 sky130_fd_sc_hd__a31o_2 _17331_ (.A1(_12874_),
    .A2(_13280_),
    .A3(_13281_),
    .B1(_13282_),
    .X(_13283_));
 sky130_fd_sc_hd__o211a_2 _17332_ (.A1(\decode.regfile.registers_16[13] ),
    .A2(_12576_),
    .B1(_12579_),
    .C1(_13283_),
    .X(_13284_));
 sky130_fd_sc_hd__o21a_2 _17333_ (.A1(_13265_),
    .A2(_13284_),
    .B1(_12566_),
    .X(_13285_));
 sky130_fd_sc_hd__o221a_2 _17334_ (.A1(\decode.regfile.registers_19[13] ),
    .A2(_12679_),
    .B1(_13264_),
    .B2(_13285_),
    .C1(_12545_),
    .X(_13286_));
 sky130_fd_sc_hd__or2_2 _17335_ (.A(\decode.regfile.registers_21[13] ),
    .B(_12681_),
    .X(_13287_));
 sky130_fd_sc_hd__o211a_2 _17336_ (.A1(_13263_),
    .A2(_13286_),
    .B1(_13164_),
    .C1(_13287_),
    .X(_13288_));
 sky130_fd_sc_hd__buf_1 _17337_ (.A(_12686_),
    .X(_13289_));
 sky130_fd_sc_hd__a211o_2 _17338_ (.A1(\decode.regfile.registers_22[13] ),
    .A2(_12528_),
    .B1(_13288_),
    .C1(_13289_),
    .X(_13290_));
 sky130_fd_sc_hd__or4_2 _17339_ (.A(_13081_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[13] ),
    .D(_13041_),
    .X(_13291_));
 sky130_fd_sc_hd__o2111a_2 _17340_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[13] ),
    .B1(_13170_),
    .C1(_13083_),
    .D1(_12862_),
    .X(_13292_));
 sky130_fd_sc_hd__a31o_2 _17341_ (.A1(_12516_),
    .A2(_13290_),
    .A3(_13291_),
    .B1(_13292_),
    .X(_13293_));
 sky130_fd_sc_hd__buf_1 _17342_ (.A(_12512_),
    .X(_13294_));
 sky130_fd_sc_hd__or4_2 _17343_ (.A(_12915_),
    .B(\decode.regfile.registers_25[13] ),
    .C(_13045_),
    .D(_13294_),
    .X(_13295_));
 sky130_fd_sc_hd__o2111a_2 _17344_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[13] ),
    .B1(_13254_),
    .C1(_13047_),
    .D1(_13088_),
    .X(_13296_));
 sky130_fd_sc_hd__a31o_2 _17345_ (.A1(_13183_),
    .A2(_13293_),
    .A3(_13295_),
    .B1(_13296_),
    .X(_13297_));
 sky130_fd_sc_hd__or4_2 _17346_ (.A(_13091_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[13] ),
    .D(_13050_),
    .X(_13298_));
 sky130_fd_sc_hd__o21a_2 _17347_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[13] ),
    .B1(_13093_),
    .X(_13299_));
 sky130_fd_sc_hd__a31o_2 _17348_ (.A1(_13221_),
    .A2(_13297_),
    .A3(_13298_),
    .B1(_13299_),
    .X(_13300_));
 sky130_fd_sc_hd__o221a_2 _17349_ (.A1(_13099_),
    .A2(_13262_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[13] ),
    .C1(_13300_),
    .X(_13301_));
 sky130_fd_sc_hd__o221a_2 _17350_ (.A1(_12708_),
    .A2(\decode.regfile.registers_31[13] ),
    .B1(_13261_),
    .B2(_13301_),
    .C1(_13219_),
    .X(_00433_));
 sky130_fd_sc_hd__o21a_2 _17351_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[14] ),
    .B1(_13097_),
    .X(_13302_));
 sky130_fd_sc_hd__o21a_2 _17352_ (.A1(_12701_),
    .A2(\decode.regfile.registers_28[14] ),
    .B1(_12698_),
    .X(_13303_));
 sky130_fd_sc_hd__and3_2 _17353_ (.A(_11025_),
    .B(_12690_),
    .C(_12535_),
    .X(_13304_));
 sky130_fd_sc_hd__o2111a_2 _17354_ (.A1(_10926_),
    .A2(\decode.regfile.registers_22[14] ),
    .B1(_12554_),
    .C1(_11009_),
    .D1(_12546_),
    .X(_13305_));
 sky130_fd_sc_hd__a21o_2 _17355_ (.A1(\decode.regfile.registers_18[14] ),
    .A2(_12570_),
    .B1(_12560_),
    .X(_13306_));
 sky130_fd_sc_hd__a32o_2 _17356_ (.A1(_11021_),
    .A2(_12559_),
    .A3(_12534_),
    .B1(_13031_),
    .B2(\decode.regfile.registers_16[14] ),
    .X(_13307_));
 sky130_fd_sc_hd__a31o_2 _17357_ (.A1(\decode.regfile.registers_13[14] ),
    .A2(_12533_),
    .A3(_12587_),
    .B1(_12662_),
    .X(_13308_));
 sky130_fd_sc_hd__a22o_2 _17358_ (.A1(\decode.regfile.registers_11[14] ),
    .A2(_12594_),
    .B1(_12582_),
    .B2(_12550_),
    .X(_13309_));
 sky130_fd_sc_hd__a41o_2 _17359_ (.A1(\decode.regfile.registers_8[14] ),
    .A2(_10593_),
    .A3(_12549_),
    .A4(_12592_),
    .B1(_12605_),
    .X(_13310_));
 sky130_fd_sc_hd__a221oi_2 _17360_ (.A1(\decode.regfile.registers_4[14] ),
    .A2(_12617_),
    .B1(_12619_),
    .B2(\decode.regfile.registers_5[14] ),
    .C1(_12622_),
    .Y(_13311_));
 sky130_fd_sc_hd__a31o_2 _17361_ (.A1(\decode.regfile.registers_2[14] ),
    .A2(_10608_),
    .A3(_12635_),
    .B1(_12638_),
    .X(_13312_));
 sky130_fd_sc_hd__a31o_2 _17362_ (.A1(_12530_),
    .A2(_10591_),
    .A3(_12557_),
    .B1(\decode.regfile.registers_0[14] ),
    .X(_13313_));
 sky130_fd_sc_hd__o221a_2 _17363_ (.A1(\decode.regfile.registers_1[14] ),
    .A2(_12630_),
    .B1(_12829_),
    .B2(_10614_),
    .C1(_13313_),
    .X(_13314_));
 sky130_fd_sc_hd__o22a_2 _17364_ (.A1(\decode.regfile.registers_3[14] ),
    .A2(_12627_),
    .B1(_10608_),
    .B2(_12613_),
    .X(_13315_));
 sky130_fd_sc_hd__o21ai_2 _17365_ (.A1(_13312_),
    .A2(_13314_),
    .B1(_13315_),
    .Y(_13316_));
 sky130_fd_sc_hd__o2bb2a_2 _17366_ (.A1_N(_13311_),
    .A2_N(_13316_),
    .B1(_12735_),
    .B2(\decode.regfile.registers_6[14] ),
    .X(_13317_));
 sky130_fd_sc_hd__o32a_2 _17367_ (.A1(_11016_),
    .A2(_12539_),
    .A3(_12502_),
    .B1(\decode.regfile.registers_7[14] ),
    .B2(_12644_),
    .X(_13318_));
 sky130_fd_sc_hd__o21a_2 _17368_ (.A1(_12611_),
    .A2(_13317_),
    .B1(_13318_),
    .X(_13319_));
 sky130_fd_sc_hd__o22a_2 _17369_ (.A1(\decode.regfile.registers_9[14] ),
    .A2(_12602_),
    .B1(_13310_),
    .B2(_13319_),
    .X(_13320_));
 sky130_fd_sc_hd__o32a_2 _17370_ (.A1(_11018_),
    .A2(_12977_),
    .A3(_12649_),
    .B1(\decode.regfile.registers_10[14] ),
    .B2(_12652_),
    .X(_13321_));
 sky130_fd_sc_hd__o21a_2 _17371_ (.A1(_12599_),
    .A2(_13320_),
    .B1(_13321_),
    .X(_13322_));
 sky130_fd_sc_hd__o221a_2 _17372_ (.A1(\decode.regfile.registers_12[14] ),
    .A2(_12745_),
    .B1(_13309_),
    .B2(_13322_),
    .C1(_12658_),
    .X(_13323_));
 sky130_fd_sc_hd__o22a_2 _17373_ (.A1(\decode.regfile.registers_14[14] ),
    .A2(_12669_),
    .B1(_13308_),
    .B2(_13323_),
    .X(_13324_));
 sky130_fd_sc_hd__o31a_2 _17374_ (.A1(\decode.regfile.registers_15[14] ),
    .A2(_12650_),
    .A3(_12723_),
    .B1(_12574_),
    .X(_13325_));
 sky130_fd_sc_hd__o21a_2 _17375_ (.A1(_12584_),
    .A2(_13324_),
    .B1(_13325_),
    .X(_13326_));
 sky130_fd_sc_hd__o221a_2 _17376_ (.A1(\decode.regfile.registers_17[14] ),
    .A2(_12578_),
    .B1(_13307_),
    .B2(_13326_),
    .C1(_12564_),
    .X(_13327_));
 sky130_fd_sc_hd__o221a_2 _17377_ (.A1(\decode.regfile.registers_19[14] ),
    .A2(_12677_),
    .B1(_13306_),
    .B2(_13327_),
    .C1(_12543_),
    .X(_13328_));
 sky130_fd_sc_hd__a211o_2 _17378_ (.A1(\decode.regfile.registers_20[14] ),
    .A2(_12770_),
    .B1(_13328_),
    .C1(_12537_),
    .X(_13329_));
 sky130_fd_sc_hd__o211a_2 _17379_ (.A1(_12716_),
    .A2(\decode.regfile.registers_21[14] ),
    .B1(_12909_),
    .C1(_13329_),
    .X(_13330_));
 sky130_fd_sc_hd__o221a_2 _17380_ (.A1(\decode.regfile.registers_23[14] ),
    .A2(_12714_),
    .B1(_13305_),
    .B2(_13330_),
    .C1(_12515_),
    .X(_13331_));
 sky130_fd_sc_hd__a211o_2 _17381_ (.A1(\decode.regfile.registers_24[14] ),
    .A2(_12691_),
    .B1(_13304_),
    .C1(_13331_),
    .X(_13332_));
 sky130_fd_sc_hd__or4_2 _17382_ (.A(_10938_),
    .B(\decode.regfile.registers_25[14] ),
    .C(_12505_),
    .D(_12811_),
    .X(_13333_));
 sky130_fd_sc_hd__o2111a_2 _17383_ (.A1(_12494_),
    .A2(\decode.regfile.registers_26[14] ),
    .B1(_13002_),
    .C1(_11010_),
    .D1(_11026_),
    .X(_13334_));
 sky130_fd_sc_hd__a31o_2 _17384_ (.A1(_12694_),
    .A2(_13332_),
    .A3(_13333_),
    .B1(_13334_),
    .X(_13335_));
 sky130_fd_sc_hd__o311a_2 _17385_ (.A1(\decode.regfile.registers_27[14] ),
    .A2(_12507_),
    .A3(_12520_),
    .B1(_12495_),
    .C1(_13335_),
    .X(_13336_));
 sky130_fd_sc_hd__o221a_2 _17386_ (.A1(_12492_),
    .A2(\decode.regfile.registers_29[14] ),
    .B1(_13303_),
    .B2(_13336_),
    .C1(_12702_),
    .X(_13337_));
 sky130_fd_sc_hd__o221a_2 _17387_ (.A1(\decode.regfile.registers_31[14] ),
    .A2(_12709_),
    .B1(_13302_),
    .B2(_13337_),
    .C1(_13219_),
    .X(_00434_));
 sky130_fd_sc_hd__o21a_2 _17388_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[15] ),
    .B1(_13097_),
    .X(_13338_));
 sky130_fd_sc_hd__buf_1 _17389_ (.A(_12515_),
    .X(_13339_));
 sky130_fd_sc_hd__a41o_2 _17390_ (.A1(\decode.regfile.registers_15[15] ),
    .A2(_10612_),
    .A3(_10619_),
    .A4(_12589_),
    .B1(_13031_),
    .X(_13340_));
 sky130_fd_sc_hd__a41o_2 _17391_ (.A1(\decode.regfile.registers_9[15] ),
    .A2(_12776_),
    .A3(_12604_),
    .A4(_12532_),
    .B1(_12599_),
    .X(_13341_));
 sky130_fd_sc_hd__a221o_2 _17392_ (.A1(\decode.regfile.registers_4[15] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[15] ),
    .C1(_12622_),
    .X(_13342_));
 sky130_fd_sc_hd__a31o_2 _17393_ (.A1(\decode.regfile.registers_2[15] ),
    .A2(_10608_),
    .A3(_12636_),
    .B1(_12639_),
    .X(_13343_));
 sky130_fd_sc_hd__a31o_2 _17394_ (.A1(_12934_),
    .A2(_12616_),
    .A3(_12558_),
    .B1(\decode.regfile.registers_0[15] ),
    .X(_13344_));
 sky130_fd_sc_hd__o221a_2 _17395_ (.A1(\decode.regfile.registers_1[15] ),
    .A2(_12932_),
    .B1(_12933_),
    .B2(_10615_),
    .C1(_13344_),
    .X(_13345_));
 sky130_fd_sc_hd__o22a_2 _17396_ (.A1(\decode.regfile.registers_3[15] ),
    .A2(_12628_),
    .B1(_10609_),
    .B2(_12625_),
    .X(_13346_));
 sky130_fd_sc_hd__o21a_2 _17397_ (.A1(_13343_),
    .A2(_13345_),
    .B1(_13346_),
    .X(_13347_));
 sky130_fd_sc_hd__o22ai_2 _17398_ (.A1(\decode.regfile.registers_6[15] ),
    .A2(_12880_),
    .B1(_13342_),
    .B2(_13347_),
    .Y(_13348_));
 sky130_fd_sc_hd__a21oi_2 _17399_ (.A1(\decode.regfile.registers_7[15] ),
    .A2(_12611_),
    .B1(_12888_),
    .Y(_13349_));
 sky130_fd_sc_hd__o21ai_2 _17400_ (.A1(_12611_),
    .A2(_13348_),
    .B1(_13349_),
    .Y(_13350_));
 sky130_fd_sc_hd__o211a_2 _17401_ (.A1(\decode.regfile.registers_8[15] ),
    .A2(_12892_),
    .B1(_12602_),
    .C1(_13350_),
    .X(_13351_));
 sky130_fd_sc_hd__o221ai_2 _17402_ (.A1(\decode.regfile.registers_10[15] ),
    .A2(_12790_),
    .B1(_13341_),
    .B2(_13351_),
    .C1(_12792_),
    .Y(_13352_));
 sky130_fd_sc_hd__or4b_2 _17403_ (.A(_12498_),
    .B(_12504_),
    .C(_12649_),
    .D_N(\decode.regfile.registers_11[15] ),
    .X(_13353_));
 sky130_fd_sc_hd__o211ai_2 _17404_ (.A1(_12541_),
    .A2(_12772_),
    .B1(_13352_),
    .C1(_13353_),
    .Y(_13354_));
 sky130_fd_sc_hd__o32a_2 _17405_ (.A1(_12499_),
    .A2(_12489_),
    .A3(_12511_),
    .B1(\decode.regfile.registers_12[15] ),
    .B2(_12745_),
    .X(_13355_));
 sky130_fd_sc_hd__a221o_2 _17406_ (.A1(\decode.regfile.registers_13[15] ),
    .A2(_12775_),
    .B1(_13354_),
    .B2(_13355_),
    .C1(_12663_),
    .X(_13356_));
 sky130_fd_sc_hd__o221a_2 _17407_ (.A1(_12666_),
    .A2(_12773_),
    .B1(_12984_),
    .B2(\decode.regfile.registers_14[15] ),
    .C1(_13356_),
    .X(_13357_));
 sky130_fd_sc_hd__o22ai_2 _17408_ (.A1(\decode.regfile.registers_16[15] ),
    .A2(_13011_),
    .B1(_13340_),
    .B2(_13357_),
    .Y(_13358_));
 sky130_fd_sc_hd__nand2_2 _17409_ (.A(_12719_),
    .B(_13358_),
    .Y(_13359_));
 sky130_fd_sc_hd__o21a_2 _17410_ (.A1(\decode.regfile.registers_17[15] ),
    .A2(_12579_),
    .B1(_12565_),
    .X(_13360_));
 sky130_fd_sc_hd__a221o_2 _17411_ (.A1(\decode.regfile.registers_18[15] ),
    .A2(_12571_),
    .B1(_13359_),
    .B2(_13360_),
    .C1(_12561_),
    .X(_13361_));
 sky130_fd_sc_hd__o41a_2 _17412_ (.A1(\decode.regfile.registers_19[15] ),
    .A2(_10599_),
    .A3(_10589_),
    .A4(_12518_),
    .B1(_12543_),
    .X(_13362_));
 sky130_fd_sc_hd__a221o_2 _17413_ (.A1(\decode.regfile.registers_20[15] ),
    .A2(_12770_),
    .B1(_13361_),
    .B2(_13362_),
    .C1(_12537_),
    .X(_13363_));
 sky130_fd_sc_hd__o211a_2 _17414_ (.A1(_12822_),
    .A2(\decode.regfile.registers_21[15] ),
    .B1(_13164_),
    .C1(_13363_),
    .X(_13364_));
 sky130_fd_sc_hd__a211o_2 _17415_ (.A1(\decode.regfile.registers_22[15] ),
    .A2(_13100_),
    .B1(_13364_),
    .C1(_13289_),
    .X(_13365_));
 sky130_fd_sc_hd__or4_2 _17416_ (.A(_13081_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[15] ),
    .D(_13041_),
    .X(_13366_));
 sky130_fd_sc_hd__buf_1 _17417_ (.A(_12546_),
    .X(_13367_));
 sky130_fd_sc_hd__o2111a_2 _17418_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[15] ),
    .B1(_13170_),
    .C1(_13083_),
    .D1(_13367_),
    .X(_13368_));
 sky130_fd_sc_hd__a31o_2 _17419_ (.A1(_13339_),
    .A2(_13365_),
    .A3(_13366_),
    .B1(_13368_),
    .X(_13369_));
 sky130_fd_sc_hd__or4_2 _17420_ (.A(_12915_),
    .B(\decode.regfile.registers_25[15] ),
    .C(_13045_),
    .D(_13294_),
    .X(_13370_));
 sky130_fd_sc_hd__o2111a_2 _17421_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[15] ),
    .B1(_13254_),
    .C1(_13047_),
    .D1(_13088_),
    .X(_13371_));
 sky130_fd_sc_hd__a31o_2 _17422_ (.A1(_13183_),
    .A2(_13369_),
    .A3(_13370_),
    .B1(_13371_),
    .X(_13372_));
 sky130_fd_sc_hd__or4_2 _17423_ (.A(_13091_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[15] ),
    .D(_13050_),
    .X(_13373_));
 sky130_fd_sc_hd__o21a_2 _17424_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[15] ),
    .B1(_13093_),
    .X(_13374_));
 sky130_fd_sc_hd__a31o_2 _17425_ (.A1(_13221_),
    .A2(_13372_),
    .A3(_13373_),
    .B1(_13374_),
    .X(_13375_));
 sky130_fd_sc_hd__o221a_2 _17426_ (.A1(_13099_),
    .A2(_13262_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[15] ),
    .C1(_13375_),
    .X(_13376_));
 sky130_fd_sc_hd__o221a_2 _17427_ (.A1(\decode.regfile.registers_31[15] ),
    .A2(_12709_),
    .B1(_13338_),
    .B2(_13376_),
    .C1(_13219_),
    .X(_00435_));
 sky130_fd_sc_hd__o21a_2 _17428_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[16] ),
    .B1(_13097_),
    .X(_13377_));
 sky130_fd_sc_hd__a41o_2 _17429_ (.A1(\decode.regfile.registers_20[16] ),
    .A2(_11024_),
    .A3(_12552_),
    .A4(_12823_),
    .B1(_12824_),
    .X(_13378_));
 sky130_fd_sc_hd__a32o_2 _17430_ (.A1(_11021_),
    .A2(_12559_),
    .A3(_12534_),
    .B1(_12673_),
    .B2(\decode.regfile.registers_16[16] ),
    .X(_13379_));
 sky130_fd_sc_hd__a41o_2 _17431_ (.A1(\decode.regfile.registers_9[16] ),
    .A2(_12776_),
    .A3(_12592_),
    .A4(_12532_),
    .B1(_12598_),
    .X(_13380_));
 sky130_fd_sc_hd__o2bb2a_2 _17432_ (.A1_N(\decode.regfile.registers_3[16] ),
    .A2_N(_12639_),
    .B1(_10609_),
    .B2(_12625_),
    .X(_13381_));
 sky130_fd_sc_hd__inv_2 _17433_ (.A(\decode.regfile.registers_1[16] ),
    .Y(_13382_));
 sky130_fd_sc_hd__nand2_2 _17434_ (.A(_12631_),
    .B(\decode.regfile.registers_0[16] ),
    .Y(_13383_));
 sky130_fd_sc_hd__o221ai_2 _17435_ (.A1(_13382_),
    .A2(_12932_),
    .B1(_10615_),
    .B2(_12933_),
    .C1(_13383_),
    .Y(_13384_));
 sky130_fd_sc_hd__o211ai_2 _17436_ (.A1(\decode.regfile.registers_2[16] ),
    .A2(_12634_),
    .B1(_12628_),
    .C1(_13384_),
    .Y(_13385_));
 sky130_fd_sc_hd__a221oi_2 _17437_ (.A1(\decode.regfile.registers_4[16] ),
    .A2(_12548_),
    .B1(_13145_),
    .B2(\decode.regfile.registers_5[16] ),
    .C1(_12614_),
    .Y(_13386_));
 sky130_fd_sc_hd__a21oi_2 _17438_ (.A1(_13381_),
    .A2(_13385_),
    .B1(_13386_),
    .Y(_13387_));
 sky130_fd_sc_hd__a221oi_2 _17439_ (.A1(\decode.regfile.registers_7[16] ),
    .A2(_12611_),
    .B1(_12623_),
    .B2(\decode.regfile.registers_6[16] ),
    .C1(_13387_),
    .Y(_13388_));
 sky130_fd_sc_hd__o21ai_2 _17440_ (.A1(\decode.regfile.registers_8[16] ),
    .A2(_12726_),
    .B1(_12601_),
    .Y(_13389_));
 sky130_fd_sc_hd__a21oi_2 _17441_ (.A1(_13388_),
    .A2(_12726_),
    .B1(_13389_),
    .Y(_13390_));
 sky130_fd_sc_hd__o22ai_2 _17442_ (.A1(\decode.regfile.registers_10[16] ),
    .A2(_12653_),
    .B1(_13380_),
    .B2(_13390_),
    .Y(_13391_));
 sky130_fd_sc_hd__or4b_2 _17443_ (.A(_11018_),
    .B(_12977_),
    .C(_12637_),
    .D_N(\decode.regfile.registers_11[16] ),
    .X(_13392_));
 sky130_fd_sc_hd__o221ai_2 _17444_ (.A1(_12540_),
    .A2(_12722_),
    .B1(_12724_),
    .B2(_13391_),
    .C1(_13392_),
    .Y(_13393_));
 sky130_fd_sc_hd__o32a_2 _17445_ (.A1(_12498_),
    .A2(_12489_),
    .A3(_12511_),
    .B1(\decode.regfile.registers_12[16] ),
    .B2(_12590_),
    .X(_13394_));
 sky130_fd_sc_hd__a221o_2 _17446_ (.A1(\decode.regfile.registers_13[16] ),
    .A2(_12774_),
    .B1(_13393_),
    .B2(_13394_),
    .C1(_12662_),
    .X(_13395_));
 sky130_fd_sc_hd__or4_2 _17447_ (.A(\decode.regfile.registers_14[16] ),
    .B(_10603_),
    .C(_10618_),
    .D(_12722_),
    .X(_13396_));
 sky130_fd_sc_hd__a32o_2 _17448_ (.A1(_12555_),
    .A2(_10923_),
    .A3(_12876_),
    .B1(_13395_),
    .B2(_13396_),
    .X(_13397_));
 sky130_fd_sc_hd__o311a_2 _17449_ (.A1(\decode.regfile.registers_15[16] ),
    .A2(_12666_),
    .A3(_12773_),
    .B1(_12575_),
    .C1(_13397_),
    .X(_13398_));
 sky130_fd_sc_hd__o221a_2 _17450_ (.A1(\decode.regfile.registers_17[16] ),
    .A2(_12579_),
    .B1(_13379_),
    .B2(_13398_),
    .C1(_12565_),
    .X(_13399_));
 sky130_fd_sc_hd__a211o_2 _17451_ (.A1(\decode.regfile.registers_18[16] ),
    .A2(_12571_),
    .B1(_12561_),
    .C1(_13399_),
    .X(_13400_));
 sky130_fd_sc_hd__o211a_2 _17452_ (.A1(\decode.regfile.registers_19[16] ),
    .A2(_12679_),
    .B1(_12906_),
    .C1(_13400_),
    .X(_13401_));
 sky130_fd_sc_hd__o221a_2 _17453_ (.A1(\decode.regfile.registers_21[16] ),
    .A2(_12716_),
    .B1(_13378_),
    .B2(_13401_),
    .C1(_12806_),
    .X(_13402_));
 sky130_fd_sc_hd__a211o_2 _17454_ (.A1(\decode.regfile.registers_22[16] ),
    .A2(_13100_),
    .B1(_13402_),
    .C1(_13289_),
    .X(_13403_));
 sky130_fd_sc_hd__or4_2 _17455_ (.A(_13081_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[16] ),
    .D(_13041_),
    .X(_13404_));
 sky130_fd_sc_hd__o2111a_2 _17456_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[16] ),
    .B1(_13170_),
    .C1(_13083_),
    .D1(_13367_),
    .X(_13405_));
 sky130_fd_sc_hd__a31o_2 _17457_ (.A1(_13339_),
    .A2(_13403_),
    .A3(_13404_),
    .B1(_13405_),
    .X(_13406_));
 sky130_fd_sc_hd__buf_1 _17458_ (.A(_10595_),
    .X(_13407_));
 sky130_fd_sc_hd__or4_2 _17459_ (.A(_13407_),
    .B(\decode.regfile.registers_25[16] ),
    .C(_13045_),
    .D(_13294_),
    .X(_13408_));
 sky130_fd_sc_hd__o2111a_2 _17460_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[16] ),
    .B1(_13254_),
    .C1(_13047_),
    .D1(_13088_),
    .X(_13409_));
 sky130_fd_sc_hd__a31o_2 _17461_ (.A1(_13183_),
    .A2(_13406_),
    .A3(_13408_),
    .B1(_13409_),
    .X(_13410_));
 sky130_fd_sc_hd__or4_2 _17462_ (.A(_13091_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[16] ),
    .D(_13050_),
    .X(_13411_));
 sky130_fd_sc_hd__o21a_2 _17463_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[16] ),
    .B1(_13093_),
    .X(_13412_));
 sky130_fd_sc_hd__a31o_2 _17464_ (.A1(_13221_),
    .A2(_13410_),
    .A3(_13411_),
    .B1(_13412_),
    .X(_13413_));
 sky130_fd_sc_hd__o221a_2 _17465_ (.A1(_13099_),
    .A2(_13262_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[16] ),
    .C1(_13413_),
    .X(_13414_));
 sky130_fd_sc_hd__o221a_2 _17466_ (.A1(\decode.regfile.registers_31[16] ),
    .A2(_12709_),
    .B1(_13377_),
    .B2(_13414_),
    .C1(_13219_),
    .X(_00436_));
 sky130_fd_sc_hd__o21a_2 _17467_ (.A1(_13055_),
    .A2(\decode.regfile.registers_30[17] ),
    .B1(_13097_),
    .X(_13415_));
 sky130_fd_sc_hd__o2111a_2 _17468_ (.A1(_10926_),
    .A2(\decode.regfile.registers_22[17] ),
    .B1(_12554_),
    .C1(_11009_),
    .D1(_12546_),
    .X(_13416_));
 sky130_fd_sc_hd__a41o_2 _17469_ (.A1(\decode.regfile.registers_20[17] ),
    .A2(_12525_),
    .A3(_12552_),
    .A4(_12523_),
    .B1(_12824_),
    .X(_13417_));
 sky130_fd_sc_hd__o2111a_2 _17470_ (.A1(\decode.regfile.registers_18[17] ),
    .A2(_10924_),
    .B1(_12569_),
    .C1(_11023_),
    .D1(_11008_),
    .X(_13418_));
 sky130_fd_sc_hd__a41o_2 _17471_ (.A1(\decode.regfile.registers_15[17] ),
    .A2(_12555_),
    .A3(_10619_),
    .A4(_12589_),
    .B1(_13031_),
    .X(_13419_));
 sky130_fd_sc_hd__a31o_2 _17472_ (.A1(\decode.regfile.registers_13[17] ),
    .A2(_12927_),
    .A3(_12588_),
    .B1(_12663_),
    .X(_13420_));
 sky130_fd_sc_hd__a32o_2 _17473_ (.A1(\decode.regfile.registers_7[17] ),
    .A2(_12882_),
    .A3(_13020_),
    .B1(_12622_),
    .B2(\decode.regfile.registers_6[17] ),
    .X(_13421_));
 sky130_fd_sc_hd__and3_2 _17474_ (.A(\decode.regfile.registers_1[17] ),
    .B(_12635_),
    .C(_12934_),
    .X(_13422_));
 sky130_fd_sc_hd__a21oi_2 _17475_ (.A1(\decode.regfile.registers_0[17] ),
    .A2(_12778_),
    .B1(_13422_),
    .Y(_13423_));
 sky130_fd_sc_hd__a221oi_2 _17476_ (.A1(\decode.regfile.registers_2[17] ),
    .A2(_12834_),
    .B1(_12639_),
    .B2(\decode.regfile.registers_3[17] ),
    .C1(_12837_),
    .Y(_13424_));
 sky130_fd_sc_hd__o21ai_2 _17477_ (.A1(_12729_),
    .A2(_13423_),
    .B1(_13424_),
    .Y(_13425_));
 sky130_fd_sc_hd__a221o_2 _17478_ (.A1(\decode.regfile.registers_4[17] ),
    .A2(_12548_),
    .B1(_13145_),
    .B2(\decode.regfile.registers_5[17] ),
    .C1(_12625_),
    .X(_13426_));
 sky130_fd_sc_hd__nand2_2 _17479_ (.A(_13425_),
    .B(_13426_),
    .Y(_13427_));
 sky130_fd_sc_hd__nand3b_2 _17480_ (.A_N(_13421_),
    .B(_13427_),
    .C(_12726_),
    .Y(_13428_));
 sky130_fd_sc_hd__o32a_2 _17481_ (.A1(_11017_),
    .A2(_12502_),
    .A3(_12509_),
    .B1(\decode.regfile.registers_8[17] ),
    .B2(_12725_),
    .X(_13429_));
 sky130_fd_sc_hd__a22o_2 _17482_ (.A1(\decode.regfile.registers_9[17] ),
    .A2(_12606_),
    .B1(_13428_),
    .B2(_13429_),
    .X(_13430_));
 sky130_fd_sc_hd__or4b_2 _17483_ (.A(\decode.regfile.registers_10[17] ),
    .B(_10603_),
    .C(_12503_),
    .D_N(_12597_),
    .X(_13431_));
 sky130_fd_sc_hd__o211a_2 _17484_ (.A1(_12599_),
    .A2(_13430_),
    .B1(_13431_),
    .C1(_12791_),
    .X(_13432_));
 sky130_fd_sc_hd__a221o_2 _17485_ (.A1(\decode.regfile.registers_11[17] ),
    .A2(_12724_),
    .B1(_12587_),
    .B2(_12550_),
    .C1(_13432_),
    .X(_13433_));
 sky130_fd_sc_hd__o311a_2 _17486_ (.A1(\decode.regfile.registers_12[17] ),
    .A2(_12542_),
    .A3(_12772_),
    .B1(_12658_),
    .C1(_13433_),
    .X(_13434_));
 sky130_fd_sc_hd__o221a_2 _17487_ (.A1(\decode.regfile.registers_14[17] ),
    .A2(_12984_),
    .B1(_13420_),
    .B2(_13434_),
    .C1(_12874_),
    .X(_13435_));
 sky130_fd_sc_hd__o22ai_2 _17488_ (.A1(\decode.regfile.registers_16[17] ),
    .A2(_13011_),
    .B1(_13419_),
    .B2(_13435_),
    .Y(_13436_));
 sky130_fd_sc_hd__nand2_2 _17489_ (.A(_12719_),
    .B(_13436_),
    .Y(_13437_));
 sky130_fd_sc_hd__o211a_2 _17490_ (.A1(\decode.regfile.registers_17[17] ),
    .A2(_12719_),
    .B1(_12565_),
    .C1(_13437_),
    .X(_13438_));
 sky130_fd_sc_hd__o221a_2 _17491_ (.A1(\decode.regfile.registers_19[17] ),
    .A2(_12678_),
    .B1(_13418_),
    .B2(_13438_),
    .C1(_12906_),
    .X(_13439_));
 sky130_fd_sc_hd__o221a_2 _17492_ (.A1(\decode.regfile.registers_21[17] ),
    .A2(_12716_),
    .B1(_13417_),
    .B2(_13439_),
    .C1(_12909_),
    .X(_13440_));
 sky130_fd_sc_hd__o221a_2 _17493_ (.A1(\decode.regfile.registers_23[17] ),
    .A2(_12714_),
    .B1(_13416_),
    .B2(_13440_),
    .C1(_12515_),
    .X(_13441_));
 sky130_fd_sc_hd__o2111a_2 _17494_ (.A1(_12712_),
    .A2(\decode.regfile.registers_24[17] ),
    .B1(_12997_),
    .C1(_12998_),
    .D1(_11025_),
    .X(_13442_));
 sky130_fd_sc_hd__or2_2 _17495_ (.A(_13441_),
    .B(_13442_),
    .X(_13443_));
 sky130_fd_sc_hd__or4_2 _17496_ (.A(_13407_),
    .B(\decode.regfile.registers_25[17] ),
    .C(_13045_),
    .D(_13294_),
    .X(_13444_));
 sky130_fd_sc_hd__o2111a_2 _17497_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[17] ),
    .B1(_13254_),
    .C1(_13047_),
    .D1(_13088_),
    .X(_13445_));
 sky130_fd_sc_hd__a31o_2 _17498_ (.A1(_13183_),
    .A2(_13443_),
    .A3(_13444_),
    .B1(_13445_),
    .X(_13446_));
 sky130_fd_sc_hd__or4_2 _17499_ (.A(_13091_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[17] ),
    .D(_13050_),
    .X(_13447_));
 sky130_fd_sc_hd__o21a_2 _17500_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[17] ),
    .B1(_13093_),
    .X(_13448_));
 sky130_fd_sc_hd__a31o_2 _17501_ (.A1(_13221_),
    .A2(_13446_),
    .A3(_13447_),
    .B1(_13448_),
    .X(_13449_));
 sky130_fd_sc_hd__o221a_2 _17502_ (.A1(_13099_),
    .A2(_13262_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[17] ),
    .C1(_13449_),
    .X(_13450_));
 sky130_fd_sc_hd__o221a_2 _17503_ (.A1(_12708_),
    .A2(\decode.regfile.registers_31[17] ),
    .B1(_13415_),
    .B2(_13450_),
    .C1(_13219_),
    .X(_00437_));
 sky130_fd_sc_hd__buf_1 _17504_ (.A(_10930_),
    .X(_13451_));
 sky130_fd_sc_hd__o21a_2 _17505_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[18] ),
    .B1(_13097_),
    .X(_13452_));
 sky130_fd_sc_hd__or2_2 _17506_ (.A(_12712_),
    .B(\decode.regfile.registers_24[18] ),
    .X(_13453_));
 sky130_fd_sc_hd__a41o_2 _17507_ (.A1(\decode.regfile.registers_8[18] ),
    .A2(_10593_),
    .A3(_12549_),
    .A4(_12592_),
    .B1(_12606_),
    .X(_13454_));
 sky130_fd_sc_hd__a31o_2 _17508_ (.A1(_12531_),
    .A2(_10592_),
    .A3(_12558_),
    .B1(\decode.regfile.registers_0[18] ),
    .X(_13455_));
 sky130_fd_sc_hd__o221ai_2 _17509_ (.A1(\decode.regfile.registers_1[18] ),
    .A2(_12778_),
    .B1(_12830_),
    .B2(_12882_),
    .C1(_13455_),
    .Y(_13456_));
 sky130_fd_sc_hd__o21ai_2 _17510_ (.A1(\decode.regfile.registers_2[18] ),
    .A2(_10616_),
    .B1(_12729_),
    .Y(_13457_));
 sky130_fd_sc_hd__o21ai_2 _17511_ (.A1(\decode.regfile.registers_3[18] ),
    .A2(_12628_),
    .B1(_12732_),
    .Y(_13458_));
 sky130_fd_sc_hd__a21oi_2 _17512_ (.A1(_13456_),
    .A2(_13457_),
    .B1(_13458_),
    .Y(_13459_));
 sky130_fd_sc_hd__a221o_2 _17513_ (.A1(\decode.regfile.registers_4[18] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[18] ),
    .C1(_12737_),
    .X(_13460_));
 sky130_fd_sc_hd__o22ai_2 _17514_ (.A1(\decode.regfile.registers_6[18] ),
    .A2(_12735_),
    .B1(_13459_),
    .B2(_13460_),
    .Y(_13461_));
 sky130_fd_sc_hd__o21ai_2 _17515_ (.A1(\decode.regfile.registers_7[18] ),
    .A2(_12645_),
    .B1(_12726_),
    .Y(_13462_));
 sky130_fd_sc_hd__a21oi_2 _17516_ (.A1(_12645_),
    .A2(_13461_),
    .B1(_13462_),
    .Y(_13463_));
 sky130_fd_sc_hd__o22ai_2 _17517_ (.A1(\decode.regfile.registers_9[18] ),
    .A2(_12602_),
    .B1(_13454_),
    .B2(_13463_),
    .Y(_13464_));
 sky130_fd_sc_hd__nand2_2 _17518_ (.A(_12790_),
    .B(_13464_),
    .Y(_13465_));
 sky130_fd_sc_hd__o211a_2 _17519_ (.A1(\decode.regfile.registers_10[18] ),
    .A2(_12654_),
    .B1(_12878_),
    .C1(_13465_),
    .X(_13466_));
 sky130_fd_sc_hd__a221o_2 _17520_ (.A1(\decode.regfile.registers_11[18] ),
    .A2(_12595_),
    .B1(_12583_),
    .B2(_12551_),
    .C1(_13466_),
    .X(_13467_));
 sky130_fd_sc_hd__o32a_2 _17521_ (.A1(_11020_),
    .A2(_12490_),
    .A3(_12512_),
    .B1(\decode.regfile.registers_12[18] ),
    .B2(_12591_),
    .X(_13468_));
 sky130_fd_sc_hd__a221o_2 _17522_ (.A1(\decode.regfile.registers_13[18] ),
    .A2(_12775_),
    .B1(_13467_),
    .B2(_13468_),
    .C1(_12664_),
    .X(_13469_));
 sky130_fd_sc_hd__o32a_2 _17523_ (.A1(_11020_),
    .A2(_12491_),
    .A3(_12666_),
    .B1(\decode.regfile.registers_14[18] ),
    .B2(_12670_),
    .X(_13470_));
 sky130_fd_sc_hd__a221o_2 _17524_ (.A1(\decode.regfile.registers_15[18] ),
    .A2(_12585_),
    .B1(_13469_),
    .B2(_13470_),
    .C1(_12673_),
    .X(_13471_));
 sky130_fd_sc_hd__o21a_2 _17525_ (.A1(\decode.regfile.registers_16[18] ),
    .A2(_12576_),
    .B1(_12579_),
    .X(_13472_));
 sky130_fd_sc_hd__a22oi_2 _17526_ (.A1(\decode.regfile.registers_17[18] ),
    .A2(_12901_),
    .B1(_13471_),
    .B2(_13472_),
    .Y(_13473_));
 sky130_fd_sc_hd__a21oi_2 _17527_ (.A1(\decode.regfile.registers_18[18] ),
    .A2(_12571_),
    .B1(_12561_),
    .Y(_13474_));
 sky130_fd_sc_hd__o21ai_2 _17528_ (.A1(_12572_),
    .A2(_13473_),
    .B1(_13474_),
    .Y(_13475_));
 sky130_fd_sc_hd__o41a_2 _17529_ (.A1(\decode.regfile.registers_19[18] ),
    .A2(_10599_),
    .A3(_10589_),
    .A4(_12518_),
    .B1(_12543_),
    .X(_13476_));
 sky130_fd_sc_hd__a221o_2 _17530_ (.A1(\decode.regfile.registers_20[18] ),
    .A2(_12770_),
    .B1(_13475_),
    .B2(_13476_),
    .C1(_12537_),
    .X(_13477_));
 sky130_fd_sc_hd__o211a_2 _17531_ (.A1(_12682_),
    .A2(\decode.regfile.registers_21[18] ),
    .B1(_12806_),
    .C1(_13477_),
    .X(_13478_));
 sky130_fd_sc_hd__a211o_2 _17532_ (.A1(\decode.regfile.registers_22[18] ),
    .A2(_12528_),
    .B1(_13478_),
    .C1(_12687_),
    .X(_13479_));
 sky130_fd_sc_hd__o32a_2 _17533_ (.A1(_10938_),
    .A2(_12542_),
    .A3(_12505_),
    .B1(\decode.regfile.registers_23[18] ),
    .B2(_12714_),
    .X(_13480_));
 sky130_fd_sc_hd__a22o_2 _17534_ (.A1(_12691_),
    .A2(_13453_),
    .B1(_13479_),
    .B2(_13480_),
    .X(_13481_));
 sky130_fd_sc_hd__buf_1 _17535_ (.A(_12505_),
    .X(_13482_));
 sky130_fd_sc_hd__or4_2 _17536_ (.A(_13407_),
    .B(\decode.regfile.registers_25[18] ),
    .C(_13482_),
    .D(_13294_),
    .X(_13483_));
 sky130_fd_sc_hd__buf_1 _17537_ (.A(_11010_),
    .X(_13484_));
 sky130_fd_sc_hd__o2111a_2 _17538_ (.A1(_13087_),
    .A2(\decode.regfile.registers_26[18] ),
    .B1(_13254_),
    .C1(_13484_),
    .D1(_13088_),
    .X(_13485_));
 sky130_fd_sc_hd__a31o_2 _17539_ (.A1(_13183_),
    .A2(_13481_),
    .A3(_13483_),
    .B1(_13485_),
    .X(_13486_));
 sky130_fd_sc_hd__buf_1 _17540_ (.A(_12506_),
    .X(_13487_));
 sky130_fd_sc_hd__or4_2 _17541_ (.A(_13091_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[18] ),
    .D(_13487_),
    .X(_13488_));
 sky130_fd_sc_hd__o21a_2 _17542_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[18] ),
    .B1(_13093_),
    .X(_13489_));
 sky130_fd_sc_hd__a31o_2 _17543_ (.A1(_13221_),
    .A2(_13486_),
    .A3(_13488_),
    .B1(_13489_),
    .X(_13490_));
 sky130_fd_sc_hd__o221a_2 _17544_ (.A1(_13099_),
    .A2(_13262_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[18] ),
    .C1(_13490_),
    .X(_13491_));
 sky130_fd_sc_hd__o221a_2 _17545_ (.A1(\decode.regfile.registers_31[18] ),
    .A2(_12872_),
    .B1(_13452_),
    .B2(_13491_),
    .C1(_13219_),
    .X(_00438_));
 sky130_fd_sc_hd__buf_1 _17546_ (.A(_12486_),
    .X(_13492_));
 sky130_fd_sc_hd__o21a_2 _17547_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[19] ),
    .B1(_13492_),
    .X(_13493_));
 sky130_fd_sc_hd__a31o_2 _17548_ (.A1(\decode.regfile.registers_13[19] ),
    .A2(_12534_),
    .A3(_12589_),
    .B1(_12664_),
    .X(_13494_));
 sky130_fd_sc_hd__a41o_2 _17549_ (.A1(\decode.regfile.registers_9[19] ),
    .A2(_12776_),
    .A3(_12604_),
    .A4(_12532_),
    .B1(_12599_),
    .X(_13495_));
 sky130_fd_sc_hd__a31o_2 _17550_ (.A1(\decode.regfile.registers_2[19] ),
    .A2(_10609_),
    .A3(_12636_),
    .B1(_12639_),
    .X(_13496_));
 sky130_fd_sc_hd__a31o_2 _17551_ (.A1(_12934_),
    .A2(_10592_),
    .A3(_12558_),
    .B1(\decode.regfile.registers_0[19] ),
    .X(_02959_));
 sky130_fd_sc_hd__o221a_2 _17552_ (.A1(\decode.regfile.registers_1[19] ),
    .A2(_12932_),
    .B1(_12830_),
    .B2(_12882_),
    .C1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__o22ai_2 _17553_ (.A1(\decode.regfile.registers_3[19] ),
    .A2(_12629_),
    .B1(_13496_),
    .B2(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__a221oi_2 _17554_ (.A1(\decode.regfile.registers_4[19] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[19] ),
    .C1(_12737_),
    .Y(_02962_));
 sky130_fd_sc_hd__o21ai_2 _17555_ (.A1(_12838_),
    .A2(_02961_),
    .B1(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__o31a_2 _17556_ (.A1(\decode.regfile.registers_6[19] ),
    .A2(_10602_),
    .A3(_12626_),
    .B1(_12645_),
    .X(_02964_));
 sky130_fd_sc_hd__a31o_2 _17557_ (.A1(\decode.regfile.registers_7[19] ),
    .A2(_10617_),
    .A3(_13020_),
    .B1(_12843_),
    .X(_02965_));
 sky130_fd_sc_hd__a21o_2 _17558_ (.A1(_02963_),
    .A2(_02964_),
    .B1(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__o211a_2 _17559_ (.A1(\decode.regfile.registers_8[19] ),
    .A2(_12892_),
    .B1(_12602_),
    .C1(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__o221a_2 _17560_ (.A1(\decode.regfile.registers_10[19] ),
    .A2(_12790_),
    .B1(_13495_),
    .B2(_02967_),
    .C1(_12878_),
    .X(_02968_));
 sky130_fd_sc_hd__a221o_2 _17561_ (.A1(\decode.regfile.registers_11[19] ),
    .A2(_12595_),
    .B1(_12588_),
    .B2(_12551_),
    .C1(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__o311a_2 _17562_ (.A1(\decode.regfile.registers_12[19] ),
    .A2(_12542_),
    .A3(_12723_),
    .B1(_12659_),
    .C1(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__o22ai_2 _17563_ (.A1(\decode.regfile.registers_14[19] ),
    .A2(_12670_),
    .B1(_13494_),
    .B2(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__o21ai_2 _17564_ (.A1(\decode.regfile.registers_15[19] ),
    .A2(_12874_),
    .B1(_12576_),
    .Y(_02972_));
 sky130_fd_sc_hd__a21oi_2 _17565_ (.A1(_12874_),
    .A2(_02971_),
    .B1(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hd__a211o_2 _17566_ (.A1(\decode.regfile.registers_16[19] ),
    .A2(_12674_),
    .B1(_12901_),
    .C1(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__or2_2 _17567_ (.A(\decode.regfile.registers_17[19] ),
    .B(_12580_),
    .X(_02975_));
 sky130_fd_sc_hd__o2111a_2 _17568_ (.A1(\decode.regfile.registers_18[19] ),
    .A2(_10925_),
    .B1(_12569_),
    .C1(_11023_),
    .D1(_11008_),
    .X(_02976_));
 sky130_fd_sc_hd__a31o_2 _17569_ (.A1(_12566_),
    .A2(_02974_),
    .A3(_02975_),
    .B1(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__o41a_2 _17570_ (.A1(\decode.regfile.registers_19[19] ),
    .A2(_11013_),
    .A3(_10589_),
    .A4(_12519_),
    .B1(_12544_),
    .X(_02978_));
 sky130_fd_sc_hd__a221o_2 _17571_ (.A1(\decode.regfile.registers_20[19] ),
    .A2(_12771_),
    .B1(_02977_),
    .B2(_02978_),
    .C1(_12538_),
    .X(_02979_));
 sky130_fd_sc_hd__o21a_2 _17572_ (.A1(\decode.regfile.registers_21[19] ),
    .A2(_12682_),
    .B1(_12909_),
    .X(_02980_));
 sky130_fd_sc_hd__a221o_2 _17573_ (.A1(\decode.regfile.registers_22[19] ),
    .A2(_12527_),
    .B1(_02979_),
    .B2(_02980_),
    .C1(_12686_),
    .X(_02981_));
 sky130_fd_sc_hd__or4_2 _17574_ (.A(_13081_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[19] ),
    .D(_13041_),
    .X(_02982_));
 sky130_fd_sc_hd__o2111a_2 _17575_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[19] ),
    .B1(_13170_),
    .C1(_13083_),
    .D1(_13367_),
    .X(_02983_));
 sky130_fd_sc_hd__a31o_2 _17576_ (.A1(_13339_),
    .A2(_02981_),
    .A3(_02982_),
    .B1(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__or4_2 _17577_ (.A(_13407_),
    .B(\decode.regfile.registers_25[19] ),
    .C(_13482_),
    .D(_13294_),
    .X(_02985_));
 sky130_fd_sc_hd__buf_1 _17578_ (.A(_12494_),
    .X(_02986_));
 sky130_fd_sc_hd__buf_1 _17579_ (.A(_11026_),
    .X(_02987_));
 sky130_fd_sc_hd__o2111a_2 _17580_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[19] ),
    .B1(_13254_),
    .C1(_13484_),
    .D1(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__a31o_2 _17581_ (.A1(_13183_),
    .A2(_02984_),
    .A3(_02985_),
    .B1(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__buf_1 _17582_ (.A(_10939_),
    .X(_02990_));
 sky130_fd_sc_hd__or4_2 _17583_ (.A(_02990_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[19] ),
    .D(_13487_),
    .X(_02991_));
 sky130_fd_sc_hd__buf_1 _17584_ (.A(_12697_),
    .X(_02992_));
 sky130_fd_sc_hd__o21a_2 _17585_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[19] ),
    .B1(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__a31o_2 _17586_ (.A1(_13221_),
    .A2(_02989_),
    .A3(_02991_),
    .B1(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__o221a_2 _17587_ (.A1(_13099_),
    .A2(_13262_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[19] ),
    .C1(_02994_),
    .X(_02995_));
 sky130_fd_sc_hd__o221a_2 _17588_ (.A1(\decode.regfile.registers_31[19] ),
    .A2(_12872_),
    .B1(_13493_),
    .B2(_02995_),
    .C1(_13219_),
    .X(_00439_));
 sky130_fd_sc_hd__o21a_2 _17589_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[20] ),
    .B1(_13492_),
    .X(_02996_));
 sky130_fd_sc_hd__buf_1 _17590_ (.A(_10930_),
    .X(_02997_));
 sky130_fd_sc_hd__o2111a_2 _17591_ (.A1(\decode.regfile.registers_18[20] ),
    .A2(_10924_),
    .B1(_12568_),
    .C1(_12524_),
    .D1(_10612_),
    .X(_02998_));
 sky130_fd_sc_hd__a41o_2 _17592_ (.A1(\decode.regfile.registers_15[20] ),
    .A2(_12555_),
    .A3(_10923_),
    .A4(_12876_),
    .B1(_13031_),
    .X(_02999_));
 sky130_fd_sc_hd__a31o_2 _17593_ (.A1(\decode.regfile.registers_13[20] ),
    .A2(_12927_),
    .A3(_12583_),
    .B1(_12663_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_2 _17594_ (.A0(\decode.regfile.registers_1[20] ),
    .A1(\decode.regfile.registers_0[20] ),
    .S(_12631_),
    .X(_03001_));
 sky130_fd_sc_hd__a221oi_2 _17595_ (.A1(\decode.regfile.registers_2[20] ),
    .A2(_12834_),
    .B1(_12639_),
    .B2(\decode.regfile.registers_3[20] ),
    .C1(_12838_),
    .Y(_03002_));
 sky130_fd_sc_hd__a21bo_2 _17596_ (.A1(_12830_),
    .A2(_03001_),
    .B1_N(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__a221o_2 _17597_ (.A1(\decode.regfile.registers_4[20] ),
    .A2(_12548_),
    .B1(_13145_),
    .B2(\decode.regfile.registers_5[20] ),
    .C1(_12614_),
    .X(_03004_));
 sky130_fd_sc_hd__nand2_2 _17598_ (.A(_03003_),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__a221oi_2 _17599_ (.A1(\decode.regfile.registers_7[20] ),
    .A2(_12610_),
    .B1(_12623_),
    .B2(\decode.regfile.registers_6[20] ),
    .C1(_12843_),
    .Y(_03006_));
 sky130_fd_sc_hd__nand2_2 _17600_ (.A(_03005_),
    .B(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__o32a_2 _17601_ (.A1(_11017_),
    .A2(_12502_),
    .A3(_12509_),
    .B1(\decode.regfile.registers_8[20] ),
    .B2(_12725_),
    .X(_03008_));
 sky130_fd_sc_hd__a22oi_2 _17602_ (.A1(\decode.regfile.registers_9[20] ),
    .A2(_12606_),
    .B1(_03007_),
    .B2(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__nand2_2 _17603_ (.A(_03009_),
    .B(_12653_),
    .Y(_03010_));
 sky130_fd_sc_hd__o21a_2 _17604_ (.A1(\decode.regfile.registers_10[20] ),
    .A2(_12652_),
    .B1(_12791_),
    .X(_03011_));
 sky130_fd_sc_hd__a221o_2 _17605_ (.A1(\decode.regfile.registers_11[20] ),
    .A2(_12594_),
    .B1(_03010_),
    .B2(_03011_),
    .C1(_12794_),
    .X(_03012_));
 sky130_fd_sc_hd__o311a_2 _17606_ (.A1(\decode.regfile.registers_12[20] ),
    .A2(_12541_),
    .A3(_12772_),
    .B1(_12658_),
    .C1(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__o221a_2 _17607_ (.A1(\decode.regfile.registers_14[20] ),
    .A2(_12984_),
    .B1(_03000_),
    .B2(_03013_),
    .C1(_12874_),
    .X(_03014_));
 sky130_fd_sc_hd__o22a_2 _17608_ (.A1(\decode.regfile.registers_16[20] ),
    .A2(_12575_),
    .B1(_02999_),
    .B2(_03014_),
    .X(_03015_));
 sky130_fd_sc_hd__o21a_2 _17609_ (.A1(\decode.regfile.registers_17[20] ),
    .A2(_12578_),
    .B1(_12564_),
    .X(_03016_));
 sky130_fd_sc_hd__o21a_2 _17610_ (.A1(_12901_),
    .A2(_03015_),
    .B1(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__o221a_2 _17611_ (.A1(\decode.regfile.registers_19[20] ),
    .A2(_12678_),
    .B1(_02998_),
    .B2(_03017_),
    .C1(_12544_),
    .X(_03018_));
 sky130_fd_sc_hd__a211o_2 _17612_ (.A1(\decode.regfile.registers_20[20] ),
    .A2(_12771_),
    .B1(_03018_),
    .C1(_12537_),
    .X(_03019_));
 sky130_fd_sc_hd__o211a_2 _17613_ (.A1(_12822_),
    .A2(\decode.regfile.registers_21[20] ),
    .B1(_13164_),
    .C1(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__a211o_2 _17614_ (.A1(\decode.regfile.registers_22[20] ),
    .A2(_13100_),
    .B1(_03020_),
    .C1(_13289_),
    .X(_03021_));
 sky130_fd_sc_hd__or4_2 _17615_ (.A(_13081_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[20] ),
    .D(_13041_),
    .X(_03022_));
 sky130_fd_sc_hd__o2111a_2 _17616_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[20] ),
    .B1(_13170_),
    .C1(_13083_),
    .D1(_13367_),
    .X(_03023_));
 sky130_fd_sc_hd__a31o_2 _17617_ (.A1(_13339_),
    .A2(_03021_),
    .A3(_03022_),
    .B1(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__or4_2 _17618_ (.A(_13407_),
    .B(\decode.regfile.registers_25[20] ),
    .C(_13482_),
    .D(_13294_),
    .X(_03025_));
 sky130_fd_sc_hd__o2111a_2 _17619_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[20] ),
    .B1(_13254_),
    .C1(_13484_),
    .D1(_02987_),
    .X(_03026_));
 sky130_fd_sc_hd__a31o_2 _17620_ (.A1(_13183_),
    .A2(_03024_),
    .A3(_03025_),
    .B1(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__or4_2 _17621_ (.A(_02990_),
    .B(_13176_),
    .C(\decode.regfile.registers_27[20] ),
    .D(_13487_),
    .X(_03028_));
 sky130_fd_sc_hd__o21a_2 _17622_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[20] ),
    .B1(_02992_),
    .X(_03029_));
 sky130_fd_sc_hd__a31o_2 _17623_ (.A1(_13221_),
    .A2(_03027_),
    .A3(_03028_),
    .B1(_03029_),
    .X(_03030_));
 sky130_fd_sc_hd__o221a_2 _17624_ (.A1(_02997_),
    .A2(_13262_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[20] ),
    .C1(_03030_),
    .X(_03031_));
 sky130_fd_sc_hd__o221a_2 _17625_ (.A1(\decode.regfile.registers_31[20] ),
    .A2(_12872_),
    .B1(_02996_),
    .B2(_03031_),
    .C1(_13219_),
    .X(_00440_));
 sky130_fd_sc_hd__o21a_2 _17626_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[21] ),
    .B1(_13492_),
    .X(_03032_));
 sky130_fd_sc_hd__a41o_2 _17627_ (.A1(\decode.regfile.registers_15[21] ),
    .A2(_10612_),
    .A3(_10619_),
    .A4(_12589_),
    .B1(_13031_),
    .X(_03033_));
 sky130_fd_sc_hd__a41o_2 _17628_ (.A1(\decode.regfile.registers_9[21] ),
    .A2(_10594_),
    .A3(_12690_),
    .A4(_12533_),
    .B1(_12599_),
    .X(_03034_));
 sky130_fd_sc_hd__o2bb2ai_2 _17629_ (.A1_N(\decode.regfile.registers_0[21] ),
    .A2_N(_12631_),
    .B1(_12508_),
    .B2(_12933_),
    .Y(_03035_));
 sky130_fd_sc_hd__a31o_2 _17630_ (.A1(\decode.regfile.registers_1[21] ),
    .A2(_12636_),
    .A3(_13145_),
    .B1(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__o211ai_2 _17631_ (.A1(\decode.regfile.registers_2[21] ),
    .A2(_12634_),
    .B1(_12629_),
    .C1(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__nand2_2 _17632_ (.A(\decode.regfile.registers_3[21] ),
    .B(_12836_),
    .Y(_03038_));
 sky130_fd_sc_hd__mux2_2 _17633_ (.A0(\decode.regfile.registers_4[21] ),
    .A1(\decode.regfile.registers_5[21] ),
    .S(_12508_),
    .X(_03039_));
 sky130_fd_sc_hd__and4b_2 _17634_ (.A_N(_03039_),
    .B(_10602_),
    .C(_10593_),
    .D(_12522_),
    .X(_03040_));
 sky130_fd_sc_hd__a31o_2 _17635_ (.A1(_12732_),
    .A2(_03037_),
    .A3(_03038_),
    .B1(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__nand2_2 _17636_ (.A(_12880_),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__o221ai_2 _17637_ (.A1(_12649_),
    .A2(_12615_),
    .B1(_12880_),
    .B2(\decode.regfile.registers_6[21] ),
    .C1(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__a21oi_2 _17638_ (.A1(\decode.regfile.registers_7[21] ),
    .A2(_12612_),
    .B1(_12889_),
    .Y(_03044_));
 sky130_fd_sc_hd__o21ai_2 _17639_ (.A1(\decode.regfile.registers_8[21] ),
    .A2(_12892_),
    .B1(_12603_),
    .Y(_03045_));
 sky130_fd_sc_hd__a21oi_2 _17640_ (.A1(_03043_),
    .A2(_03044_),
    .B1(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__o221ai_2 _17641_ (.A1(\decode.regfile.registers_10[21] ),
    .A2(_12654_),
    .B1(_03034_),
    .B2(_03046_),
    .C1(_12878_),
    .Y(_03047_));
 sky130_fd_sc_hd__o2bb2a_2 _17642_ (.A1_N(\decode.regfile.registers_11[21] ),
    .A2_N(_12724_),
    .B1(_12722_),
    .B2(_12540_),
    .X(_03048_));
 sky130_fd_sc_hd__nand2_2 _17643_ (.A(_03047_),
    .B(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__or4_2 _17644_ (.A(\decode.regfile.registers_12[21] ),
    .B(_12489_),
    .C(_11019_),
    .D(_12541_),
    .X(_03050_));
 sky130_fd_sc_hd__a31o_2 _17645_ (.A1(\decode.regfile.registers_13[21] ),
    .A2(_12927_),
    .A3(_12587_),
    .B1(_12662_),
    .X(_03051_));
 sky130_fd_sc_hd__a31o_2 _17646_ (.A1(_12659_),
    .A2(_03049_),
    .A3(_03050_),
    .B1(_03051_),
    .X(_03052_));
 sky130_fd_sc_hd__o221a_2 _17647_ (.A1(_12666_),
    .A2(_12773_),
    .B1(_12984_),
    .B2(\decode.regfile.registers_14[21] ),
    .C1(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__o22a_2 _17648_ (.A1(\decode.regfile.registers_16[21] ),
    .A2(_13011_),
    .B1(_03033_),
    .B2(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__or2_2 _17649_ (.A(\decode.regfile.registers_17[21] ),
    .B(_12579_),
    .X(_03055_));
 sky130_fd_sc_hd__o211a_2 _17650_ (.A1(_12901_),
    .A2(_03054_),
    .B1(_03055_),
    .C1(_12826_),
    .X(_03056_));
 sky130_fd_sc_hd__a211o_2 _17651_ (.A1(\decode.regfile.registers_18[21] ),
    .A2(_12572_),
    .B1(_12562_),
    .C1(_03056_),
    .X(_03057_));
 sky130_fd_sc_hd__o41a_2 _17652_ (.A1(\decode.regfile.registers_19[21] ),
    .A2(_11013_),
    .A3(_10589_),
    .A4(_12519_),
    .B1(_12544_),
    .X(_03058_));
 sky130_fd_sc_hd__a221o_2 _17653_ (.A1(\decode.regfile.registers_20[21] ),
    .A2(_12771_),
    .B1(_03057_),
    .B2(_03058_),
    .C1(_12538_),
    .X(_03059_));
 sky130_fd_sc_hd__o21a_2 _17654_ (.A1(\decode.regfile.registers_21[21] ),
    .A2(_12822_),
    .B1(_12909_),
    .X(_03060_));
 sky130_fd_sc_hd__a221o_2 _17655_ (.A1(\decode.regfile.registers_22[21] ),
    .A2(_12527_),
    .B1(_03059_),
    .B2(_03060_),
    .C1(_12686_),
    .X(_03061_));
 sky130_fd_sc_hd__or4_2 _17656_ (.A(_13081_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[21] ),
    .D(_12995_),
    .X(_03062_));
 sky130_fd_sc_hd__o2111a_2 _17657_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[21] ),
    .B1(_13170_),
    .C1(_13083_),
    .D1(_13367_),
    .X(_03063_));
 sky130_fd_sc_hd__a31o_2 _17658_ (.A1(_13339_),
    .A2(_03061_),
    .A3(_03062_),
    .B1(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__or4_2 _17659_ (.A(_13407_),
    .B(\decode.regfile.registers_25[21] ),
    .C(_13482_),
    .D(_13294_),
    .X(_03065_));
 sky130_fd_sc_hd__o2111a_2 _17660_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[21] ),
    .B1(_13254_),
    .C1(_13484_),
    .D1(_02987_),
    .X(_03066_));
 sky130_fd_sc_hd__a31o_2 _17661_ (.A1(_13183_),
    .A2(_03064_),
    .A3(_03065_),
    .B1(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__buf_1 _17662_ (.A(_12667_),
    .X(_03068_));
 sky130_fd_sc_hd__or4_2 _17663_ (.A(_02990_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[21] ),
    .D(_13487_),
    .X(_03069_));
 sky130_fd_sc_hd__o21a_2 _17664_ (.A1(_13215_),
    .A2(\decode.regfile.registers_28[21] ),
    .B1(_02992_),
    .X(_03070_));
 sky130_fd_sc_hd__a31o_2 _17665_ (.A1(_13221_),
    .A2(_03067_),
    .A3(_03069_),
    .B1(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__o221a_2 _17666_ (.A1(_02997_),
    .A2(_13262_),
    .B1(_13182_),
    .B2(\decode.regfile.registers_29[21] ),
    .C1(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__buf_1 _17667_ (.A(_12704_),
    .X(_03073_));
 sky130_fd_sc_hd__o221a_2 _17668_ (.A1(\decode.regfile.registers_31[21] ),
    .A2(_12872_),
    .B1(_03032_),
    .B2(_03072_),
    .C1(_03073_),
    .X(_00441_));
 sky130_fd_sc_hd__o21a_2 _17669_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[22] ),
    .B1(_13492_),
    .X(_03074_));
 sky130_fd_sc_hd__a21o_2 _17670_ (.A1(\decode.regfile.registers_18[22] ),
    .A2(_12571_),
    .B1(_12561_),
    .X(_03075_));
 sky130_fd_sc_hd__and4_2 _17671_ (.A(\decode.regfile.registers_17[22] ),
    .B(_11021_),
    .C(_12559_),
    .D(_12534_),
    .X(_03076_));
 sky130_fd_sc_hd__a41o_2 _17672_ (.A1(\decode.regfile.registers_15[22] ),
    .A2(_10611_),
    .A3(_10923_),
    .A4(_12876_),
    .B1(_12672_),
    .X(_03077_));
 sky130_fd_sc_hd__a21oi_2 _17673_ (.A1(_12636_),
    .A2(_13145_),
    .B1(\decode.regfile.registers_0[22] ),
    .Y(_03078_));
 sky130_fd_sc_hd__a31o_2 _17674_ (.A1(_12138_),
    .A2(_12636_),
    .A3(_12531_),
    .B1(_12728_),
    .X(_03079_));
 sky130_fd_sc_hd__a221oi_2 _17675_ (.A1(\decode.regfile.registers_2[22] ),
    .A2(_12835_),
    .B1(_12639_),
    .B2(\decode.regfile.registers_3[22] ),
    .C1(_12838_),
    .Y(_03080_));
 sky130_fd_sc_hd__o21ai_2 _17676_ (.A1(_03078_),
    .A2(_03079_),
    .B1(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__a221o_2 _17677_ (.A1(\decode.regfile.registers_4[22] ),
    .A2(_12548_),
    .B1(_13145_),
    .B2(\decode.regfile.registers_5[22] ),
    .C1(_12625_),
    .X(_03082_));
 sky130_fd_sc_hd__a32o_2 _17678_ (.A1(\decode.regfile.registers_7[22] ),
    .A2(_12882_),
    .A3(_13020_),
    .B1(_12622_),
    .B2(\decode.regfile.registers_6[22] ),
    .X(_03083_));
 sky130_fd_sc_hd__a21oi_2 _17679_ (.A1(_03081_),
    .A2(_03082_),
    .B1(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__a21oi_2 _17680_ (.A1(\decode.regfile.registers_8[22] ),
    .A2(_12843_),
    .B1(_12606_),
    .Y(_03085_));
 sky130_fd_sc_hd__o21ai_2 _17681_ (.A1(_12888_),
    .A2(_03084_),
    .B1(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__o41a_2 _17682_ (.A1(\decode.regfile.registers_9[22] ),
    .A2(_11017_),
    .A3(_12502_),
    .A4(_12509_),
    .B1(_12652_),
    .X(_03087_));
 sky130_fd_sc_hd__a22o_2 _17683_ (.A1(\decode.regfile.registers_10[22] ),
    .A2(_12598_),
    .B1(_03086_),
    .B2(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__a22o_2 _17684_ (.A1(\decode.regfile.registers_11[22] ),
    .A2(_12594_),
    .B1(_12582_),
    .B2(_12550_),
    .X(_03089_));
 sky130_fd_sc_hd__a21o_2 _17685_ (.A1(_12792_),
    .A2(_03088_),
    .B1(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__o32a_2 _17686_ (.A1(_12498_),
    .A2(_12489_),
    .A3(_12510_),
    .B1(\decode.regfile.registers_12[22] ),
    .B2(_12590_),
    .X(_03091_));
 sky130_fd_sc_hd__a221o_2 _17687_ (.A1(\decode.regfile.registers_13[22] ),
    .A2(_12774_),
    .B1(_03090_),
    .B2(_03091_),
    .C1(_12662_),
    .X(_03092_));
 sky130_fd_sc_hd__o221a_2 _17688_ (.A1(_12650_),
    .A2(_12723_),
    .B1(_12669_),
    .B2(\decode.regfile.registers_14[22] ),
    .C1(_03092_),
    .X(_03093_));
 sky130_fd_sc_hd__o221a_2 _17689_ (.A1(\decode.regfile.registers_16[22] ),
    .A2(_12575_),
    .B1(_03077_),
    .B2(_03093_),
    .C1(_12578_),
    .X(_03094_));
 sky130_fd_sc_hd__o21a_2 _17690_ (.A1(_03076_),
    .A2(_03094_),
    .B1(_12565_),
    .X(_03095_));
 sky130_fd_sc_hd__o221a_2 _17691_ (.A1(\decode.regfile.registers_19[22] ),
    .A2(_12678_),
    .B1(_03075_),
    .B2(_03095_),
    .C1(_12544_),
    .X(_03096_));
 sky130_fd_sc_hd__a211o_2 _17692_ (.A1(\decode.regfile.registers_20[22] ),
    .A2(_12771_),
    .B1(_03096_),
    .C1(_12537_),
    .X(_03097_));
 sky130_fd_sc_hd__o211a_2 _17693_ (.A1(_12822_),
    .A2(\decode.regfile.registers_21[22] ),
    .B1(_13164_),
    .C1(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__a211o_2 _17694_ (.A1(\decode.regfile.registers_22[22] ),
    .A2(_13100_),
    .B1(_03098_),
    .C1(_13289_),
    .X(_03099_));
 sky130_fd_sc_hd__or4_2 _17695_ (.A(_11014_),
    .B(_13168_),
    .C(\decode.regfile.registers_23[22] ),
    .D(_12995_),
    .X(_03100_));
 sky130_fd_sc_hd__o2111a_2 _17696_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[22] ),
    .B1(_13170_),
    .C1(_12998_),
    .D1(_13367_),
    .X(_03101_));
 sky130_fd_sc_hd__a31o_2 _17697_ (.A1(_13339_),
    .A2(_03099_),
    .A3(_03100_),
    .B1(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__or4_2 _17698_ (.A(_13407_),
    .B(\decode.regfile.registers_25[22] ),
    .C(_13482_),
    .D(_13294_),
    .X(_03103_));
 sky130_fd_sc_hd__o2111a_2 _17699_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[22] ),
    .B1(_13254_),
    .C1(_13484_),
    .D1(_02987_),
    .X(_03104_));
 sky130_fd_sc_hd__a31o_2 _17700_ (.A1(_12968_),
    .A2(_03102_),
    .A3(_03103_),
    .B1(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__or4_2 _17701_ (.A(_02990_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[22] ),
    .D(_13487_),
    .X(_03106_));
 sky130_fd_sc_hd__o21a_2 _17702_ (.A1(_10929_),
    .A2(\decode.regfile.registers_28[22] ),
    .B1(_02992_),
    .X(_03107_));
 sky130_fd_sc_hd__a31o_2 _17703_ (.A1(_13221_),
    .A2(_03105_),
    .A3(_03106_),
    .B1(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__o221a_2 _17704_ (.A1(_02997_),
    .A2(_13262_),
    .B1(_12965_),
    .B2(\decode.regfile.registers_29[22] ),
    .C1(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__o221a_2 _17705_ (.A1(_12708_),
    .A2(\decode.regfile.registers_31[22] ),
    .B1(_03074_),
    .B2(_03109_),
    .C1(_03073_),
    .X(_00442_));
 sky130_fd_sc_hd__o21a_2 _17706_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[23] ),
    .B1(_13492_),
    .X(_03110_));
 sky130_fd_sc_hd__a41o_2 _17707_ (.A1(\decode.regfile.registers_20[23] ),
    .A2(_12525_),
    .A3(_12552_),
    .A4(_12823_),
    .B1(_12824_),
    .X(_03111_));
 sky130_fd_sc_hd__o2111a_2 _17708_ (.A1(\decode.regfile.registers_18[23] ),
    .A2(_10925_),
    .B1(_12569_),
    .C1(_11023_),
    .D1(_11008_),
    .X(_03112_));
 sky130_fd_sc_hd__and4_2 _17709_ (.A(\decode.regfile.registers_17[23] ),
    .B(_11022_),
    .C(_12567_),
    .D(_12586_),
    .X(_03113_));
 sky130_fd_sc_hd__a41o_2 _17710_ (.A1(\decode.regfile.registers_15[23] ),
    .A2(_10612_),
    .A3(_10619_),
    .A4(_12589_),
    .B1(_13031_),
    .X(_03114_));
 sky130_fd_sc_hd__a31o_2 _17711_ (.A1(\decode.regfile.registers_13[23] ),
    .A2(_12927_),
    .A3(_12588_),
    .B1(_12663_),
    .X(_03115_));
 sky130_fd_sc_hd__o21ai_2 _17712_ (.A1(\decode.regfile.registers_10[23] ),
    .A2(_12790_),
    .B1(_12878_),
    .Y(_03116_));
 sky130_fd_sc_hd__mux2_2 _17713_ (.A0(\decode.regfile.registers_4[23] ),
    .A1(\decode.regfile.registers_5[23] ),
    .S(_12882_),
    .X(_03117_));
 sky130_fd_sc_hd__a31o_2 _17714_ (.A1(\decode.regfile.registers_3[23] ),
    .A2(_10616_),
    .A3(_12729_),
    .B1(_12838_),
    .X(_03118_));
 sky130_fd_sc_hd__and3_2 _17715_ (.A(\decode.regfile.registers_1[23] ),
    .B(_12635_),
    .C(_12530_),
    .X(_03119_));
 sky130_fd_sc_hd__a211o_2 _17716_ (.A1(\decode.regfile.registers_0[23] ),
    .A2(_12932_),
    .B1(_12834_),
    .C1(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__o211a_2 _17717_ (.A1(\decode.regfile.registers_2[23] ),
    .A2(_12634_),
    .B1(_12628_),
    .C1(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__o32a_2 _17718_ (.A1(_10610_),
    .A2(_12626_),
    .A3(_03117_),
    .B1(_03118_),
    .B2(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__o22ai_2 _17719_ (.A1(\decode.regfile.registers_6[23] ),
    .A2(_12735_),
    .B1(_12623_),
    .B2(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__a21oi_2 _17720_ (.A1(\decode.regfile.registers_7[23] ),
    .A2(_12612_),
    .B1(_12889_),
    .Y(_03124_));
 sky130_fd_sc_hd__o21ai_2 _17721_ (.A1(_12612_),
    .A2(_03123_),
    .B1(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__o32a_2 _17722_ (.A1(_11018_),
    .A2(_12977_),
    .A3(_12510_),
    .B1(\decode.regfile.registers_8[23] ),
    .B2(_12892_),
    .X(_03126_));
 sky130_fd_sc_hd__a221oi_2 _17723_ (.A1(\decode.regfile.registers_9[23] ),
    .A2(_12607_),
    .B1(_03125_),
    .B2(_03126_),
    .C1(_12600_),
    .Y(_03127_));
 sky130_fd_sc_hd__or4b_2 _17724_ (.A(_12498_),
    .B(_12504_),
    .C(_12649_),
    .D_N(\decode.regfile.registers_11[23] ),
    .X(_03128_));
 sky130_fd_sc_hd__o211ai_2 _17725_ (.A1(_03116_),
    .A2(_03127_),
    .B1(_12591_),
    .C1(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__o311a_2 _17726_ (.A1(\decode.regfile.registers_12[23] ),
    .A2(_12542_),
    .A3(_12772_),
    .B1(_12658_),
    .C1(_03129_),
    .X(_03130_));
 sky130_fd_sc_hd__o221a_2 _17727_ (.A1(\decode.regfile.registers_14[23] ),
    .A2(_12984_),
    .B1(_03115_),
    .B2(_03130_),
    .C1(_12874_),
    .X(_03131_));
 sky130_fd_sc_hd__o221a_2 _17728_ (.A1(\decode.regfile.registers_16[23] ),
    .A2(_13011_),
    .B1(_03114_),
    .B2(_03131_),
    .C1(_12579_),
    .X(_03132_));
 sky130_fd_sc_hd__o21a_2 _17729_ (.A1(_03113_),
    .A2(_03132_),
    .B1(_12566_),
    .X(_03133_));
 sky130_fd_sc_hd__o221a_2 _17730_ (.A1(\decode.regfile.registers_19[23] ),
    .A2(_12678_),
    .B1(_03112_),
    .B2(_03133_),
    .C1(_12906_),
    .X(_03134_));
 sky130_fd_sc_hd__o221a_2 _17731_ (.A1(\decode.regfile.registers_21[23] ),
    .A2(_12716_),
    .B1(_03111_),
    .B2(_03134_),
    .C1(_13164_),
    .X(_03135_));
 sky130_fd_sc_hd__a211o_2 _17732_ (.A1(\decode.regfile.registers_22[23] ),
    .A2(_13100_),
    .B1(_03135_),
    .C1(_13289_),
    .X(_03136_));
 sky130_fd_sc_hd__or4_2 _17733_ (.A(_11014_),
    .B(_10936_),
    .C(\decode.regfile.registers_23[23] ),
    .D(_12995_),
    .X(_03137_));
 sky130_fd_sc_hd__o2111a_2 _17734_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[23] ),
    .B1(_12997_),
    .C1(_12998_),
    .D1(_13367_),
    .X(_03138_));
 sky130_fd_sc_hd__a31o_2 _17735_ (.A1(_13339_),
    .A2(_03136_),
    .A3(_03137_),
    .B1(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__or4_2 _17736_ (.A(_13407_),
    .B(\decode.regfile.registers_25[23] ),
    .C(_13482_),
    .D(_13294_),
    .X(_03140_));
 sky130_fd_sc_hd__o2111a_2 _17737_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[23] ),
    .B1(_13002_),
    .C1(_13484_),
    .D1(_02987_),
    .X(_03141_));
 sky130_fd_sc_hd__a31o_2 _17738_ (.A1(_12968_),
    .A2(_03139_),
    .A3(_03140_),
    .B1(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__or4_2 _17739_ (.A(_02990_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[23] ),
    .D(_13487_),
    .X(_03143_));
 sky130_fd_sc_hd__o21a_2 _17740_ (.A1(_10929_),
    .A2(\decode.regfile.registers_28[23] ),
    .B1(_02992_),
    .X(_03144_));
 sky130_fd_sc_hd__a31o_2 _17741_ (.A1(_12967_),
    .A2(_03142_),
    .A3(_03143_),
    .B1(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__o221a_2 _17742_ (.A1(_02997_),
    .A2(_13262_),
    .B1(_12965_),
    .B2(\decode.regfile.registers_29[23] ),
    .C1(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__o221a_2 _17743_ (.A1(_12708_),
    .A2(\decode.regfile.registers_31[23] ),
    .B1(_03110_),
    .B2(_03146_),
    .C1(_03073_),
    .X(_00443_));
 sky130_fd_sc_hd__o21a_2 _17744_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[24] ),
    .B1(_13492_),
    .X(_03147_));
 sky130_fd_sc_hd__a41o_2 _17745_ (.A1(\decode.regfile.registers_20[24] ),
    .A2(_12525_),
    .A3(_12552_),
    .A4(_12823_),
    .B1(_12824_),
    .X(_03148_));
 sky130_fd_sc_hd__o21ai_2 _17746_ (.A1(\decode.regfile.registers_19[24] ),
    .A2(_12679_),
    .B1(_12906_),
    .Y(_03149_));
 sky130_fd_sc_hd__a32o_2 _17747_ (.A1(_11022_),
    .A2(_12568_),
    .A3(_12535_),
    .B1(_12674_),
    .B2(\decode.regfile.registers_16[24] ),
    .X(_03150_));
 sky130_fd_sc_hd__a31o_2 _17748_ (.A1(\decode.regfile.registers_13[24] ),
    .A2(_12534_),
    .A3(_12876_),
    .B1(_12664_),
    .X(_03151_));
 sky130_fd_sc_hd__a221o_2 _17749_ (.A1(\decode.regfile.registers_7[24] ),
    .A2(_12611_),
    .B1(_12623_),
    .B2(\decode.regfile.registers_6[24] ),
    .C1(_12888_),
    .X(_03152_));
 sky130_fd_sc_hd__a31o_2 _17750_ (.A1(\decode.regfile.registers_3[24] ),
    .A2(_10616_),
    .A3(_12729_),
    .B1(_12838_),
    .X(_03153_));
 sky130_fd_sc_hd__and3_2 _17751_ (.A(\decode.regfile.registers_1[24] ),
    .B(_12635_),
    .C(_12530_),
    .X(_03154_));
 sky130_fd_sc_hd__a211o_2 _17752_ (.A1(\decode.regfile.registers_0[24] ),
    .A2(_12932_),
    .B1(_12834_),
    .C1(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__o211a_2 _17753_ (.A1(\decode.regfile.registers_2[24] ),
    .A2(_12634_),
    .B1(_12628_),
    .C1(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__o31a_2 _17754_ (.A1(\decode.regfile.registers_5[24] ),
    .A2(_12509_),
    .A3(_12614_),
    .B1(_12735_),
    .X(_03157_));
 sky130_fd_sc_hd__or4_2 _17755_ (.A(\decode.regfile.registers_4[24] ),
    .B(_10609_),
    .C(_12882_),
    .D(_12614_),
    .X(_03158_));
 sky130_fd_sc_hd__o211a_2 _17756_ (.A1(_03153_),
    .A2(_03156_),
    .B1(_03157_),
    .C1(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__o22a_2 _17757_ (.A1(\decode.regfile.registers_8[24] ),
    .A2(_12726_),
    .B1(_03152_),
    .B2(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__and4_2 _17758_ (.A(\decode.regfile.registers_9[24] ),
    .B(_12604_),
    .C(_12532_),
    .D(_12776_),
    .X(_03161_));
 sky130_fd_sc_hd__a211o_2 _17759_ (.A1(_03160_),
    .A2(_12603_),
    .B1(_12600_),
    .C1(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__o21a_2 _17760_ (.A1(\decode.regfile.registers_10[24] ),
    .A2(_12790_),
    .B1(_12792_),
    .X(_03163_));
 sky130_fd_sc_hd__a221o_2 _17761_ (.A1(\decode.regfile.registers_11[24] ),
    .A2(_12595_),
    .B1(_03162_),
    .B2(_03163_),
    .C1(_12794_),
    .X(_03164_));
 sky130_fd_sc_hd__o311a_2 _17762_ (.A1(\decode.regfile.registers_12[24] ),
    .A2(_12542_),
    .A3(_12723_),
    .B1(_12659_),
    .C1(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__o22a_2 _17763_ (.A1(\decode.regfile.registers_14[24] ),
    .A2(_12670_),
    .B1(_03151_),
    .B2(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__o31a_2 _17764_ (.A1(\decode.regfile.registers_15[24] ),
    .A2(_12667_),
    .A3(_12773_),
    .B1(_13011_),
    .X(_03167_));
 sky130_fd_sc_hd__o21a_2 _17765_ (.A1(_12585_),
    .A2(_03166_),
    .B1(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__o22a_2 _17766_ (.A1(\decode.regfile.registers_17[24] ),
    .A2(_12580_),
    .B1(_03150_),
    .B2(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__o2111a_2 _17767_ (.A1(\decode.regfile.registers_18[24] ),
    .A2(_10925_),
    .B1(_12569_),
    .C1(_11023_),
    .D1(_11009_),
    .X(_03170_));
 sky130_fd_sc_hd__a21oi_2 _17768_ (.A1(_03169_),
    .A2(_12566_),
    .B1(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__nor2_2 _17769_ (.A(_03149_),
    .B(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__o221a_2 _17770_ (.A1(\decode.regfile.registers_21[24] ),
    .A2(_12716_),
    .B1(_03148_),
    .B2(_03172_),
    .C1(_13164_),
    .X(_03173_));
 sky130_fd_sc_hd__a211o_2 _17771_ (.A1(\decode.regfile.registers_22[24] ),
    .A2(_13100_),
    .B1(_03173_),
    .C1(_13289_),
    .X(_03174_));
 sky130_fd_sc_hd__or4_2 _17772_ (.A(_11014_),
    .B(_10936_),
    .C(\decode.regfile.registers_23[24] ),
    .D(_12995_),
    .X(_03175_));
 sky130_fd_sc_hd__o2111a_2 _17773_ (.A1(_13250_),
    .A2(\decode.regfile.registers_24[24] ),
    .B1(_12997_),
    .C1(_12998_),
    .D1(_13367_),
    .X(_03176_));
 sky130_fd_sc_hd__a31o_2 _17774_ (.A1(_13339_),
    .A2(_03174_),
    .A3(_03175_),
    .B1(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__or4_2 _17775_ (.A(_13407_),
    .B(\decode.regfile.registers_25[24] ),
    .C(_13482_),
    .D(_12811_),
    .X(_03178_));
 sky130_fd_sc_hd__o2111a_2 _17776_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[24] ),
    .B1(_13002_),
    .C1(_13484_),
    .D1(_02987_),
    .X(_03179_));
 sky130_fd_sc_hd__a31o_2 _17777_ (.A1(_12968_),
    .A2(_03177_),
    .A3(_03178_),
    .B1(_03179_),
    .X(_03180_));
 sky130_fd_sc_hd__or4_2 _17778_ (.A(_02990_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[24] ),
    .D(_13487_),
    .X(_03181_));
 sky130_fd_sc_hd__o21a_2 _17779_ (.A1(_10929_),
    .A2(\decode.regfile.registers_28[24] ),
    .B1(_02992_),
    .X(_03182_));
 sky130_fd_sc_hd__a31o_2 _17780_ (.A1(_12967_),
    .A2(_03180_),
    .A3(_03181_),
    .B1(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__o221a_2 _17781_ (.A1(_02997_),
    .A2(_12767_),
    .B1(_12965_),
    .B2(\decode.regfile.registers_29[24] ),
    .C1(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__o221a_2 _17782_ (.A1(\decode.regfile.registers_31[24] ),
    .A2(_12872_),
    .B1(_03147_),
    .B2(_03184_),
    .C1(_03073_),
    .X(_00444_));
 sky130_fd_sc_hd__o21a_2 _17783_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[25] ),
    .B1(_13492_),
    .X(_03185_));
 sky130_fd_sc_hd__a41o_2 _17784_ (.A1(\decode.regfile.registers_20[25] ),
    .A2(_12525_),
    .A3(_12552_),
    .A4(_12823_),
    .B1(_12824_),
    .X(_03186_));
 sky130_fd_sc_hd__o21ai_2 _17785_ (.A1(\decode.regfile.registers_19[25] ),
    .A2(_12679_),
    .B1(_12906_),
    .Y(_03187_));
 sky130_fd_sc_hd__a41o_2 _17786_ (.A1(\decode.regfile.registers_17[25] ),
    .A2(_12524_),
    .A3(_12568_),
    .A4(_12535_),
    .B1(_12571_),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_2 _17787_ (.A0(\decode.regfile.registers_4[25] ),
    .A1(\decode.regfile.registers_5[25] ),
    .S(_10616_),
    .X(_03189_));
 sky130_fd_sc_hd__o2bb2a_2 _17788_ (.A1_N(\decode.regfile.registers_3[25] ),
    .A2_N(_12836_),
    .B1(_10610_),
    .B2(_12626_),
    .X(_03190_));
 sky130_fd_sc_hd__a31o_2 _17789_ (.A1(\decode.regfile.registers_1[25] ),
    .A2(_12636_),
    .A3(_13145_),
    .B1(_12835_),
    .X(_03191_));
 sky130_fd_sc_hd__a21o_2 _17790_ (.A1(\decode.regfile.registers_0[25] ),
    .A2(_12778_),
    .B1(_03191_),
    .X(_03192_));
 sky130_fd_sc_hd__o211ai_2 _17791_ (.A1(\decode.regfile.registers_2[25] ),
    .A2(_12634_),
    .B1(_12629_),
    .C1(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__a2bb2oi_2 _17792_ (.A1_N(_12732_),
    .A2_N(_03189_),
    .B1(_03190_),
    .B2(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__o32a_2 _17793_ (.A1(\decode.regfile.registers_6[25] ),
    .A2(_10603_),
    .A3(_12615_),
    .B1(_12623_),
    .B2(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__o32a_2 _17794_ (.A1(_12498_),
    .A2(_12540_),
    .A3(_12977_),
    .B1(\decode.regfile.registers_7[25] ),
    .B2(_12645_),
    .X(_03196_));
 sky130_fd_sc_hd__o21ai_2 _17795_ (.A1(_12612_),
    .A2(_03195_),
    .B1(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__a21oi_2 _17796_ (.A1(\decode.regfile.registers_8[25] ),
    .A2(_12889_),
    .B1(_12607_),
    .Y(_03198_));
 sky130_fd_sc_hd__nand2_2 _17797_ (.A(_03197_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__o41a_2 _17798_ (.A1(\decode.regfile.registers_9[25] ),
    .A2(_11019_),
    .A3(_12504_),
    .A4(_12511_),
    .B1(_12654_),
    .X(_03200_));
 sky130_fd_sc_hd__a22oi_2 _17799_ (.A1(\decode.regfile.registers_10[25] ),
    .A2(_12600_),
    .B1(_03199_),
    .B2(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__o2bb2a_2 _17800_ (.A1_N(\decode.regfile.registers_11[25] ),
    .A2_N(_12595_),
    .B1(_12772_),
    .B2(_12541_),
    .X(_03202_));
 sky130_fd_sc_hd__o21ai_2 _17801_ (.A1(_12595_),
    .A2(_03201_),
    .B1(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__o32a_2 _17802_ (.A1(_11020_),
    .A2(_12490_),
    .A3(_12512_),
    .B1(\decode.regfile.registers_12[25] ),
    .B2(_12591_),
    .X(_03204_));
 sky130_fd_sc_hd__a221oi_2 _17803_ (.A1(\decode.regfile.registers_13[25] ),
    .A2(_12775_),
    .B1(_03203_),
    .B2(_03204_),
    .C1(_12664_),
    .Y(_03205_));
 sky130_fd_sc_hd__nor2_2 _17804_ (.A(\decode.regfile.registers_14[25] ),
    .B(_12670_),
    .Y(_03206_));
 sky130_fd_sc_hd__a21oi_2 _17805_ (.A1(\decode.regfile.registers_15[25] ),
    .A2(_12585_),
    .B1(_12673_),
    .Y(_03207_));
 sky130_fd_sc_hd__o31ai_2 _17806_ (.A1(_12585_),
    .A2(_03205_),
    .A3(_03206_),
    .B1(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__o211a_2 _17807_ (.A1(\decode.regfile.registers_16[25] ),
    .A2(_12576_),
    .B1(_12719_),
    .C1(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__o22a_2 _17808_ (.A1(\decode.regfile.registers_18[25] ),
    .A2(_12566_),
    .B1(_03188_),
    .B2(_03209_),
    .X(_03210_));
 sky130_fd_sc_hd__nor2_2 _17809_ (.A(_12562_),
    .B(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__nor2_2 _17810_ (.A(_03187_),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__o221a_2 _17811_ (.A1(\decode.regfile.registers_21[25] ),
    .A2(_12716_),
    .B1(_03186_),
    .B2(_03212_),
    .C1(_13164_),
    .X(_03213_));
 sky130_fd_sc_hd__a211o_2 _17812_ (.A1(\decode.regfile.registers_22[25] ),
    .A2(_13100_),
    .B1(_03213_),
    .C1(_13289_),
    .X(_03214_));
 sky130_fd_sc_hd__or4_2 _17813_ (.A(_11014_),
    .B(_10936_),
    .C(\decode.regfile.registers_23[25] ),
    .D(_12995_),
    .X(_03215_));
 sky130_fd_sc_hd__o2111a_2 _17814_ (.A1(_12712_),
    .A2(\decode.regfile.registers_24[25] ),
    .B1(_12997_),
    .C1(_12998_),
    .D1(_13367_),
    .X(_03216_));
 sky130_fd_sc_hd__a31o_2 _17815_ (.A1(_13339_),
    .A2(_03214_),
    .A3(_03215_),
    .B1(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__or4_2 _17816_ (.A(_13407_),
    .B(\decode.regfile.registers_25[25] ),
    .C(_13482_),
    .D(_12811_),
    .X(_03218_));
 sky130_fd_sc_hd__o2111a_2 _17817_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[25] ),
    .B1(_13002_),
    .C1(_13484_),
    .D1(_02987_),
    .X(_03219_));
 sky130_fd_sc_hd__a31o_2 _17818_ (.A1(_12968_),
    .A2(_03217_),
    .A3(_03218_),
    .B1(_03219_),
    .X(_03220_));
 sky130_fd_sc_hd__or4_2 _17819_ (.A(_02990_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[25] ),
    .D(_13487_),
    .X(_03221_));
 sky130_fd_sc_hd__o21a_2 _17820_ (.A1(_10929_),
    .A2(\decode.regfile.registers_28[25] ),
    .B1(_02992_),
    .X(_03222_));
 sky130_fd_sc_hd__a31o_2 _17821_ (.A1(_12967_),
    .A2(_03220_),
    .A3(_03221_),
    .B1(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__o221a_2 _17822_ (.A1(_02997_),
    .A2(_12767_),
    .B1(_12965_),
    .B2(\decode.regfile.registers_29[25] ),
    .C1(_03223_),
    .X(_03224_));
 sky130_fd_sc_hd__o221a_2 _17823_ (.A1(\decode.regfile.registers_31[25] ),
    .A2(_12872_),
    .B1(_03185_),
    .B2(_03224_),
    .C1(_03073_),
    .X(_00445_));
 sky130_fd_sc_hd__o21a_2 _17824_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[26] ),
    .B1(_13492_),
    .X(_03225_));
 sky130_fd_sc_hd__a41o_2 _17825_ (.A1(\decode.regfile.registers_20[26] ),
    .A2(_12546_),
    .A3(_12553_),
    .A4(_12554_),
    .B1(_12538_),
    .X(_03226_));
 sky130_fd_sc_hd__a21o_2 _17826_ (.A1(\decode.regfile.registers_18[26] ),
    .A2(_12572_),
    .B1(_12562_),
    .X(_03227_));
 sky130_fd_sc_hd__a32o_2 _17827_ (.A1(_12524_),
    .A2(_12568_),
    .A3(_12535_),
    .B1(_12674_),
    .B2(\decode.regfile.registers_16[26] ),
    .X(_03228_));
 sky130_fd_sc_hd__a22o_2 _17828_ (.A1(\decode.regfile.registers_11[26] ),
    .A2(_12724_),
    .B1(_12587_),
    .B2(_12551_),
    .X(_03229_));
 sky130_fd_sc_hd__a21oi_2 _17829_ (.A1(\decode.regfile.registers_8[26] ),
    .A2(_12889_),
    .B1(_12607_),
    .Y(_03230_));
 sky130_fd_sc_hd__a221o_2 _17830_ (.A1(\decode.regfile.registers_4[26] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[26] ),
    .C1(_12737_),
    .X(_03231_));
 sky130_fd_sc_hd__a31o_2 _17831_ (.A1(_12530_),
    .A2(_10591_),
    .A3(_12557_),
    .B1(\decode.regfile.registers_0[26] ),
    .X(_03232_));
 sky130_fd_sc_hd__o221a_2 _17832_ (.A1(\decode.regfile.registers_1[26] ),
    .A2(_12631_),
    .B1(_12933_),
    .B2(_12508_),
    .C1(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__a211o_2 _17833_ (.A1(\decode.regfile.registers_2[26] ),
    .A2(_12835_),
    .B1(_12836_),
    .C1(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__o221a_2 _17834_ (.A1(_10610_),
    .A2(_12626_),
    .B1(_12629_),
    .B2(\decode.regfile.registers_3[26] ),
    .C1(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__o32a_2 _17835_ (.A1(\decode.regfile.registers_6[26] ),
    .A2(_10603_),
    .A3(_12615_),
    .B1(_03231_),
    .B2(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__o32a_2 _17836_ (.A1(_12497_),
    .A2(_12539_),
    .A3(_12503_),
    .B1(\decode.regfile.registers_7[26] ),
    .B2(_12645_),
    .X(_03237_));
 sky130_fd_sc_hd__o21ai_2 _17837_ (.A1(_12612_),
    .A2(_03236_),
    .B1(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__a2bb2o_2 _17838_ (.A1_N(\decode.regfile.registers_9[26] ),
    .A2_N(_12603_),
    .B1(_03230_),
    .B2(_03238_),
    .X(_03239_));
 sky130_fd_sc_hd__o21ai_2 _17839_ (.A1(\decode.regfile.registers_10[26] ),
    .A2(_12654_),
    .B1(_12878_),
    .Y(_03240_));
 sky130_fd_sc_hd__a21oi_2 _17840_ (.A1(_12654_),
    .A2(_03239_),
    .B1(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__o32a_2 _17841_ (.A1(\decode.regfile.registers_12[26] ),
    .A2(_12542_),
    .A3(_12723_),
    .B1(_03229_),
    .B2(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__and3_2 _17842_ (.A(\decode.regfile.registers_13[26] ),
    .B(_12534_),
    .C(_12588_),
    .X(_03243_));
 sky130_fd_sc_hd__a211o_2 _17843_ (.A1(_03242_),
    .A2(_12659_),
    .B1(_12664_),
    .C1(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__o32a_2 _17844_ (.A1(_11021_),
    .A2(_12491_),
    .A3(_12666_),
    .B1(\decode.regfile.registers_14[26] ),
    .B2(_12670_),
    .X(_03245_));
 sky130_fd_sc_hd__a22o_2 _17845_ (.A1(\decode.regfile.registers_15[26] ),
    .A2(_12585_),
    .B1(_03244_),
    .B2(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__o41a_2 _17846_ (.A1(_10595_),
    .A2(_10599_),
    .A3(_10588_),
    .A4(_12542_),
    .B1(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__o221a_2 _17847_ (.A1(\decode.regfile.registers_17[26] ),
    .A2(_12580_),
    .B1(_03228_),
    .B2(_03247_),
    .C1(_12566_),
    .X(_03248_));
 sky130_fd_sc_hd__o221a_2 _17848_ (.A1(\decode.regfile.registers_19[26] ),
    .A2(_12679_),
    .B1(_03227_),
    .B2(_03248_),
    .C1(_12545_),
    .X(_03249_));
 sky130_fd_sc_hd__o221ai_2 _17849_ (.A1(\decode.regfile.registers_21[26] ),
    .A2(_12682_),
    .B1(_03226_),
    .B2(_03249_),
    .C1(_12806_),
    .Y(_03250_));
 sky130_fd_sc_hd__a21oi_2 _17850_ (.A1(\decode.regfile.registers_22[26] ),
    .A2(_12527_),
    .B1(_12687_),
    .Y(_03251_));
 sky130_fd_sc_hd__nand2_2 _17851_ (.A(_03250_),
    .B(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__or4_2 _17852_ (.A(_11014_),
    .B(_10936_),
    .C(\decode.regfile.registers_23[26] ),
    .D(_12995_),
    .X(_03253_));
 sky130_fd_sc_hd__o2111a_2 _17853_ (.A1(_12712_),
    .A2(\decode.regfile.registers_24[26] ),
    .B1(_12997_),
    .C1(_12998_),
    .D1(_13367_),
    .X(_03254_));
 sky130_fd_sc_hd__a31o_2 _17854_ (.A1(_13339_),
    .A2(_03252_),
    .A3(_03253_),
    .B1(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__or4_2 _17855_ (.A(_10938_),
    .B(\decode.regfile.registers_25[26] ),
    .C(_13482_),
    .D(_12811_),
    .X(_03256_));
 sky130_fd_sc_hd__o2111a_2 _17856_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[26] ),
    .B1(_13002_),
    .C1(_13484_),
    .D1(_02987_),
    .X(_03257_));
 sky130_fd_sc_hd__a31o_2 _17857_ (.A1(_12968_),
    .A2(_03255_),
    .A3(_03256_),
    .B1(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__or4_2 _17858_ (.A(_02990_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[26] ),
    .D(_13487_),
    .X(_03259_));
 sky130_fd_sc_hd__o21a_2 _17859_ (.A1(_10929_),
    .A2(\decode.regfile.registers_28[26] ),
    .B1(_02992_),
    .X(_03260_));
 sky130_fd_sc_hd__a31o_2 _17860_ (.A1(_12967_),
    .A2(_03258_),
    .A3(_03259_),
    .B1(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__o221a_2 _17861_ (.A1(_02997_),
    .A2(_12767_),
    .B1(_12965_),
    .B2(\decode.regfile.registers_29[26] ),
    .C1(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__o221a_2 _17862_ (.A1(\decode.regfile.registers_31[26] ),
    .A2(_12872_),
    .B1(_03225_),
    .B2(_03262_),
    .C1(_03073_),
    .X(_00446_));
 sky130_fd_sc_hd__o21a_2 _17863_ (.A1(_13451_),
    .A2(\decode.regfile.registers_30[27] ),
    .B1(_13492_),
    .X(_03263_));
 sky130_fd_sc_hd__a21o_2 _17864_ (.A1(\decode.regfile.registers_18[27] ),
    .A2(_12571_),
    .B1(_12560_),
    .X(_03264_));
 sky130_fd_sc_hd__and4_2 _17865_ (.A(\decode.regfile.registers_17[27] ),
    .B(_11021_),
    .C(_12559_),
    .D(_12534_),
    .X(_03265_));
 sky130_fd_sc_hd__a41o_2 _17866_ (.A1(\decode.regfile.registers_15[27] ),
    .A2(_10611_),
    .A3(_10618_),
    .A4(_12588_),
    .B1(_12672_),
    .X(_03266_));
 sky130_fd_sc_hd__o2111a_2 _17867_ (.A1(\decode.regfile.registers_10[27] ),
    .A2(_10617_),
    .B1(_12776_),
    .C1(_10610_),
    .D1(_12604_),
    .X(_03267_));
 sky130_fd_sc_hd__a221o_2 _17868_ (.A1(\decode.regfile.registers_7[27] ),
    .A2(_12610_),
    .B1(_12622_),
    .B2(\decode.regfile.registers_6[27] ),
    .C1(_12843_),
    .X(_03268_));
 sky130_fd_sc_hd__a31o_2 _17869_ (.A1(\decode.regfile.registers_3[27] ),
    .A2(_10615_),
    .A3(_12728_),
    .B1(_12837_),
    .X(_03269_));
 sky130_fd_sc_hd__or2b_2 _17870_ (.A(_10614_),
    .B_N(\decode.regfile.registers_2[27] ),
    .X(_03270_));
 sky130_fd_sc_hd__nand2_2 _17871_ (.A(_12630_),
    .B(\decode.regfile.registers_0[27] ),
    .Y(_03271_));
 sky130_fd_sc_hd__o221a_2 _17872_ (.A1(_12315_),
    .A2(_12630_),
    .B1(_12829_),
    .B2(_10614_),
    .C1(_03271_),
    .X(_03272_));
 sky130_fd_sc_hd__a21oi_2 _17873_ (.A1(_12729_),
    .A2(_03270_),
    .B1(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__a221o_2 _17874_ (.A1(\decode.regfile.registers_4[27] ),
    .A2(_12548_),
    .B1(_12531_),
    .B2(\decode.regfile.registers_5[27] ),
    .C1(_12625_),
    .X(_03274_));
 sky130_fd_sc_hd__o21a_2 _17875_ (.A1(_03269_),
    .A2(_03273_),
    .B1(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__o22ai_2 _17876_ (.A1(\decode.regfile.registers_8[27] ),
    .A2(_12725_),
    .B1(_03268_),
    .B2(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand2_2 _17877_ (.A(_12601_),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__o211a_2 _17878_ (.A1(_12602_),
    .A2(\decode.regfile.registers_9[27] ),
    .B1(_12652_),
    .C1(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__o22ai_2 _17879_ (.A1(\decode.regfile.registers_11[27] ),
    .A2(_12792_),
    .B1(_03267_),
    .B2(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__o21ai_2 _17880_ (.A1(_12541_),
    .A2(_12722_),
    .B1(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__or4_2 _17881_ (.A(\decode.regfile.registers_12[27] ),
    .B(_12489_),
    .C(_12498_),
    .D(_12540_),
    .X(_03281_));
 sky130_fd_sc_hd__a31o_2 _17882_ (.A1(\decode.regfile.registers_13[27] ),
    .A2(_12533_),
    .A3(_12582_),
    .B1(_12662_),
    .X(_03282_));
 sky130_fd_sc_hd__a31o_2 _17883_ (.A1(_12658_),
    .A2(_03280_),
    .A3(_03281_),
    .B1(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__o221a_2 _17884_ (.A1(_12650_),
    .A2(_12723_),
    .B1(_12669_),
    .B2(\decode.regfile.registers_14[27] ),
    .C1(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__o221a_2 _17885_ (.A1(\decode.regfile.registers_16[27] ),
    .A2(_12575_),
    .B1(_03266_),
    .B2(_03284_),
    .C1(_12578_),
    .X(_03285_));
 sky130_fd_sc_hd__o21a_2 _17886_ (.A1(_03265_),
    .A2(_03285_),
    .B1(_12565_),
    .X(_03286_));
 sky130_fd_sc_hd__o221a_2 _17887_ (.A1(\decode.regfile.registers_19[27] ),
    .A2(_12678_),
    .B1(_03264_),
    .B2(_03286_),
    .C1(_12544_),
    .X(_03287_));
 sky130_fd_sc_hd__a211o_2 _17888_ (.A1(\decode.regfile.registers_20[27] ),
    .A2(_12770_),
    .B1(_03287_),
    .C1(_12537_),
    .X(_03288_));
 sky130_fd_sc_hd__o211a_2 _17889_ (.A1(_12822_),
    .A2(\decode.regfile.registers_21[27] ),
    .B1(_13164_),
    .C1(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__a211o_2 _17890_ (.A1(\decode.regfile.registers_22[27] ),
    .A2(_13100_),
    .B1(_03289_),
    .C1(_13289_),
    .X(_03290_));
 sky130_fd_sc_hd__or4_2 _17891_ (.A(_11014_),
    .B(_10936_),
    .C(\decode.regfile.registers_23[27] ),
    .D(_12995_),
    .X(_03291_));
 sky130_fd_sc_hd__o2111a_2 _17892_ (.A1(_12712_),
    .A2(\decode.regfile.registers_24[27] ),
    .B1(_12997_),
    .C1(_12998_),
    .D1(_11025_),
    .X(_03292_));
 sky130_fd_sc_hd__a31o_2 _17893_ (.A1(_12515_),
    .A2(_03290_),
    .A3(_03291_),
    .B1(_03292_),
    .X(_03293_));
 sky130_fd_sc_hd__or4_2 _17894_ (.A(_10938_),
    .B(\decode.regfile.registers_25[27] ),
    .C(_13482_),
    .D(_12811_),
    .X(_03294_));
 sky130_fd_sc_hd__o2111a_2 _17895_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[27] ),
    .B1(_13002_),
    .C1(_13484_),
    .D1(_02987_),
    .X(_03295_));
 sky130_fd_sc_hd__a31o_2 _17896_ (.A1(_12968_),
    .A2(_03293_),
    .A3(_03294_),
    .B1(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__or4_2 _17897_ (.A(_02990_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[27] ),
    .D(_13487_),
    .X(_03297_));
 sky130_fd_sc_hd__o21a_2 _17898_ (.A1(_10929_),
    .A2(\decode.regfile.registers_28[27] ),
    .B1(_02992_),
    .X(_03298_));
 sky130_fd_sc_hd__a31o_2 _17899_ (.A1(_12967_),
    .A2(_03296_),
    .A3(_03297_),
    .B1(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__o221a_2 _17900_ (.A1(_02997_),
    .A2(_12767_),
    .B1(_12965_),
    .B2(\decode.regfile.registers_29[27] ),
    .C1(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__o221a_2 _17901_ (.A1(\decode.regfile.registers_31[27] ),
    .A2(_12872_),
    .B1(_03263_),
    .B2(_03300_),
    .C1(_03073_),
    .X(_00447_));
 sky130_fd_sc_hd__o21a_2 _17902_ (.A1(_12765_),
    .A2(\decode.regfile.registers_30[28] ),
    .B1(_13492_),
    .X(_03301_));
 sky130_fd_sc_hd__o2111a_2 _17903_ (.A1(_10927_),
    .A2(\decode.regfile.registers_24[28] ),
    .B1(_10933_),
    .C1(_12759_),
    .D1(_12862_),
    .X(_03302_));
 sky130_fd_sc_hd__o2111a_2 _17904_ (.A1(_10926_),
    .A2(\decode.regfile.registers_22[28] ),
    .B1(_12554_),
    .C1(_11009_),
    .D1(_12546_),
    .X(_03303_));
 sky130_fd_sc_hd__a41o_2 _17905_ (.A1(\decode.regfile.registers_20[28] ),
    .A2(_11024_),
    .A3(_12553_),
    .A4(_12554_),
    .B1(_12537_),
    .X(_03304_));
 sky130_fd_sc_hd__a41o_2 _17906_ (.A1(\decode.regfile.registers_15[28] ),
    .A2(_12555_),
    .A3(_10619_),
    .A4(_12876_),
    .B1(_13031_),
    .X(_03305_));
 sky130_fd_sc_hd__a31o_2 _17907_ (.A1(\decode.regfile.registers_13[28] ),
    .A2(_12927_),
    .A3(_12583_),
    .B1(_12663_),
    .X(_03306_));
 sky130_fd_sc_hd__o2111a_2 _17908_ (.A1(\decode.regfile.registers_10[28] ),
    .A2(_10617_),
    .B1(_12776_),
    .C1(_10611_),
    .D1(_12604_),
    .X(_03307_));
 sky130_fd_sc_hd__a221oi_2 _17909_ (.A1(\decode.regfile.registers_2[28] ),
    .A2(_12834_),
    .B1(_12638_),
    .B2(\decode.regfile.registers_3[28] ),
    .C1(_12837_),
    .Y(_03308_));
 sky130_fd_sc_hd__a31o_2 _17910_ (.A1(_12530_),
    .A2(_12616_),
    .A3(_12557_),
    .B1(\decode.regfile.registers_0[28] ),
    .X(_03309_));
 sky130_fd_sc_hd__o211ai_2 _17911_ (.A1(\decode.regfile.registers_1[28] ),
    .A2(_12631_),
    .B1(_12933_),
    .C1(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__nand2_2 _17912_ (.A(_03308_),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__a221o_2 _17913_ (.A1(\decode.regfile.registers_4[28] ),
    .A2(_12547_),
    .B1(_12531_),
    .B2(\decode.regfile.registers_5[28] ),
    .C1(_12625_),
    .X(_03312_));
 sky130_fd_sc_hd__a32o_2 _17914_ (.A1(\decode.regfile.registers_7[28] ),
    .A2(_10615_),
    .A3(_13020_),
    .B1(_12621_),
    .B2(\decode.regfile.registers_6[28] ),
    .X(_03313_));
 sky130_fd_sc_hd__a21o_2 _17915_ (.A1(_03311_),
    .A2(_03312_),
    .B1(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__and4_2 _17916_ (.A(\decode.regfile.registers_8[28] ),
    .B(_12592_),
    .C(_10593_),
    .D(_12549_),
    .X(_03315_));
 sky130_fd_sc_hd__a211o_2 _17917_ (.A1(_12726_),
    .A2(_03314_),
    .B1(_03315_),
    .C1(_12606_),
    .X(_03316_));
 sky130_fd_sc_hd__o211a_2 _17918_ (.A1(_12602_),
    .A2(\decode.regfile.registers_9[28] ),
    .B1(_12653_),
    .C1(_03316_),
    .X(_03317_));
 sky130_fd_sc_hd__o22a_2 _17919_ (.A1(\decode.regfile.registers_11[28] ),
    .A2(_12792_),
    .B1(_03307_),
    .B2(_03317_),
    .X(_03318_));
 sky130_fd_sc_hd__or4_2 _17920_ (.A(\decode.regfile.registers_12[28] ),
    .B(_12489_),
    .C(_11019_),
    .D(_12540_),
    .X(_03319_));
 sky130_fd_sc_hd__o221a_2 _17921_ (.A1(_12512_),
    .A2(_12772_),
    .B1(_12794_),
    .B2(_03318_),
    .C1(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__o221a_2 _17922_ (.A1(\decode.regfile.registers_14[28] ),
    .A2(_12984_),
    .B1(_03306_),
    .B2(_03320_),
    .C1(_12874_),
    .X(_03321_));
 sky130_fd_sc_hd__o221a_2 _17923_ (.A1(\decode.regfile.registers_16[28] ),
    .A2(_13011_),
    .B1(_03305_),
    .B2(_03321_),
    .C1(_12578_),
    .X(_03322_));
 sky130_fd_sc_hd__a41o_2 _17924_ (.A1(\decode.regfile.registers_17[28] ),
    .A2(_12524_),
    .A3(_12568_),
    .A4(_12535_),
    .B1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__o2111a_2 _17925_ (.A1(\decode.regfile.registers_18[28] ),
    .A2(_10924_),
    .B1(_12568_),
    .C1(_12524_),
    .D1(_11008_),
    .X(_03324_));
 sky130_fd_sc_hd__a21o_2 _17926_ (.A1(_12566_),
    .A2(_03323_),
    .B1(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__o211a_2 _17927_ (.A1(\decode.regfile.registers_19[28] ),
    .A2(_12679_),
    .B1(_12545_),
    .C1(_03325_),
    .X(_03326_));
 sky130_fd_sc_hd__o221a_2 _17928_ (.A1(\decode.regfile.registers_21[28] ),
    .A2(_12682_),
    .B1(_03304_),
    .B2(_03326_),
    .C1(_12806_),
    .X(_03327_));
 sky130_fd_sc_hd__o221a_2 _17929_ (.A1(\decode.regfile.registers_23[28] ),
    .A2(_12714_),
    .B1(_03303_),
    .B2(_03327_),
    .C1(_12515_),
    .X(_03328_));
 sky130_fd_sc_hd__o22a_2 _17930_ (.A1(_12513_),
    .A2(\decode.regfile.registers_25[28] ),
    .B1(_03302_),
    .B2(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__o2111a_2 _17931_ (.A1(_10928_),
    .A2(\decode.regfile.registers_26[28] ),
    .B1(_12814_),
    .C1(_11011_),
    .D1(_11027_),
    .X(_03330_));
 sky130_fd_sc_hd__a21o_2 _17932_ (.A1(_03329_),
    .A2(_12695_),
    .B1(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__or4_2 _17933_ (.A(_02990_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[28] ),
    .D(_12506_),
    .X(_03332_));
 sky130_fd_sc_hd__o21a_2 _17934_ (.A1(_10929_),
    .A2(\decode.regfile.registers_28[28] ),
    .B1(_02992_),
    .X(_03333_));
 sky130_fd_sc_hd__a31o_2 _17935_ (.A1(_12967_),
    .A2(_03331_),
    .A3(_03332_),
    .B1(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__o221a_2 _17936_ (.A1(_02997_),
    .A2(_12767_),
    .B1(_12965_),
    .B2(\decode.regfile.registers_29[28] ),
    .C1(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__o221a_2 _17937_ (.A1(_12708_),
    .A2(\decode.regfile.registers_31[28] ),
    .B1(_03301_),
    .B2(_03335_),
    .C1(_03073_),
    .X(_00448_));
 sky130_fd_sc_hd__o21a_2 _17938_ (.A1(_12765_),
    .A2(\decode.regfile.registers_30[29] ),
    .B1(_12486_),
    .X(_03336_));
 sky130_fd_sc_hd__o2111a_2 _17939_ (.A1(_10926_),
    .A2(\decode.regfile.registers_22[29] ),
    .B1(_12554_),
    .C1(_11009_),
    .D1(_12546_),
    .X(_03337_));
 sky130_fd_sc_hd__a41o_2 _17940_ (.A1(\decode.regfile.registers_20[29] ),
    .A2(_12525_),
    .A3(_12552_),
    .A4(_12523_),
    .B1(_12536_),
    .X(_03338_));
 sky130_fd_sc_hd__a41o_2 _17941_ (.A1(\decode.regfile.registers_17[29] ),
    .A2(_11022_),
    .A3(_12567_),
    .A4(_12586_),
    .B1(_12570_),
    .X(_03339_));
 sky130_fd_sc_hd__o21ai_2 _17942_ (.A1(\decode.regfile.registers_10[29] ),
    .A2(_12790_),
    .B1(_12792_),
    .Y(_03340_));
 sky130_fd_sc_hd__mux2_2 _17943_ (.A0(\decode.regfile.registers_4[29] ),
    .A1(\decode.regfile.registers_5[29] ),
    .S(_10615_),
    .X(_03341_));
 sky130_fd_sc_hd__nand2_2 _17944_ (.A(_12631_),
    .B(\decode.regfile.registers_0[29] ),
    .Y(_03342_));
 sky130_fd_sc_hd__o221ai_2 _17945_ (.A1(_12387_),
    .A2(_12932_),
    .B1(_10615_),
    .B2(_12933_),
    .C1(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__o211ai_2 _17946_ (.A1(\decode.regfile.registers_2[29] ),
    .A2(_12634_),
    .B1(_12628_),
    .C1(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__o2bb2a_2 _17947_ (.A1_N(\decode.regfile.registers_3[29] ),
    .A2_N(_12639_),
    .B1(_10609_),
    .B2(_12625_),
    .X(_03345_));
 sky130_fd_sc_hd__a2bb2o_2 _17948_ (.A1_N(_12732_),
    .A2_N(_03341_),
    .B1(_03344_),
    .B2(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__nand2_2 _17949_ (.A(_12880_),
    .B(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__o221ai_2 _17950_ (.A1(_12649_),
    .A2(_12615_),
    .B1(_12880_),
    .B2(\decode.regfile.registers_6[29] ),
    .C1(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__a21oi_2 _17951_ (.A1(\decode.regfile.registers_7[29] ),
    .A2(_12611_),
    .B1(_12889_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand2_2 _17952_ (.A(_03348_),
    .B(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__o32a_2 _17953_ (.A1(_11018_),
    .A2(_12977_),
    .A3(_12510_),
    .B1(\decode.regfile.registers_8[29] ),
    .B2(_12892_),
    .X(_03351_));
 sky130_fd_sc_hd__a221oi_2 _17954_ (.A1(\decode.regfile.registers_9[29] ),
    .A2(_12607_),
    .B1(_03350_),
    .B2(_03351_),
    .C1(_12600_),
    .Y(_03352_));
 sky130_fd_sc_hd__or4b_2 _17955_ (.A(_12498_),
    .B(_12977_),
    .C(_12649_),
    .D_N(\decode.regfile.registers_11[29] ),
    .X(_03353_));
 sky130_fd_sc_hd__o211ai_2 _17956_ (.A1(_03340_),
    .A2(_03352_),
    .B1(_12591_),
    .C1(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__o32a_2 _17957_ (.A1(_11019_),
    .A2(_12489_),
    .A3(_12511_),
    .B1(\decode.regfile.registers_12[29] ),
    .B2(_12745_),
    .X(_03355_));
 sky130_fd_sc_hd__a221o_2 _17958_ (.A1(\decode.regfile.registers_13[29] ),
    .A2(_12775_),
    .B1(_03354_),
    .B2(_03355_),
    .C1(_12663_),
    .X(_03356_));
 sky130_fd_sc_hd__o32a_2 _17959_ (.A1(_11020_),
    .A2(_12491_),
    .A3(_12650_),
    .B1(\decode.regfile.registers_14[29] ),
    .B2(_12669_),
    .X(_03357_));
 sky130_fd_sc_hd__a221o_2 _17960_ (.A1(\decode.regfile.registers_15[29] ),
    .A2(_12584_),
    .B1(_03356_),
    .B2(_03357_),
    .C1(_13031_),
    .X(_03358_));
 sky130_fd_sc_hd__o211a_2 _17961_ (.A1(\decode.regfile.registers_16[29] ),
    .A2(_13011_),
    .B1(_12579_),
    .C1(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__o22a_2 _17962_ (.A1(\decode.regfile.registers_18[29] ),
    .A2(_12565_),
    .B1(_03339_),
    .B2(_03359_),
    .X(_03360_));
 sky130_fd_sc_hd__or4_2 _17963_ (.A(\decode.regfile.registers_19[29] ),
    .B(_10599_),
    .C(_10588_),
    .D(_12518_),
    .X(_03361_));
 sky130_fd_sc_hd__o211a_2 _17964_ (.A1(_12561_),
    .A2(_03360_),
    .B1(_03361_),
    .C1(_12906_),
    .X(_03362_));
 sky130_fd_sc_hd__o221a_2 _17965_ (.A1(\decode.regfile.registers_21[29] ),
    .A2(_12716_),
    .B1(_03338_),
    .B2(_03362_),
    .C1(_12909_),
    .X(_03363_));
 sky130_fd_sc_hd__o221a_2 _17966_ (.A1(\decode.regfile.registers_23[29] ),
    .A2(_12714_),
    .B1(_03337_),
    .B2(_03363_),
    .C1(_12514_),
    .X(_03364_));
 sky130_fd_sc_hd__o2111a_2 _17967_ (.A1(_12712_),
    .A2(\decode.regfile.registers_24[29] ),
    .B1(_12997_),
    .C1(_12690_),
    .D1(_11025_),
    .X(_03365_));
 sky130_fd_sc_hd__or2_2 _17968_ (.A(_03364_),
    .B(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__or4_2 _17969_ (.A(_10938_),
    .B(\decode.regfile.registers_25[29] ),
    .C(_12505_),
    .D(_12811_),
    .X(_03367_));
 sky130_fd_sc_hd__o2111a_2 _17970_ (.A1(_02986_),
    .A2(\decode.regfile.registers_26[29] ),
    .B1(_13002_),
    .C1(_11010_),
    .D1(_02987_),
    .X(_03368_));
 sky130_fd_sc_hd__a31o_2 _17971_ (.A1(_12968_),
    .A2(_03366_),
    .A3(_03367_),
    .B1(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__or4_2 _17972_ (.A(_10939_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[29] ),
    .D(_12506_),
    .X(_03370_));
 sky130_fd_sc_hd__o21a_2 _17973_ (.A1(_10929_),
    .A2(\decode.regfile.registers_28[29] ),
    .B1(_12697_),
    .X(_03371_));
 sky130_fd_sc_hd__a31o_2 _17974_ (.A1(_12967_),
    .A2(_03369_),
    .A3(_03370_),
    .B1(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__o221a_2 _17975_ (.A1(_02997_),
    .A2(_12767_),
    .B1(_12965_),
    .B2(\decode.regfile.registers_29[29] ),
    .C1(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__o221a_2 _17976_ (.A1(_12708_),
    .A2(\decode.regfile.registers_31[29] ),
    .B1(_03336_),
    .B2(_03373_),
    .C1(_03073_),
    .X(_00449_));
 sky130_fd_sc_hd__o21a_2 _17977_ (.A1(_10931_),
    .A2(\decode.regfile.registers_30[30] ),
    .B1(_12487_),
    .X(_03374_));
 sky130_fd_sc_hd__o21a_2 _17978_ (.A1(_10930_),
    .A2(\decode.regfile.registers_28[30] ),
    .B1(_12698_),
    .X(_03375_));
 sky130_fd_sc_hd__a41o_2 _17979_ (.A1(\decode.regfile.registers_20[30] ),
    .A2(_12525_),
    .A3(_12552_),
    .A4(_12823_),
    .B1(_12824_),
    .X(_03376_));
 sky130_fd_sc_hd__o2111a_2 _17980_ (.A1(\decode.regfile.registers_18[30] ),
    .A2(_10925_),
    .B1(_12569_),
    .C1(_11023_),
    .D1(_11008_),
    .X(_03377_));
 sky130_fd_sc_hd__a32o_2 _17981_ (.A1(_11022_),
    .A2(_12567_),
    .A3(_12586_),
    .B1(_12673_),
    .B2(\decode.regfile.registers_16[30] ),
    .X(_03378_));
 sky130_fd_sc_hd__o211a_2 _17982_ (.A1(\decode.regfile.registers_14[30] ),
    .A2(_10619_),
    .B1(_12589_),
    .C1(_10612_),
    .X(_03379_));
 sky130_fd_sc_hd__and3_2 _17983_ (.A(\decode.regfile.registers_13[30] ),
    .B(_12927_),
    .C(_12583_),
    .X(_03380_));
 sky130_fd_sc_hd__a221oi_2 _17984_ (.A1(\decode.regfile.registers_2[30] ),
    .A2(_12834_),
    .B1(_12639_),
    .B2(\decode.regfile.registers_3[30] ),
    .C1(_12837_),
    .Y(_03381_));
 sky130_fd_sc_hd__a31o_2 _17985_ (.A1(_12934_),
    .A2(_10592_),
    .A3(_12558_),
    .B1(\decode.regfile.registers_0[30] ),
    .X(_03382_));
 sky130_fd_sc_hd__o211ai_2 _17986_ (.A1(\decode.regfile.registers_1[30] ),
    .A2(_12932_),
    .B1(_12830_),
    .C1(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__a221oi_2 _17987_ (.A1(\decode.regfile.registers_4[30] ),
    .A2(_12548_),
    .B1(_13145_),
    .B2(\decode.regfile.registers_5[30] ),
    .C1(_12625_),
    .Y(_03384_));
 sky130_fd_sc_hd__a21oi_2 _17988_ (.A1(_03381_),
    .A2(_03383_),
    .B1(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__a221oi_2 _17989_ (.A1(\decode.regfile.registers_7[30] ),
    .A2(_12610_),
    .B1(_12737_),
    .B2(\decode.regfile.registers_6[30] ),
    .C1(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__a21oi_2 _17990_ (.A1(\decode.regfile.registers_8[30] ),
    .A2(_12843_),
    .B1(_12605_),
    .Y(_03387_));
 sky130_fd_sc_hd__o21ai_2 _17991_ (.A1(_12888_),
    .A2(_03386_),
    .B1(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__o211a_2 _17992_ (.A1(_12602_),
    .A2(\decode.regfile.registers_9[30] ),
    .B1(_12652_),
    .C1(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__a211o_2 _17993_ (.A1(\decode.regfile.registers_10[30] ),
    .A2(_12599_),
    .B1(_12594_),
    .C1(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__o41a_2 _17994_ (.A1(\decode.regfile.registers_11[30] ),
    .A2(_12499_),
    .A3(_12504_),
    .A4(_12650_),
    .B1(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__o32a_2 _17995_ (.A1(_12499_),
    .A2(_12490_),
    .A3(_12511_),
    .B1(\decode.regfile.registers_12[30] ),
    .B2(_12745_),
    .X(_03392_));
 sky130_fd_sc_hd__o21a_2 _17996_ (.A1(_12794_),
    .A2(_03391_),
    .B1(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__o32a_2 _17997_ (.A1(_10604_),
    .A2(_10619_),
    .A3(_12773_),
    .B1(_03380_),
    .B2(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__o221a_2 _17998_ (.A1(\decode.regfile.registers_15[30] ),
    .A2(_12874_),
    .B1(_03379_),
    .B2(_03394_),
    .C1(_12576_),
    .X(_03395_));
 sky130_fd_sc_hd__o221a_2 _17999_ (.A1(\decode.regfile.registers_17[30] ),
    .A2(_12719_),
    .B1(_03378_),
    .B2(_03395_),
    .C1(_12826_),
    .X(_03396_));
 sky130_fd_sc_hd__o221a_2 _18000_ (.A1(\decode.regfile.registers_19[30] ),
    .A2(_12678_),
    .B1(_03377_),
    .B2(_03396_),
    .C1(_12906_),
    .X(_03397_));
 sky130_fd_sc_hd__o221a_2 _18001_ (.A1(\decode.regfile.registers_21[30] ),
    .A2(_12716_),
    .B1(_03376_),
    .B2(_03397_),
    .C1(_13164_),
    .X(_03398_));
 sky130_fd_sc_hd__a211o_2 _18002_ (.A1(\decode.regfile.registers_22[30] ),
    .A2(_13100_),
    .B1(_03398_),
    .C1(_13289_),
    .X(_03399_));
 sky130_fd_sc_hd__or4_2 _18003_ (.A(_11014_),
    .B(_10936_),
    .C(\decode.regfile.registers_23[30] ),
    .D(_12995_),
    .X(_03400_));
 sky130_fd_sc_hd__o2111a_2 _18004_ (.A1(_12712_),
    .A2(\decode.regfile.registers_24[30] ),
    .B1(_12997_),
    .C1(_12998_),
    .D1(_11025_),
    .X(_03401_));
 sky130_fd_sc_hd__a31o_2 _18005_ (.A1(_12515_),
    .A2(_03399_),
    .A3(_03400_),
    .B1(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__or4_2 _18006_ (.A(_10938_),
    .B(\decode.regfile.registers_25[30] ),
    .C(_12505_),
    .D(_12811_),
    .X(_03403_));
 sky130_fd_sc_hd__o2111a_2 _18007_ (.A1(_12494_),
    .A2(\decode.regfile.registers_26[30] ),
    .B1(_13002_),
    .C1(_11010_),
    .D1(_11026_),
    .X(_03404_));
 sky130_fd_sc_hd__a31o_2 _18008_ (.A1(_12968_),
    .A2(_03402_),
    .A3(_03403_),
    .B1(_03404_),
    .X(_03405_));
 sky130_fd_sc_hd__o311a_2 _18009_ (.A1(\decode.regfile.registers_27[30] ),
    .A2(_12507_),
    .A3(_12520_),
    .B1(_12967_),
    .C1(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__o221a_2 _18010_ (.A1(_12493_),
    .A2(\decode.regfile.registers_29[30] ),
    .B1(_03375_),
    .B2(_03406_),
    .C1(_12702_),
    .X(_03407_));
 sky130_fd_sc_hd__or4_2 _18011_ (.A(\decode.regfile.registers_31[30] ),
    .B(_12491_),
    .C(_12706_),
    .D(_10940_),
    .X(_03408_));
 sky130_fd_sc_hd__o211a_2 _18012_ (.A1(_03374_),
    .A2(_03407_),
    .B1(_12704_),
    .C1(_03408_),
    .X(_00450_));
 sky130_fd_sc_hd__o21a_2 _18013_ (.A1(_12765_),
    .A2(\decode.regfile.registers_30[31] ),
    .B1(_12486_),
    .X(_03409_));
 sky130_fd_sc_hd__a31o_2 _18014_ (.A1(\decode.regfile.registers_7[31] ),
    .A2(_10617_),
    .A3(_13020_),
    .B1(_12888_),
    .X(_03410_));
 sky130_fd_sc_hd__and2b_2 _18015_ (.A_N(_10616_),
    .B(\decode.regfile.registers_6[31] ),
    .X(_03411_));
 sky130_fd_sc_hd__a221o_2 _18016_ (.A1(\decode.regfile.registers_4[31] ),
    .A2(_12618_),
    .B1(_12620_),
    .B2(\decode.regfile.registers_5[31] ),
    .C1(_12737_),
    .X(_03412_));
 sky130_fd_sc_hd__a31o_2 _18017_ (.A1(_12934_),
    .A2(_10592_),
    .A3(_12558_),
    .B1(\decode.regfile.registers_0[31] ),
    .X(_03413_));
 sky130_fd_sc_hd__o211ai_2 _18018_ (.A1(\decode.regfile.registers_1[31] ),
    .A2(_12778_),
    .B1(_12634_),
    .C1(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__o21ai_2 _18019_ (.A1(\decode.regfile.registers_2[31] ),
    .A2(_12882_),
    .B1(_12729_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2_2 _18020_ (.A(_03414_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__o221a_2 _18021_ (.A1(_10609_),
    .A2(_12614_),
    .B1(_12629_),
    .B2(\decode.regfile.registers_3[31] ),
    .C1(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__o32a_2 _18022_ (.A1(_10603_),
    .A2(_12615_),
    .A3(_03411_),
    .B1(_03412_),
    .B2(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__o22ai_2 _18023_ (.A1(\decode.regfile.registers_8[31] ),
    .A2(_12892_),
    .B1(_03410_),
    .B2(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand2_2 _18024_ (.A(_12603_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__o41a_2 _18025_ (.A1(\decode.regfile.registers_9[31] ),
    .A2(_12498_),
    .A3(_12977_),
    .A4(_12510_),
    .B1(_12653_),
    .X(_03421_));
 sky130_fd_sc_hd__a22oi_2 _18026_ (.A1(\decode.regfile.registers_10[31] ),
    .A2(_12600_),
    .B1(_03420_),
    .B2(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__or4b_2 _18027_ (.A(_11019_),
    .B(_12504_),
    .C(_12649_),
    .D_N(\decode.regfile.registers_11[31] ),
    .X(_03423_));
 sky130_fd_sc_hd__o211ai_2 _18028_ (.A1(_12595_),
    .A2(_03422_),
    .B1(_03423_),
    .C1(_12591_),
    .Y(_03424_));
 sky130_fd_sc_hd__o32a_2 _18029_ (.A1(_12499_),
    .A2(_12490_),
    .A3(_12512_),
    .B1(\decode.regfile.registers_12[31] ),
    .B2(_12745_),
    .X(_03425_));
 sky130_fd_sc_hd__a32o_2 _18030_ (.A1(\decode.regfile.registers_13[31] ),
    .A2(_12927_),
    .A3(_12588_),
    .B1(_03424_),
    .B2(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__o211a_2 _18031_ (.A1(\decode.regfile.registers_14[31] ),
    .A2(_10923_),
    .B1(_12876_),
    .C1(_12555_),
    .X(_03427_));
 sky130_fd_sc_hd__a21o_2 _18032_ (.A1(_12670_),
    .A2(_03426_),
    .B1(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__o311a_2 _18033_ (.A1(\decode.regfile.registers_15[31] ),
    .A2(_12667_),
    .A3(_12773_),
    .B1(_13011_),
    .C1(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__a211o_2 _18034_ (.A1(\decode.regfile.registers_16[31] ),
    .A2(_12674_),
    .B1(_12901_),
    .C1(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__o21a_2 _18035_ (.A1(\decode.regfile.registers_17[31] ),
    .A2(_12719_),
    .B1(_12826_),
    .X(_03431_));
 sky130_fd_sc_hd__a221o_2 _18036_ (.A1(\decode.regfile.registers_18[31] ),
    .A2(_12572_),
    .B1(_03430_),
    .B2(_03431_),
    .C1(_12562_),
    .X(_03432_));
 sky130_fd_sc_hd__o41a_2 _18037_ (.A1(\decode.regfile.registers_19[31] ),
    .A2(_11013_),
    .A3(_10589_),
    .A4(_12519_),
    .B1(_12544_),
    .X(_03433_));
 sky130_fd_sc_hd__a221o_2 _18038_ (.A1(\decode.regfile.registers_20[31] ),
    .A2(_12771_),
    .B1(_03432_),
    .B2(_03433_),
    .C1(_12538_),
    .X(_03434_));
 sky130_fd_sc_hd__o21a_2 _18039_ (.A1(\decode.regfile.registers_21[31] ),
    .A2(_12822_),
    .B1(_12909_),
    .X(_03435_));
 sky130_fd_sc_hd__a221o_2 _18040_ (.A1(\decode.regfile.registers_22[31] ),
    .A2(_12527_),
    .B1(_03434_),
    .B2(_03435_),
    .C1(_12686_),
    .X(_03436_));
 sky130_fd_sc_hd__or4_2 _18041_ (.A(_11014_),
    .B(_10936_),
    .C(\decode.regfile.registers_23[31] ),
    .D(_12995_),
    .X(_03437_));
 sky130_fd_sc_hd__o2111a_2 _18042_ (.A1(_12712_),
    .A2(\decode.regfile.registers_24[31] ),
    .B1(_12997_),
    .C1(_12998_),
    .D1(_11025_),
    .X(_03438_));
 sky130_fd_sc_hd__a31o_2 _18043_ (.A1(_12515_),
    .A2(_03436_),
    .A3(_03437_),
    .B1(_03438_),
    .X(_03439_));
 sky130_fd_sc_hd__or4_2 _18044_ (.A(_10938_),
    .B(\decode.regfile.registers_25[31] ),
    .C(_12505_),
    .D(_12811_),
    .X(_03440_));
 sky130_fd_sc_hd__o2111a_2 _18045_ (.A1(_12494_),
    .A2(\decode.regfile.registers_26[31] ),
    .B1(_13002_),
    .C1(_11010_),
    .D1(_11026_),
    .X(_03441_));
 sky130_fd_sc_hd__a31o_2 _18046_ (.A1(_12968_),
    .A2(_03439_),
    .A3(_03440_),
    .B1(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__or4_2 _18047_ (.A(_10939_),
    .B(_03068_),
    .C(\decode.regfile.registers_27[31] ),
    .D(_12506_),
    .X(_03443_));
 sky130_fd_sc_hd__o21a_2 _18048_ (.A1(_10929_),
    .A2(\decode.regfile.registers_28[31] ),
    .B1(_12697_),
    .X(_03444_));
 sky130_fd_sc_hd__a31o_2 _18049_ (.A1(_12967_),
    .A2(_03442_),
    .A3(_03443_),
    .B1(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__o221a_2 _18050_ (.A1(_10930_),
    .A2(_12767_),
    .B1(_12965_),
    .B2(\decode.regfile.registers_29[31] ),
    .C1(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__o221a_2 _18051_ (.A1(\decode.regfile.registers_31[31] ),
    .A2(_12872_),
    .B1(_03409_),
    .B2(_03446_),
    .C1(_03073_),
    .X(_00451_));
 sky130_fd_sc_hd__and3_2 _18052_ (.A(_10965_),
    .B(_10998_),
    .C(_10969_),
    .X(_03447_));
 sky130_fd_sc_hd__buf_1 _18053_ (.A(_03447_),
    .X(_00452_));
 sky130_fd_sc_hd__and3_2 _18054_ (.A(_10583_),
    .B(_10584_),
    .C(_10998_),
    .X(_03448_));
 sky130_fd_sc_hd__buf_1 _18055_ (.A(_03448_),
    .X(_00453_));
 sky130_fd_sc_hd__buf_1 _18056_ (.A(_09954_),
    .X(_03449_));
 sky130_fd_sc_hd__and4bb_2 _18057_ (.A_N(_10965_),
    .B_N(_10972_),
    .C(_10969_),
    .D(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__buf_1 _18058_ (.A(_03450_),
    .X(_00454_));
 sky130_fd_sc_hd__and4b_2 _18059_ (.A_N(\decode.control.io_opcode[3] ),
    .B(_10583_),
    .C(_10584_),
    .D(_10998_),
    .X(_03451_));
 sky130_fd_sc_hd__buf_1 _18060_ (.A(_03451_),
    .X(_00455_));
 sky130_fd_sc_hd__buf_1 _18061_ (.A(_10910_),
    .X(_03452_));
 sky130_fd_sc_hd__o31ai_2 _18062_ (.A1(_10965_),
    .A2(_10964_),
    .A3(_10951_),
    .B1(_10582_),
    .Y(_03453_));
 sky130_fd_sc_hd__and4b_2 _18063_ (.A_N(_03452_),
    .B(_10916_),
    .C(_03453_),
    .D(_10018_),
    .X(_03454_));
 sky130_fd_sc_hd__buf_1 _18064_ (.A(_03454_),
    .X(_00456_));
 sky130_fd_sc_hd__o21a_2 _18065_ (.A1(_10943_),
    .A2(_10941_),
    .B1(_10581_),
    .X(_03455_));
 sky130_fd_sc_hd__a221o_2 _18066_ (.A1(_10964_),
    .A2(_10665_),
    .B1(_10969_),
    .B2(_10965_),
    .C1(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__and4b_2 _18067_ (.A_N(_03452_),
    .B(_10916_),
    .C(_03456_),
    .D(_10018_),
    .X(_03457_));
 sky130_fd_sc_hd__buf_1 _18068_ (.A(_03457_),
    .X(_00457_));
 sky130_fd_sc_hd__and3b_2 _18069_ (.A_N(_10579_),
    .B(_10964_),
    .C(_10580_),
    .X(_03458_));
 sky130_fd_sc_hd__o41a_2 _18070_ (.A1(_10997_),
    .A2(_03458_),
    .A3(_10969_),
    .A4(_03453_),
    .B1(_10999_),
    .X(_00458_));
 sky130_fd_sc_hd__and4bb_2 _18071_ (.A_N(_10972_),
    .B_N(_10579_),
    .C(_10948_),
    .D(_10018_),
    .X(_03459_));
 sky130_fd_sc_hd__buf_1 _18072_ (.A(_03459_),
    .X(_00459_));
 sky130_fd_sc_hd__and4bb_2 _18073_ (.A_N(_10965_),
    .B_N(_10972_),
    .C(_11000_),
    .D(_10018_),
    .X(_03460_));
 sky130_fd_sc_hd__buf_1 _18074_ (.A(_03460_),
    .X(_00460_));
 sky130_fd_sc_hd__and3_2 _18075_ (.A(_10579_),
    .B(_10667_),
    .C(_10973_),
    .X(_03461_));
 sky130_fd_sc_hd__buf_1 _18076_ (.A(_03461_),
    .X(_00461_));
 sky130_fd_sc_hd__o211a_2 _18077_ (.A1(_10944_),
    .A2(_10941_),
    .B1(_10581_),
    .C1(_10946_),
    .X(_03462_));
 sky130_fd_sc_hd__o41a_2 _18078_ (.A1(_10997_),
    .A2(_10969_),
    .A3(_11034_),
    .A4(_03462_),
    .B1(_10999_),
    .X(_00462_));
 sky130_fd_sc_hd__buf_1 _18079_ (.A(_10575_),
    .X(_03463_));
 sky130_fd_sc_hd__buf_1 _18080_ (.A(_10910_),
    .X(_03464_));
 sky130_fd_sc_hd__buf_1 _18081_ (.A(_10915_),
    .X(_03465_));
 sky130_fd_sc_hd__and4bb_2 _18082_ (.A_N(_03463_),
    .B_N(_03464_),
    .C(_03465_),
    .D(\decode.io_id_pc[0] ),
    .X(_03466_));
 sky130_fd_sc_hd__buf_1 _18083_ (.A(_03466_),
    .X(_00463_));
 sky130_fd_sc_hd__buf_1 _18084_ (.A(_10910_),
    .X(_03467_));
 sky130_fd_sc_hd__and4bb_2 _18085_ (.A_N(_03463_),
    .B_N(_03467_),
    .C(_03465_),
    .D(\decode.io_id_pc[1] ),
    .X(_03468_));
 sky130_fd_sc_hd__buf_1 _18086_ (.A(_03468_),
    .X(_00464_));
 sky130_fd_sc_hd__buf_1 _18087_ (.A(_10575_),
    .X(_03469_));
 sky130_fd_sc_hd__and4bb_2 _18088_ (.A_N(_03469_),
    .B_N(_03467_),
    .C(_03465_),
    .D(\decode.io_id_pc[2] ),
    .X(_03470_));
 sky130_fd_sc_hd__buf_1 _18089_ (.A(_03470_),
    .X(_00465_));
 sky130_fd_sc_hd__and4bb_2 _18090_ (.A_N(_03469_),
    .B_N(_03467_),
    .C(_03465_),
    .D(\decode.io_id_pc[3] ),
    .X(_03471_));
 sky130_fd_sc_hd__buf_1 _18091_ (.A(_03471_),
    .X(_00466_));
 sky130_fd_sc_hd__and4bb_2 _18092_ (.A_N(_03469_),
    .B_N(_03467_),
    .C(_03465_),
    .D(\decode.io_id_pc[4] ),
    .X(_03472_));
 sky130_fd_sc_hd__buf_1 _18093_ (.A(_03472_),
    .X(_00467_));
 sky130_fd_sc_hd__and4bb_2 _18094_ (.A_N(_03469_),
    .B_N(_03467_),
    .C(_03465_),
    .D(\decode.io_id_pc[5] ),
    .X(_03473_));
 sky130_fd_sc_hd__buf_1 _18095_ (.A(_03473_),
    .X(_00468_));
 sky130_fd_sc_hd__buf_1 _18096_ (.A(_10915_),
    .X(_03474_));
 sky130_fd_sc_hd__and4bb_2 _18097_ (.A_N(_03469_),
    .B_N(_03467_),
    .C(_03474_),
    .D(\decode.io_id_pc[6] ),
    .X(_03475_));
 sky130_fd_sc_hd__buf_1 _18098_ (.A(_03475_),
    .X(_00469_));
 sky130_fd_sc_hd__and4bb_2 _18099_ (.A_N(_03469_),
    .B_N(_03467_),
    .C(_03474_),
    .D(\decode.io_id_pc[7] ),
    .X(_03476_));
 sky130_fd_sc_hd__buf_1 _18100_ (.A(_03476_),
    .X(_00470_));
 sky130_fd_sc_hd__and4bb_2 _18101_ (.A_N(_03469_),
    .B_N(_03467_),
    .C(_03474_),
    .D(\decode.io_id_pc[8] ),
    .X(_03477_));
 sky130_fd_sc_hd__buf_1 _18102_ (.A(_03477_),
    .X(_00471_));
 sky130_fd_sc_hd__and4bb_2 _18103_ (.A_N(_03469_),
    .B_N(_03467_),
    .C(_03474_),
    .D(\decode.io_id_pc[9] ),
    .X(_03478_));
 sky130_fd_sc_hd__buf_1 _18104_ (.A(_03478_),
    .X(_00472_));
 sky130_fd_sc_hd__and4bb_2 _18105_ (.A_N(_03469_),
    .B_N(_03467_),
    .C(_03474_),
    .D(\decode.io_id_pc[10] ),
    .X(_03479_));
 sky130_fd_sc_hd__buf_1 _18106_ (.A(_03479_),
    .X(_00473_));
 sky130_fd_sc_hd__buf_1 _18107_ (.A(_10909_),
    .X(_03480_));
 sky130_fd_sc_hd__and4bb_2 _18108_ (.A_N(_03469_),
    .B_N(_03480_),
    .C(_03474_),
    .D(\decode.io_id_pc[11] ),
    .X(_03481_));
 sky130_fd_sc_hd__buf_1 _18109_ (.A(_03481_),
    .X(_00474_));
 sky130_fd_sc_hd__buf_1 _18110_ (.A(_10575_),
    .X(_03482_));
 sky130_fd_sc_hd__and4bb_2 _18111_ (.A_N(_03482_),
    .B_N(_03480_),
    .C(_03474_),
    .D(\decode.io_id_pc[12] ),
    .X(_03483_));
 sky130_fd_sc_hd__buf_1 _18112_ (.A(_03483_),
    .X(_00475_));
 sky130_fd_sc_hd__and4bb_2 _18113_ (.A_N(_03482_),
    .B_N(_03480_),
    .C(_03474_),
    .D(\decode.io_id_pc[13] ),
    .X(_03484_));
 sky130_fd_sc_hd__buf_1 _18114_ (.A(_03484_),
    .X(_00476_));
 sky130_fd_sc_hd__and4bb_2 _18115_ (.A_N(_03482_),
    .B_N(_03480_),
    .C(_03474_),
    .D(\decode.io_id_pc[14] ),
    .X(_03485_));
 sky130_fd_sc_hd__buf_1 _18116_ (.A(_03485_),
    .X(_00477_));
 sky130_fd_sc_hd__and4bb_2 _18117_ (.A_N(_03482_),
    .B_N(_03480_),
    .C(_03474_),
    .D(\decode.io_id_pc[15] ),
    .X(_03486_));
 sky130_fd_sc_hd__buf_1 _18118_ (.A(_03486_),
    .X(_00478_));
 sky130_fd_sc_hd__buf_1 _18119_ (.A(_10915_),
    .X(_03487_));
 sky130_fd_sc_hd__and4bb_2 _18120_ (.A_N(_03482_),
    .B_N(_03480_),
    .C(_03487_),
    .D(\decode.io_id_pc[16] ),
    .X(_03488_));
 sky130_fd_sc_hd__buf_1 _18121_ (.A(_03488_),
    .X(_00479_));
 sky130_fd_sc_hd__and4bb_2 _18122_ (.A_N(_03482_),
    .B_N(_03480_),
    .C(_03487_),
    .D(\decode.io_id_pc[17] ),
    .X(_03489_));
 sky130_fd_sc_hd__buf_1 _18123_ (.A(_03489_),
    .X(_00480_));
 sky130_fd_sc_hd__and4bb_2 _18124_ (.A_N(_03482_),
    .B_N(_03480_),
    .C(_03487_),
    .D(\decode.io_id_pc[18] ),
    .X(_03490_));
 sky130_fd_sc_hd__buf_1 _18125_ (.A(_03490_),
    .X(_00481_));
 sky130_fd_sc_hd__and4bb_2 _18126_ (.A_N(_03482_),
    .B_N(_03480_),
    .C(_03487_),
    .D(\decode.io_id_pc[19] ),
    .X(_03491_));
 sky130_fd_sc_hd__buf_1 _18127_ (.A(_03491_),
    .X(_00482_));
 sky130_fd_sc_hd__and4bb_2 _18128_ (.A_N(_03482_),
    .B_N(_03480_),
    .C(_03487_),
    .D(\decode.io_id_pc[20] ),
    .X(_03492_));
 sky130_fd_sc_hd__buf_1 _18129_ (.A(_03492_),
    .X(_00483_));
 sky130_fd_sc_hd__buf_1 _18130_ (.A(_10909_),
    .X(_03493_));
 sky130_fd_sc_hd__and4bb_2 _18131_ (.A_N(_03482_),
    .B_N(_03493_),
    .C(_03487_),
    .D(\decode.io_id_pc[21] ),
    .X(_03494_));
 sky130_fd_sc_hd__buf_1 _18132_ (.A(_03494_),
    .X(_00484_));
 sky130_fd_sc_hd__buf_1 _18133_ (.A(_10575_),
    .X(_03495_));
 sky130_fd_sc_hd__and4bb_2 _18134_ (.A_N(_03495_),
    .B_N(_03493_),
    .C(_03487_),
    .D(\decode.io_id_pc[22] ),
    .X(_03496_));
 sky130_fd_sc_hd__buf_1 _18135_ (.A(_03496_),
    .X(_00485_));
 sky130_fd_sc_hd__and4bb_2 _18136_ (.A_N(_03495_),
    .B_N(_03493_),
    .C(_03487_),
    .D(\decode.io_id_pc[23] ),
    .X(_03497_));
 sky130_fd_sc_hd__buf_1 _18137_ (.A(_03497_),
    .X(_00486_));
 sky130_fd_sc_hd__and4bb_2 _18138_ (.A_N(_03495_),
    .B_N(_03493_),
    .C(_03487_),
    .D(\decode.io_id_pc[24] ),
    .X(_03498_));
 sky130_fd_sc_hd__buf_1 _18139_ (.A(_03498_),
    .X(_00487_));
 sky130_fd_sc_hd__and4bb_2 _18140_ (.A_N(_03495_),
    .B_N(_03493_),
    .C(_03487_),
    .D(\decode.io_id_pc[25] ),
    .X(_03499_));
 sky130_fd_sc_hd__buf_1 _18141_ (.A(_03499_),
    .X(_00488_));
 sky130_fd_sc_hd__buf_1 _18142_ (.A(_10915_),
    .X(_03500_));
 sky130_fd_sc_hd__and4bb_2 _18143_ (.A_N(_03495_),
    .B_N(_03493_),
    .C(_03500_),
    .D(\decode.io_id_pc[26] ),
    .X(_03501_));
 sky130_fd_sc_hd__buf_1 _18144_ (.A(_03501_),
    .X(_00489_));
 sky130_fd_sc_hd__and4bb_2 _18145_ (.A_N(_03495_),
    .B_N(_03493_),
    .C(_03500_),
    .D(\decode.io_id_pc[27] ),
    .X(_03502_));
 sky130_fd_sc_hd__buf_1 _18146_ (.A(_03502_),
    .X(_00490_));
 sky130_fd_sc_hd__and4bb_2 _18147_ (.A_N(_03495_),
    .B_N(_03493_),
    .C(_03500_),
    .D(\decode.io_id_pc[28] ),
    .X(_03503_));
 sky130_fd_sc_hd__buf_1 _18148_ (.A(_03503_),
    .X(_00491_));
 sky130_fd_sc_hd__and4bb_2 _18149_ (.A_N(_03495_),
    .B_N(_03493_),
    .C(_03500_),
    .D(\decode.io_id_pc[29] ),
    .X(_03504_));
 sky130_fd_sc_hd__buf_1 _18150_ (.A(_03504_),
    .X(_00492_));
 sky130_fd_sc_hd__and4bb_2 _18151_ (.A_N(_03495_),
    .B_N(_03493_),
    .C(_03500_),
    .D(\decode.io_id_pc[30] ),
    .X(_03505_));
 sky130_fd_sc_hd__buf_1 _18152_ (.A(_03505_),
    .X(_00493_));
 sky130_fd_sc_hd__and4bb_2 _18153_ (.A_N(_03495_),
    .B_N(_10910_),
    .C(_03500_),
    .D(\decode.io_id_pc[31] ),
    .X(_03506_));
 sky130_fd_sc_hd__buf_1 _18154_ (.A(_03506_),
    .X(_00494_));
 sky130_fd_sc_hd__nor4_2 _18155_ (.A(_11251_),
    .B(_10577_),
    .C(_10673_),
    .D(_10911_),
    .Y(_00495_));
 sky130_fd_sc_hd__nor4_2 _18156_ (.A(_11067_),
    .B(_10577_),
    .C(_10673_),
    .D(_10911_),
    .Y(_00496_));
 sky130_fd_sc_hd__and4bb_2 _18157_ (.A_N(_03463_),
    .B_N(_03464_),
    .C(_03465_),
    .D(_10657_),
    .X(_03507_));
 sky130_fd_sc_hd__buf_1 _18158_ (.A(_03507_),
    .X(_00497_));
 sky130_fd_sc_hd__and4bb_2 _18159_ (.A_N(_03463_),
    .B_N(_03464_),
    .C(_03465_),
    .D(_10662_),
    .X(_03508_));
 sky130_fd_sc_hd__buf_1 _18160_ (.A(_03508_),
    .X(_00498_));
 sky130_fd_sc_hd__nor4_2 _18161_ (.A(_11062_),
    .B(_10577_),
    .C(_10673_),
    .D(_10911_),
    .Y(_00499_));
 sky130_fd_sc_hd__and4bb_2 _18162_ (.A_N(_10912_),
    .B_N(_03464_),
    .C(_10921_),
    .D(\decode.control.io_funct7[0] ),
    .X(_03509_));
 sky130_fd_sc_hd__buf_1 _18163_ (.A(_03509_),
    .X(_00500_));
 sky130_fd_sc_hd__and4bb_2 _18164_ (.A_N(_03463_),
    .B_N(_03464_),
    .C(_10921_),
    .D(\decode.control.io_funct7[1] ),
    .X(_03510_));
 sky130_fd_sc_hd__buf_1 _18165_ (.A(_03510_),
    .X(_00501_));
 sky130_fd_sc_hd__and4bb_2 _18166_ (.A_N(_03463_),
    .B_N(_03464_),
    .C(_10921_),
    .D(\decode.control.io_funct7[2] ),
    .X(_03511_));
 sky130_fd_sc_hd__buf_1 _18167_ (.A(_03511_),
    .X(_00502_));
 sky130_fd_sc_hd__and4bb_2 _18168_ (.A_N(_03463_),
    .B_N(_03464_),
    .C(_10921_),
    .D(\decode.control.io_funct7[3] ),
    .X(_03512_));
 sky130_fd_sc_hd__buf_1 _18169_ (.A(_03512_),
    .X(_00503_));
 sky130_fd_sc_hd__and4bb_2 _18170_ (.A_N(_03463_),
    .B_N(_03464_),
    .C(_10921_),
    .D(\decode.control.io_funct7[4] ),
    .X(_03513_));
 sky130_fd_sc_hd__buf_1 _18171_ (.A(_03513_),
    .X(_00504_));
 sky130_fd_sc_hd__and4bb_2 _18172_ (.A_N(_03463_),
    .B_N(_03464_),
    .C(_03465_),
    .D(\decode.control.io_funct7[5] ),
    .X(_03514_));
 sky130_fd_sc_hd__buf_1 _18173_ (.A(_03514_),
    .X(_00505_));
 sky130_fd_sc_hd__and4bb_2 _18174_ (.A_N(_03463_),
    .B_N(_03464_),
    .C(_03465_),
    .D(\decode.control.io_funct7[6] ),
    .X(_03515_));
 sky130_fd_sc_hd__buf_1 _18175_ (.A(_03515_),
    .X(_00506_));
 sky130_fd_sc_hd__and3_2 _18176_ (.A(_12553_),
    .B(_12569_),
    .C(_10940_),
    .X(_03516_));
 sky130_fd_sc_hd__buf_1 _18177_ (.A(_10576_),
    .X(_03517_));
 sky130_fd_sc_hd__nand4_2 _18178_ (.A(_10579_),
    .B(\decode.control.io_opcode[5] ),
    .C(\decode.control.io_opcode[4] ),
    .D(_10580_),
    .Y(_03518_));
 sky130_fd_sc_hd__a2111oi_2 _18179_ (.A1(_10944_),
    .A2(_03516_),
    .B1(_03517_),
    .C1(_03518_),
    .D1(_10972_),
    .Y(_00507_));
 sky130_fd_sc_hd__or4_2 _18180_ (.A(\decode.immGen._imm_T_10[4] ),
    .B(\decode.immGen._imm_T_10[2] ),
    .C(\decode.immGen._imm_T_10[1] ),
    .D(\decode.immGen._imm_T_10[0] ),
    .X(_03519_));
 sky130_fd_sc_hd__or2b_2 _18181_ (.A(_10944_),
    .B_N(_10941_),
    .X(_03520_));
 sky130_fd_sc_hd__o311a_2 _18182_ (.A1(\decode.immGen._imm_T_10[3] ),
    .A2(_03519_),
    .A3(_03520_),
    .B1(_10581_),
    .C1(_11004_),
    .X(_00508_));
 sky130_fd_sc_hd__nor3_2 _18183_ (.A(\decode.control.io_funct3[2] ),
    .B(_10943_),
    .C(\decode.control.io_funct3[0] ),
    .Y(_03521_));
 sky130_fd_sc_hd__and4bb_2 _18184_ (.A_N(\decode.control.io_funct3[2] ),
    .B_N(_10944_),
    .C(_10941_),
    .D(\decode.control.io_funct7[5] ),
    .X(_03522_));
 sky130_fd_sc_hd__or4_2 _18185_ (.A(\decode.control.io_funct7[6] ),
    .B(\decode.control.io_funct7[4] ),
    .C(\decode.control.io_funct7[3] ),
    .D(\decode.control.io_funct7[1] ),
    .X(_03523_));
 sky130_fd_sc_hd__and2b_2 _18186_ (.A_N(_10943_),
    .B(\decode.control.io_funct3[0] ),
    .X(_03524_));
 sky130_fd_sc_hd__o31a_2 _18187_ (.A1(\decode.control.io_funct7[2] ),
    .A2(\decode.control.io_funct7[0] ),
    .A3(_03523_),
    .B1(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__or4b_2 _18188_ (.A(_10579_),
    .B(_10578_),
    .C(\decode.control.io_opcode[5] ),
    .D_N(\decode.control.io_opcode[4] ),
    .X(_03526_));
 sky130_fd_sc_hd__o31a_2 _18189_ (.A1(_03522_),
    .A2(_03525_),
    .A3(_03526_),
    .B1(_10582_),
    .X(_03527_));
 sky130_fd_sc_hd__and2b_2 _18190_ (.A_N(\decode.control.io_funct3[2] ),
    .B(\decode.control.io_funct3[0] ),
    .X(_03528_));
 sky130_fd_sc_hd__or3_2 _18191_ (.A(\decode.control.io_funct7[2] ),
    .B(\decode.control.io_funct7[1] ),
    .C(\decode.control.io_funct7[0] ),
    .X(_03529_));
 sky130_fd_sc_hd__or4b_2 _18192_ (.A(\decode.control.io_funct7[6] ),
    .B(_03529_),
    .C(\decode.control.io_funct7[5] ),
    .D_N(\decode.control.io_funct7[3] ),
    .X(_03530_));
 sky130_fd_sc_hd__o31a_2 _18193_ (.A1(\decode.control.io_funct7[5] ),
    .A2(\decode.control.io_funct7[2] ),
    .A3(_03523_),
    .B1(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__o22a_2 _18194_ (.A1(\decode.control.io_opcode[3] ),
    .A2(_10585_),
    .B1(_03518_),
    .B2(_03531_),
    .X(_03532_));
 sky130_fd_sc_hd__and3b_2 _18195_ (.A_N(_10946_),
    .B(_03532_),
    .C(_03526_),
    .X(_03533_));
 sky130_fd_sc_hd__o31a_2 _18196_ (.A1(_10965_),
    .A2(_10964_),
    .A3(_10951_),
    .B1(_10946_),
    .X(_03534_));
 sky130_fd_sc_hd__nor4_2 _18197_ (.A(\decode.control.io_funct7[6] ),
    .B(\decode.control.io_funct7[4] ),
    .C(\decode.control.io_funct7[3] ),
    .D(_03529_),
    .Y(_03535_));
 sky130_fd_sc_hd__o21ai_2 _18198_ (.A1(_10943_),
    .A2(_03528_),
    .B1(\decode.control.io_funct7[5] ),
    .Y(_03536_));
 sky130_fd_sc_hd__or3b_2 _18199_ (.A(_10943_),
    .B(\decode.control.io_funct3[0] ),
    .C_N(\decode.control.io_funct3[2] ),
    .X(_03537_));
 sky130_fd_sc_hd__nor2_2 _18200_ (.A(\decode.control.io_funct7[5] ),
    .B(_03523_),
    .Y(_03538_));
 sky130_fd_sc_hd__and4b_2 _18201_ (.A_N(\decode.control.io_funct7[0] ),
    .B(_03521_),
    .C(_03538_),
    .D(\decode.control.io_funct7[2] ),
    .X(_03539_));
 sky130_fd_sc_hd__a31o_2 _18202_ (.A1(_03535_),
    .A2(_03536_),
    .A3(_03537_),
    .B1(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__or2b_2 _18203_ (.A(\decode.control.io_funct3[2] ),
    .B_N(_10943_),
    .X(_03541_));
 sky130_fd_sc_hd__a21oi_2 _18204_ (.A1(_10943_),
    .A2(_10941_),
    .B1(\decode.control.io_funct3[2] ),
    .Y(_03542_));
 sky130_fd_sc_hd__a221o_2 _18205_ (.A1(_03541_),
    .A2(_10949_),
    .B1(_11000_),
    .B2(_03542_),
    .C1(_11006_),
    .X(_03543_));
 sky130_fd_sc_hd__a31oi_2 _18206_ (.A1(_03540_),
    .A2(_03458_),
    .A3(_10965_),
    .B1(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__o41a_2 _18207_ (.A1(_10944_),
    .A2(_03528_),
    .A3(_03533_),
    .A4(_03534_),
    .B1(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__o211a_2 _18208_ (.A1(_03521_),
    .A2(_03527_),
    .B1(_03545_),
    .C1(_10999_),
    .X(_00509_));
 sky130_fd_sc_hd__buf_1 _18209_ (.A(_10672_),
    .X(_03546_));
 sky130_fd_sc_hd__or3b_2 _18210_ (.A(_12494_),
    .B(_03518_),
    .C_N(_03521_),
    .X(_03547_));
 sky130_fd_sc_hd__or4_2 _18211_ (.A(\decode.immGen._imm_T_10[3] ),
    .B(_03519_),
    .C(_03530_),
    .D(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__or4b_2 _18212_ (.A(_11347_),
    .B(_03529_),
    .C(_11011_),
    .D_N(_12636_),
    .X(_03549_));
 sky130_fd_sc_hd__or4_2 _18213_ (.A(\decode.control.io_funct7[4] ),
    .B(_11100_),
    .C(_03548_),
    .D(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__buf_1 _18214_ (.A(_10910_),
    .X(_03551_));
 sky130_fd_sc_hd__nor4_2 _18215_ (.A(_10577_),
    .B(_03546_),
    .C(_03550_),
    .D(_03551_),
    .Y(_00510_));
 sky130_fd_sc_hd__nor3_2 _18216_ (.A(_11149_),
    .B(_03548_),
    .C(_03549_),
    .Y(_03552_));
 sky130_fd_sc_hd__and3_2 _18217_ (.A(\decode.control.io_funct7[4] ),
    .B(_10998_),
    .C(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__buf_1 _18218_ (.A(_03553_),
    .X(_00511_));
 sky130_fd_sc_hd__buf_1 _18219_ (.A(\csr.mcycle[19] ),
    .X(_03554_));
 sky130_fd_sc_hd__buf_1 _18220_ (.A(\csr.mcycle[22] ),
    .X(_03555_));
 sky130_fd_sc_hd__and4_2 _18221_ (.A(\csr.mcycle[14] ),
    .B(\csr.mcycle[16] ),
    .C(\csr.mcycle[15] ),
    .D(\csr.mcycle[17] ),
    .X(_03556_));
 sky130_fd_sc_hd__and3_2 _18222_ (.A(\csr.mcycle[0] ),
    .B(\csr.mcycle[2] ),
    .C(\csr.mcycle[1] ),
    .X(_03557_));
 sky130_fd_sc_hd__and4_2 _18223_ (.A(\csr.mcycle[4] ),
    .B(\csr.mcycle[3] ),
    .C(\csr.mcycle[5] ),
    .D(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__and4_2 _18224_ (.A(\csr.mcycle[6] ),
    .B(\csr.mcycle[8] ),
    .C(\csr.mcycle[7] ),
    .D(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__and3_2 _18225_ (.A(\csr.mcycle[12] ),
    .B(\csr.mcycle[11] ),
    .C(\csr.mcycle[13] ),
    .X(_03560_));
 sky130_fd_sc_hd__and4_2 _18226_ (.A(\csr.mcycle[10] ),
    .B(\csr.mcycle[9] ),
    .C(_03559_),
    .D(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__and3_2 _18227_ (.A(\csr.mcycle[18] ),
    .B(_03556_),
    .C(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__and4_2 _18228_ (.A(\csr.mcycle[20] ),
    .B(_03554_),
    .C(_03555_),
    .D(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__and4_2 _18229_ (.A(\csr.mcycle[21] ),
    .B(\csr.mcycle[24] ),
    .C(\csr.mcycle[23] ),
    .D(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__and3_2 _18230_ (.A(\csr.mcycle[28] ),
    .B(\csr.mcycle[27] ),
    .C(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__and4_2 _18231_ (.A(\csr.mcycle[26] ),
    .B(\csr.mcycle[25] ),
    .C(\csr.mcycle[30] ),
    .D(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__nand2_2 _18232_ (.A(\csr.mcycle[29] ),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__or4_2 _18233_ (.A(\csr._mcycle_T_3[63] ),
    .B(\csr._mcycle_T_3[62] ),
    .C(\csr._mcycle_T_3[61] ),
    .D(\csr._mcycle_T_3[58] ),
    .X(_03568_));
 sky130_fd_sc_hd__or4_2 _18234_ (.A(\csr._mcycle_T_3[53] ),
    .B(\csr._mcycle_T_3[52] ),
    .C(\csr._mcycle_T_3[51] ),
    .D(\csr._mcycle_T_3[50] ),
    .X(_03569_));
 sky130_fd_sc_hd__or4_2 _18235_ (.A(\csr._mcycle_T_3[57] ),
    .B(\csr._mcycle_T_3[56] ),
    .C(\csr._mcycle_T_3[55] ),
    .D(\csr._mcycle_T_3[54] ),
    .X(_03570_));
 sky130_fd_sc_hd__or4_2 _18236_ (.A(\csr._mcycle_T_3[45] ),
    .B(\csr._mcycle_T_3[44] ),
    .C(\csr._mcycle_T_3[43] ),
    .D(\csr._mcycle_T_3[42] ),
    .X(_03571_));
 sky130_fd_sc_hd__or4_2 _18237_ (.A(\csr._mcycle_T_3[49] ),
    .B(\csr._mcycle_T_3[48] ),
    .C(\csr._mcycle_T_3[47] ),
    .D(\csr._mcycle_T_3[46] ),
    .X(_03572_));
 sky130_fd_sc_hd__or4_2 _18238_ (.A(_03569_),
    .B(_03570_),
    .C(_03571_),
    .D(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__nor4_2 _18239_ (.A(\csr._mcycle_T_3[60] ),
    .B(\csr._mcycle_T_3[59] ),
    .C(_03568_),
    .D(_03573_),
    .Y(_03574_));
 sky130_fd_sc_hd__or3_2 _18240_ (.A(\csr._mcycle_T_3[33] ),
    .B(\csr._mcycle_T_3[32] ),
    .C(\csr.mcycle[31] ),
    .X(_03575_));
 sky130_fd_sc_hd__or4_2 _18241_ (.A(\csr._mcycle_T_3[37] ),
    .B(\csr._mcycle_T_3[36] ),
    .C(\csr._mcycle_T_3[35] ),
    .D(\csr._mcycle_T_3[34] ),
    .X(_03576_));
 sky130_fd_sc_hd__or4_2 _18242_ (.A(\csr._mcycle_T_3[41] ),
    .B(\csr._mcycle_T_3[40] ),
    .C(\csr._mcycle_T_3[39] ),
    .D(\csr._mcycle_T_3[38] ),
    .X(_03577_));
 sky130_fd_sc_hd__nor3_2 _18243_ (.A(_03575_),
    .B(_03576_),
    .C(_03577_),
    .Y(_03578_));
 sky130_fd_sc_hd__buf_1 _18244_ (.A(_10575_),
    .X(_03579_));
 sky130_fd_sc_hd__buf_1 _18245_ (.A(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__a31oi_2 _18246_ (.A1(_03567_),
    .A2(_03574_),
    .A3(_03578_),
    .B1(_03580_),
    .Y(_00512_));
 sky130_fd_sc_hd__buf_1 _18247_ (.A(_10910_),
    .X(_03581_));
 sky130_fd_sc_hd__buf_1 _18248_ (.A(_09954_),
    .X(_03582_));
 sky130_fd_sc_hd__buf_1 _18249_ (.A(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__and3b_2 _18250_ (.A_N(_03581_),
    .B(_03583_),
    .C(\decode.id_ex_funct3_reg[0] ),
    .X(_03584_));
 sky130_fd_sc_hd__buf_1 _18251_ (.A(_03584_),
    .X(_00513_));
 sky130_fd_sc_hd__inv_2 _18252_ (.A(\decode.id_ex_funct3_reg[1] ),
    .Y(_03585_));
 sky130_fd_sc_hd__or4_2 _18253_ (.A(reset),
    .B(_10971_),
    .C(_10757_),
    .D(_10908_),
    .X(_03586_));
 sky130_fd_sc_hd__buf_1 _18254_ (.A(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__buf_1 _18255_ (.A(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__nor2_2 _18256_ (.A(_03585_),
    .B(_03588_),
    .Y(_00514_));
 sky130_fd_sc_hd__and3b_2 _18257_ (.A_N(_03581_),
    .B(_03583_),
    .C(\decode.id_ex_funct3_reg[2] ),
    .X(_03589_));
 sky130_fd_sc_hd__buf_1 _18258_ (.A(_03589_),
    .X(_00515_));
 sky130_fd_sc_hd__nor2_2 _18259_ (.A(\csr.io_trapped ),
    .B(\csr.io_mret ),
    .Y(_03590_));
 sky130_fd_sc_hd__inv_2 _18260_ (.A(_10756_),
    .Y(_03591_));
 sky130_fd_sc_hd__buf_1 _18261_ (.A(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__o2111a_2 _18262_ (.A1(\fetch.bht.bhtTable_tag_MPORT_en ),
    .A2(_10907_),
    .B1(_03590_),
    .C1(_03592_),
    .D1(_09953_),
    .X(_03593_));
 sky130_fd_sc_hd__buf_1 _18263_ (.A(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__buf_1 _18264_ (.A(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__buf_1 _18265_ (.A(_03595_),
    .X(_03596_));
 sky130_fd_sc_hd__and2_2 _18266_ (.A(\decode.id_ex_rs2_data_reg[0] ),
    .B(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__buf_1 _18267_ (.A(_03597_),
    .X(_00516_));
 sky130_fd_sc_hd__inv_2 _18268_ (.A(\decode.id_ex_rs2_data_reg[1] ),
    .Y(_03598_));
 sky130_fd_sc_hd__buf_1 _18269_ (.A(_03588_),
    .X(_03599_));
 sky130_fd_sc_hd__nor2_2 _18270_ (.A(_03598_),
    .B(_03599_),
    .Y(_00517_));
 sky130_fd_sc_hd__and2_2 _18271_ (.A(\decode.id_ex_rs2_data_reg[2] ),
    .B(_03596_),
    .X(_03600_));
 sky130_fd_sc_hd__buf_1 _18272_ (.A(_03600_),
    .X(_00518_));
 sky130_fd_sc_hd__and2_2 _18273_ (.A(\decode.id_ex_rs2_data_reg[3] ),
    .B(_03596_),
    .X(_03601_));
 sky130_fd_sc_hd__buf_1 _18274_ (.A(_03601_),
    .X(_00519_));
 sky130_fd_sc_hd__and2_2 _18275_ (.A(\decode.id_ex_rs2_data_reg[4] ),
    .B(_03596_),
    .X(_03602_));
 sky130_fd_sc_hd__buf_1 _18276_ (.A(_03602_),
    .X(_00520_));
 sky130_fd_sc_hd__and2_2 _18277_ (.A(\decode.id_ex_rs2_data_reg[5] ),
    .B(_03596_),
    .X(_03603_));
 sky130_fd_sc_hd__buf_1 _18278_ (.A(_03603_),
    .X(_00521_));
 sky130_fd_sc_hd__and2_2 _18279_ (.A(\decode.id_ex_rs2_data_reg[6] ),
    .B(_03596_),
    .X(_03604_));
 sky130_fd_sc_hd__buf_1 _18280_ (.A(_03604_),
    .X(_00522_));
 sky130_fd_sc_hd__buf_1 _18281_ (.A(_03595_),
    .X(_03605_));
 sky130_fd_sc_hd__and2_2 _18282_ (.A(\decode.id_ex_rs2_data_reg[7] ),
    .B(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__buf_1 _18283_ (.A(_03606_),
    .X(_00523_));
 sky130_fd_sc_hd__and2_2 _18284_ (.A(\decode.id_ex_rs2_data_reg[8] ),
    .B(_03605_),
    .X(_03607_));
 sky130_fd_sc_hd__buf_1 _18285_ (.A(_03607_),
    .X(_00524_));
 sky130_fd_sc_hd__and2_2 _18286_ (.A(\decode.id_ex_rs2_data_reg[9] ),
    .B(_03605_),
    .X(_03608_));
 sky130_fd_sc_hd__buf_1 _18287_ (.A(_03608_),
    .X(_00525_));
 sky130_fd_sc_hd__and2_2 _18288_ (.A(\decode.id_ex_rs2_data_reg[10] ),
    .B(_03605_),
    .X(_03609_));
 sky130_fd_sc_hd__buf_1 _18289_ (.A(_03609_),
    .X(_00526_));
 sky130_fd_sc_hd__and2_2 _18290_ (.A(\decode.id_ex_rs2_data_reg[11] ),
    .B(_03605_),
    .X(_03610_));
 sky130_fd_sc_hd__buf_1 _18291_ (.A(_03610_),
    .X(_00527_));
 sky130_fd_sc_hd__and2_2 _18292_ (.A(\decode.id_ex_rs2_data_reg[12] ),
    .B(_03605_),
    .X(_03611_));
 sky130_fd_sc_hd__buf_1 _18293_ (.A(_03611_),
    .X(_00528_));
 sky130_fd_sc_hd__and2_2 _18294_ (.A(\decode.id_ex_rs2_data_reg[13] ),
    .B(_03605_),
    .X(_03612_));
 sky130_fd_sc_hd__buf_1 _18295_ (.A(_03612_),
    .X(_00529_));
 sky130_fd_sc_hd__and2_2 _18296_ (.A(\decode.id_ex_rs2_data_reg[14] ),
    .B(_03605_),
    .X(_03613_));
 sky130_fd_sc_hd__buf_1 _18297_ (.A(_03613_),
    .X(_00530_));
 sky130_fd_sc_hd__and2_2 _18298_ (.A(\decode.id_ex_rs2_data_reg[15] ),
    .B(_03605_),
    .X(_03614_));
 sky130_fd_sc_hd__buf_1 _18299_ (.A(_03614_),
    .X(_00531_));
 sky130_fd_sc_hd__and2_2 _18300_ (.A(\decode.id_ex_rs2_data_reg[16] ),
    .B(_03605_),
    .X(_03615_));
 sky130_fd_sc_hd__buf_1 _18301_ (.A(_03615_),
    .X(_00532_));
 sky130_fd_sc_hd__buf_1 _18302_ (.A(_03595_),
    .X(_03616_));
 sky130_fd_sc_hd__and2_2 _18303_ (.A(\decode.id_ex_rs2_data_reg[17] ),
    .B(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__buf_1 _18304_ (.A(_03617_),
    .X(_00533_));
 sky130_fd_sc_hd__and2_2 _18305_ (.A(\decode.id_ex_rs2_data_reg[18] ),
    .B(_03616_),
    .X(_03618_));
 sky130_fd_sc_hd__buf_1 _18306_ (.A(_03618_),
    .X(_00534_));
 sky130_fd_sc_hd__and2_2 _18307_ (.A(\decode.id_ex_rs2_data_reg[19] ),
    .B(_03616_),
    .X(_03619_));
 sky130_fd_sc_hd__buf_1 _18308_ (.A(_03619_),
    .X(_00535_));
 sky130_fd_sc_hd__and2_2 _18309_ (.A(\decode.id_ex_rs2_data_reg[20] ),
    .B(_03616_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_1 _18310_ (.A(_03620_),
    .X(_00536_));
 sky130_fd_sc_hd__and2_2 _18311_ (.A(\decode.id_ex_rs2_data_reg[21] ),
    .B(_03616_),
    .X(_03621_));
 sky130_fd_sc_hd__buf_1 _18312_ (.A(_03621_),
    .X(_00537_));
 sky130_fd_sc_hd__and2_2 _18313_ (.A(\decode.id_ex_rs2_data_reg[22] ),
    .B(_03616_),
    .X(_03622_));
 sky130_fd_sc_hd__buf_1 _18314_ (.A(_03622_),
    .X(_00538_));
 sky130_fd_sc_hd__and2_2 _18315_ (.A(\decode.id_ex_rs2_data_reg[23] ),
    .B(_03616_),
    .X(_03623_));
 sky130_fd_sc_hd__buf_1 _18316_ (.A(_03623_),
    .X(_00539_));
 sky130_fd_sc_hd__and2_2 _18317_ (.A(\decode.id_ex_rs2_data_reg[24] ),
    .B(_03616_),
    .X(_03624_));
 sky130_fd_sc_hd__buf_1 _18318_ (.A(_03624_),
    .X(_00540_));
 sky130_fd_sc_hd__and2_2 _18319_ (.A(\decode.id_ex_rs2_data_reg[25] ),
    .B(_03616_),
    .X(_03625_));
 sky130_fd_sc_hd__buf_1 _18320_ (.A(_03625_),
    .X(_00541_));
 sky130_fd_sc_hd__and2_2 _18321_ (.A(\decode.id_ex_rs2_data_reg[26] ),
    .B(_03616_),
    .X(_03626_));
 sky130_fd_sc_hd__buf_1 _18322_ (.A(_03626_),
    .X(_00542_));
 sky130_fd_sc_hd__buf_1 _18323_ (.A(_03594_),
    .X(_03627_));
 sky130_fd_sc_hd__and2_2 _18324_ (.A(\decode.id_ex_rs2_data_reg[27] ),
    .B(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__buf_1 _18325_ (.A(_03628_),
    .X(_00543_));
 sky130_fd_sc_hd__and2_2 _18326_ (.A(\decode.id_ex_rs2_data_reg[28] ),
    .B(_03627_),
    .X(_03629_));
 sky130_fd_sc_hd__buf_1 _18327_ (.A(_03629_),
    .X(_00544_));
 sky130_fd_sc_hd__and2_2 _18328_ (.A(\decode.id_ex_rs2_data_reg[29] ),
    .B(_03627_),
    .X(_03630_));
 sky130_fd_sc_hd__buf_1 _18329_ (.A(_03630_),
    .X(_00545_));
 sky130_fd_sc_hd__and2_2 _18330_ (.A(\decode.id_ex_rs2_data_reg[30] ),
    .B(_03627_),
    .X(_03631_));
 sky130_fd_sc_hd__buf_1 _18331_ (.A(_03631_),
    .X(_00546_));
 sky130_fd_sc_hd__and2_2 _18332_ (.A(\decode.id_ex_rs2_data_reg[31] ),
    .B(_03627_),
    .X(_03632_));
 sky130_fd_sc_hd__buf_1 _18333_ (.A(_03632_),
    .X(_00547_));
 sky130_fd_sc_hd__buf_1 _18334_ (.A(\decode.id_ex_aluop_reg[1] ),
    .X(_03633_));
 sky130_fd_sc_hd__buf_1 _18335_ (.A(\decode.id_ex_aluop_reg[2] ),
    .X(_03634_));
 sky130_fd_sc_hd__buf_1 _18336_ (.A(\decode.id_ex_aluop_reg[3] ),
    .X(_03635_));
 sky130_fd_sc_hd__or3b_2 _18337_ (.A(_03633_),
    .B(_03634_),
    .C_N(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__buf_1 _18338_ (.A(\decode.id_ex_aluop_reg[0] ),
    .X(_03637_));
 sky130_fd_sc_hd__buf_1 _18339_ (.A(_03637_),
    .X(_03638_));
 sky130_fd_sc_hd__buf_1 _18340_ (.A(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__inv_2 _18341_ (.A(\execute.io_mem_rd[3] ),
    .Y(_03640_));
 sky130_fd_sc_hd__nand2_2 _18342_ (.A(_03640_),
    .B(\decode.id_ex_ex_rs1_reg[3] ),
    .Y(_03641_));
 sky130_fd_sc_hd__inv_2 _18343_ (.A(\execute.io_mem_rd[0] ),
    .Y(_03642_));
 sky130_fd_sc_hd__nand2_2 _18344_ (.A(_03642_),
    .B(\decode.id_ex_ex_rs1_reg[0] ),
    .Y(_03643_));
 sky130_fd_sc_hd__and3_2 _18345_ (.A(_09921_),
    .B(_03641_),
    .C(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__or2b_2 _18346_ (.A(\execute.io_mem_rd[2] ),
    .B_N(\decode.id_ex_ex_rs1_reg[2] ),
    .X(_03645_));
 sky130_fd_sc_hd__or2b_2 _18347_ (.A(\decode.id_ex_ex_rs1_reg[2] ),
    .B_N(\execute.io_mem_rd[2] ),
    .X(_03646_));
 sky130_fd_sc_hd__or2b_2 _18348_ (.A(\decode.id_ex_ex_rs1_reg[1] ),
    .B_N(\execute.io_mem_rd[1] ),
    .X(_03647_));
 sky130_fd_sc_hd__or2b_2 _18349_ (.A(\execute.io_mem_rd[1] ),
    .B_N(\decode.id_ex_ex_rs1_reg[1] ),
    .X(_03648_));
 sky130_fd_sc_hd__o2111a_2 _18350_ (.A1(_03642_),
    .A2(\decode.id_ex_ex_rs1_reg[0] ),
    .B1(_03646_),
    .C1(_03647_),
    .D1(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__and2_2 _18351_ (.A(\execute.io_mem_regwrite ),
    .B(\decode.id_ex_ex_use_rs1_reg ),
    .X(_03650_));
 sky130_fd_sc_hd__nand2_2 _18352_ (.A(_09920_),
    .B(\decode.id_ex_ex_rs1_reg[4] ),
    .Y(_03651_));
 sky130_fd_sc_hd__inv_2 _18353_ (.A(\decode.id_ex_ex_rs1_reg[4] ),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2_2 _18354_ (.A(_03652_),
    .B(\execute.io_mem_rd[4] ),
    .Y(_03653_));
 sky130_fd_sc_hd__o2111a_2 _18355_ (.A1(_03640_),
    .A2(\decode.id_ex_ex_rs1_reg[3] ),
    .B1(_03650_),
    .C1(_03651_),
    .D1(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__nand4_2 _18356_ (.A(_03644_),
    .B(_03645_),
    .C(_03649_),
    .D(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__buf_1 _18357_ (.A(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__nand2_2 _18358_ (.A(\execute.io_mem_memtoreg[1] ),
    .B(\execute.io_mem_memtoreg[0] ),
    .Y(_03657_));
 sky130_fd_sc_hd__buf_1 _18359_ (.A(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_1 _18360_ (.A(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__inv_2 _18361_ (.A(\execute.io_mem_memtoreg[1] ),
    .Y(_03660_));
 sky130_fd_sc_hd__inv_2 _18362_ (.A(\execute.io_mem_memtoreg[0] ),
    .Y(_03661_));
 sky130_fd_sc_hd__nand2_2 _18363_ (.A(_03660_),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__nand2_2 _18364_ (.A(_03657_),
    .B(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__buf_1 _18365_ (.A(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__buf_1 _18366_ (.A(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__buf_1 _18367_ (.A(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__o22a_2 _18368_ (.A1(\execute.csr_read_data_out_reg[31] ),
    .A2(_03659_),
    .B1(io_memory_address[31]),
    .B2(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__o31a_2 _18369_ (.A1(\execute.io_mem_memtoreg[1] ),
    .A2(\execute.io_mem_memtoreg[0] ),
    .A3(\execute.io_reg_pc[31] ),
    .B1(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__inv_2 _18370_ (.A(\decode.id_ex_islui_reg ),
    .Y(_03669_));
 sky130_fd_sc_hd__buf_1 _18371_ (.A(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__or2b_2 _18372_ (.A(_09929_),
    .B_N(\decode.id_ex_ex_rs1_reg[2] ),
    .X(_03671_));
 sky130_fd_sc_hd__nor2_2 _18373_ (.A(\decode.io_wb_rd[2] ),
    .B(\decode.io_wb_rd[3] ),
    .Y(_03672_));
 sky130_fd_sc_hd__nand3b_2 _18374_ (.A_N(\decode.io_wb_rd[4] ),
    .B(_10196_),
    .C(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__o22a_2 _18375_ (.A1(\decode.io_wb_rd[4] ),
    .A2(_03652_),
    .B1(\decode.id_ex_ex_rs1_reg[1] ),
    .B2(_09931_),
    .X(_03674_));
 sky130_fd_sc_hd__o2111ai_2 _18376_ (.A1(_09935_),
    .A2(\decode.id_ex_ex_rs1_reg[3] ),
    .B1(_03671_),
    .C1(_03673_),
    .D1(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__nand2_2 _18377_ (.A(_09934_),
    .B(\decode.id_ex_ex_rs1_reg[3] ),
    .Y(_03676_));
 sky130_fd_sc_hd__or2b_2 _18378_ (.A(\decode.io_wb_rd[1] ),
    .B_N(\decode.id_ex_ex_rs1_reg[1] ),
    .X(_03677_));
 sky130_fd_sc_hd__or2b_2 _18379_ (.A(\decode.io_wb_rd[0] ),
    .B_N(\decode.id_ex_ex_rs1_reg[0] ),
    .X(_03678_));
 sky130_fd_sc_hd__nand3_2 _18380_ (.A(_03676_),
    .B(_03677_),
    .C(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__inv_2 _18381_ (.A(\decode.id_ex_ex_rs1_reg[2] ),
    .Y(_03680_));
 sky130_fd_sc_hd__nand2_2 _18382_ (.A(\decode.io_wb_regwrite ),
    .B(\decode.id_ex_ex_use_rs1_reg ),
    .Y(_03681_));
 sky130_fd_sc_hd__a21oi_2 _18383_ (.A1(_03680_),
    .A2(_09929_),
    .B1(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__or2b_2 _18384_ (.A(\decode.id_ex_ex_rs1_reg[0] ),
    .B_N(\decode.io_wb_rd[0] ),
    .X(_03683_));
 sky130_fd_sc_hd__nand2_2 _18385_ (.A(_03652_),
    .B(\decode.io_wb_rd[4] ),
    .Y(_03684_));
 sky130_fd_sc_hd__nand4b_2 _18386_ (.A_N(_03679_),
    .B(_03682_),
    .C(_03683_),
    .D(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__o21ai_2 _18387_ (.A1(_03675_),
    .A2(_03685_),
    .B1(_03655_),
    .Y(_03686_));
 sky130_fd_sc_hd__buf_1 _18388_ (.A(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__buf_1 _18389_ (.A(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__buf_1 _18390_ (.A(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__o22a_2 _18391_ (.A1(\memory.csr_read_data_out_reg[31] ),
    .A2(_09988_),
    .B1(_10144_),
    .B2(_10145_),
    .X(_03690_));
 sky130_fd_sc_hd__or2b_2 _18392_ (.A(\decode.io_wb_rd[4] ),
    .B_N(\decode.id_ex_ex_rs1_reg[4] ),
    .X(_03691_));
 sky130_fd_sc_hd__or2b_2 _18393_ (.A(\decode.id_ex_ex_rs1_reg[1] ),
    .B_N(\decode.io_wb_rd[1] ),
    .X(_03692_));
 sky130_fd_sc_hd__nand4_2 _18394_ (.A(_03691_),
    .B(_03692_),
    .C(_03683_),
    .D(_03671_),
    .Y(_03693_));
 sky130_fd_sc_hd__or2b_2 _18395_ (.A(\decode.id_ex_ex_rs1_reg[3] ),
    .B_N(_10194_),
    .X(_03694_));
 sky130_fd_sc_hd__nand4b_2 _18396_ (.A_N(_03681_),
    .B(_03676_),
    .C(_03694_),
    .D(_03677_),
    .Y(_03695_));
 sky130_fd_sc_hd__a22oi_2 _18397_ (.A1(_03680_),
    .A2(_09929_),
    .B1(\decode.io_wb_rd[4] ),
    .B2(_03652_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand3_2 _18398_ (.A(_03696_),
    .B(_03678_),
    .C(_03673_),
    .Y(_03697_));
 sky130_fd_sc_hd__nor3_2 _18399_ (.A(_03693_),
    .B(_03695_),
    .C(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__nand2_2 _18400_ (.A(_03655_),
    .B(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__buf_1 _18401_ (.A(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__buf_1 _18402_ (.A(_03700_),
    .X(_03701_));
 sky130_fd_sc_hd__o22a_2 _18403_ (.A1(\decode.id_ex_rs1_data_reg[31] ),
    .A2(_03689_),
    .B1(_03690_),
    .B2(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__o211a_2 _18404_ (.A1(_03656_),
    .A2(_03668_),
    .B1(_03670_),
    .C1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__buf_1 _18405_ (.A(_03703_),
    .X(_03704_));
 sky130_fd_sc_hd__buf_1 _18406_ (.A(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__buf_1 _18407_ (.A(\decode.id_ex_immsrc_reg ),
    .X(_03706_));
 sky130_fd_sc_hd__buf_1 _18408_ (.A(_03706_),
    .X(_03707_));
 sky130_fd_sc_hd__buf_1 _18409_ (.A(_03707_),
    .X(_03708_));
 sky130_fd_sc_hd__buf_1 _18410_ (.A(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__buf_1 _18411_ (.A(\csr.io_csr_address[1] ),
    .X(_03710_));
 sky130_fd_sc_hd__nor2_2 _18412_ (.A(\execute.io_mem_rd[1] ),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__and2_2 _18413_ (.A(\execute.io_mem_rd[1] ),
    .B(_03710_),
    .X(_03712_));
 sky130_fd_sc_hd__nand2_2 _18414_ (.A(_03640_),
    .B(\csr.io_csr_address[3] ),
    .Y(_03713_));
 sky130_fd_sc_hd__o211ai_2 _18415_ (.A1(_03711_),
    .A2(_03712_),
    .B1(_09921_),
    .C1(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__buf_1 _18416_ (.A(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__xnor2_2 _18417_ (.A(\execute.io_mem_rd[2] ),
    .B(\csr.io_csr_address[2] ),
    .Y(_03716_));
 sky130_fd_sc_hd__xnor2_2 _18418_ (.A(\execute.io_mem_rd[4] ),
    .B(\csr.io_csr_address[4] ),
    .Y(_03717_));
 sky130_fd_sc_hd__buf_1 _18419_ (.A(\csr.io_csr_address[0] ),
    .X(_03718_));
 sky130_fd_sc_hd__inv_2 _18420_ (.A(\csr.io_csr_address[3] ),
    .Y(_03719_));
 sky130_fd_sc_hd__a22oi_2 _18421_ (.A1(_03642_),
    .A2(_03718_),
    .B1(\execute.io_mem_rd[3] ),
    .B2(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__inv_2 _18422_ (.A(\csr.io_csr_address[0] ),
    .Y(_03721_));
 sky130_fd_sc_hd__nand2_2 _18423_ (.A(\decode.id_ex_ex_use_rs2_reg ),
    .B(\execute.io_mem_regwrite ),
    .Y(_03722_));
 sky130_fd_sc_hd__a21oi_2 _18424_ (.A1(_03721_),
    .A2(\execute.io_mem_rd[0] ),
    .B1(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__nand4_2 _18425_ (.A(_03716_),
    .B(_03717_),
    .C(_03720_),
    .D(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__buf_1 _18426_ (.A(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__inv_2 _18427_ (.A(\decode.id_ex_immsrc_reg ),
    .Y(_03726_));
 sky130_fd_sc_hd__buf_1 _18428_ (.A(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__buf_1 _18429_ (.A(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__o31a_2 _18430_ (.A1(_03715_),
    .A2(_03725_),
    .A3(_03668_),
    .B1(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__or2b_2 _18431_ (.A(\decode.io_wb_rd[4] ),
    .B_N(\csr.io_csr_address[4] ),
    .X(_03730_));
 sky130_fd_sc_hd__or2b_2 _18432_ (.A(\decode.io_wb_rd[0] ),
    .B_N(\csr.io_csr_address[0] ),
    .X(_03731_));
 sky130_fd_sc_hd__or2b_2 _18433_ (.A(\csr.io_csr_address[4] ),
    .B_N(\decode.io_wb_rd[4] ),
    .X(_03732_));
 sky130_fd_sc_hd__or2b_2 _18434_ (.A(\csr.io_csr_address[0] ),
    .B_N(\decode.io_wb_rd[0] ),
    .X(_03733_));
 sky130_fd_sc_hd__nand4_2 _18435_ (.A(_03730_),
    .B(_03731_),
    .C(_03732_),
    .D(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__and2_2 _18436_ (.A(\decode.io_wb_regwrite ),
    .B(\decode.id_ex_ex_use_rs2_reg ),
    .X(_03735_));
 sky130_fd_sc_hd__or2b_2 _18437_ (.A(\decode.io_wb_rd[1] ),
    .B_N(_03710_),
    .X(_03736_));
 sky130_fd_sc_hd__inv_2 _18438_ (.A(\csr.io_csr_address[1] ),
    .Y(_03737_));
 sky130_fd_sc_hd__nand2_2 _18439_ (.A(_03737_),
    .B(\decode.io_wb_rd[1] ),
    .Y(_03738_));
 sky130_fd_sc_hd__o2111a_2 _18440_ (.A1(\decode.io_wb_rd[3] ),
    .A2(_03719_),
    .B1(_03735_),
    .C1(_03736_),
    .D1(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__or2b_2 _18441_ (.A(\decode.io_wb_rd[2] ),
    .B_N(\csr.io_csr_address[2] ),
    .X(_03740_));
 sky130_fd_sc_hd__inv_2 _18442_ (.A(\csr.io_csr_address[2] ),
    .Y(_03741_));
 sky130_fd_sc_hd__nand2_2 _18443_ (.A(_03741_),
    .B(\decode.io_wb_rd[2] ),
    .Y(_03742_));
 sky130_fd_sc_hd__o211a_2 _18444_ (.A1(_09934_),
    .A2(\csr.io_csr_address[3] ),
    .B1(_03740_),
    .C1(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__nand4b_2 _18445_ (.A_N(_03734_),
    .B(_03739_),
    .C(_03743_),
    .D(_03673_),
    .Y(_03744_));
 sky130_fd_sc_hd__o21ai_2 _18446_ (.A1(_03714_),
    .A2(_03724_),
    .B1(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__buf_1 _18447_ (.A(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__buf_1 _18448_ (.A(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__and2_2 _18449_ (.A(\decode.id_ex_ex_use_rs2_reg ),
    .B(\execute.io_mem_regwrite ),
    .X(_03748_));
 sky130_fd_sc_hd__or2b_2 _18450_ (.A(\execute.io_mem_rd[2] ),
    .B_N(\csr.io_csr_address[2] ),
    .X(_03749_));
 sky130_fd_sc_hd__nand2_2 _18451_ (.A(_03741_),
    .B(\execute.io_mem_rd[2] ),
    .Y(_03750_));
 sky130_fd_sc_hd__o2111a_2 _18452_ (.A1(_03718_),
    .A2(_03642_),
    .B1(_03748_),
    .C1(_03749_),
    .D1(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__o211a_2 _18453_ (.A1(_03711_),
    .A2(_03712_),
    .B1(_09921_),
    .C1(_03713_),
    .X(_03752_));
 sky130_fd_sc_hd__nand2_2 _18454_ (.A(\execute.io_mem_rd[4] ),
    .B(\csr.io_csr_address[4] ),
    .Y(_03753_));
 sky130_fd_sc_hd__or2_2 _18455_ (.A(\execute.io_mem_rd[4] ),
    .B(\csr.io_csr_address[4] ),
    .X(_03754_));
 sky130_fd_sc_hd__buf_1 _18456_ (.A(_03719_),
    .X(_03755_));
 sky130_fd_sc_hd__o2bb2ai_2 _18457_ (.A1_N(\execute.io_mem_rd[3] ),
    .A2_N(_03755_),
    .B1(\execute.io_mem_rd[0] ),
    .B2(_03721_),
    .Y(_03756_));
 sky130_fd_sc_hd__a21oi_2 _18458_ (.A1(_03753_),
    .A2(_03754_),
    .B1(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__nand3_2 _18459_ (.A(_03751_),
    .B(_03752_),
    .C(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__buf_1 _18460_ (.A(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__and4_2 _18461_ (.A(_03673_),
    .B(_03732_),
    .C(_03733_),
    .D(_03742_),
    .X(_03760_));
 sky130_fd_sc_hd__nand2_2 _18462_ (.A(_03719_),
    .B(\decode.io_wb_rd[3] ),
    .Y(_03761_));
 sky130_fd_sc_hd__and4_2 _18463_ (.A(_03730_),
    .B(_03731_),
    .C(_03740_),
    .D(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__nand4_2 _18464_ (.A(_03759_),
    .B(_03739_),
    .C(_03760_),
    .D(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__buf_1 _18465_ (.A(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__o22a_2 _18466_ (.A1(\decode.id_ex_rs2_data_reg[31] ),
    .A2(_03747_),
    .B1(_03690_),
    .B2(_03764_),
    .X(_03765_));
 sky130_fd_sc_hd__a22oi_2 _18467_ (.A1(_03709_),
    .A2(\decode.id_ex_imm_reg[31] ),
    .B1(_03729_),
    .B2(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__and3_2 _18468_ (.A(_03639_),
    .B(_03705_),
    .C(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__o2111ai_2 _18469_ (.A1(\decode.id_ex_ex_rs1_reg[0] ),
    .A2(_03642_),
    .B1(_03647_),
    .C1(_03646_),
    .D1(_03648_),
    .Y(_03768_));
 sky130_fd_sc_hd__nand4_2 _18470_ (.A(_09921_),
    .B(_03645_),
    .C(_03641_),
    .D(_03643_),
    .Y(_03769_));
 sky130_fd_sc_hd__o2111ai_2 _18471_ (.A1(\decode.id_ex_ex_rs1_reg[3] ),
    .A2(_03640_),
    .B1(_03650_),
    .C1(_03653_),
    .D1(_03651_),
    .Y(_03770_));
 sky130_fd_sc_hd__o31a_2 _18472_ (.A1(_03768_),
    .A2(_03769_),
    .A3(_03770_),
    .B1(_03698_),
    .X(_03771_));
 sky130_fd_sc_hd__buf_1 _18473_ (.A(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__buf_1 _18474_ (.A(\decode.id_ex_islui_reg ),
    .X(_03773_));
 sky130_fd_sc_hd__buf_1 _18475_ (.A(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__buf_1 _18476_ (.A(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__buf_1 _18477_ (.A(_03662_),
    .X(_03776_));
 sky130_fd_sc_hd__buf_1 _18478_ (.A(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__or3_2 _18479_ (.A(\execute.csr_read_data_out_reg[29] ),
    .B(_03661_),
    .C(_03660_),
    .X(_03778_));
 sky130_fd_sc_hd__o221a_2 _18480_ (.A1(\execute.io_reg_pc[29] ),
    .A2(_03777_),
    .B1(_03666_),
    .B2(io_memory_address[29]),
    .C1(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__o22ai_2 _18481_ (.A1(_03656_),
    .A2(_03779_),
    .B1(\decode.id_ex_rs1_data_reg[29] ),
    .B2(_03689_),
    .Y(_03780_));
 sky130_fd_sc_hd__a211oi_2 _18482_ (.A1(_10135_),
    .A2(_03772_),
    .B1(_03775_),
    .C1(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__o2111ai_2 _18483_ (.A1(_10194_),
    .A2(_03755_),
    .B1(_03735_),
    .C1(_03736_),
    .D1(_03738_),
    .Y(_03782_));
 sky130_fd_sc_hd__nand4_2 _18484_ (.A(_03673_),
    .B(_03740_),
    .C(_03761_),
    .D(_03742_),
    .Y(_03783_));
 sky130_fd_sc_hd__nor3_2 _18485_ (.A(_03734_),
    .B(_03782_),
    .C(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__o21a_2 _18486_ (.A1(_03715_),
    .A2(_03725_),
    .B1(_03784_),
    .X(_03785_));
 sky130_fd_sc_hd__o221a_2 _18487_ (.A1(_03759_),
    .A2(_03779_),
    .B1(\decode.id_ex_rs2_data_reg[29] ),
    .B2(_03747_),
    .C1(_03727_),
    .X(_03786_));
 sky130_fd_sc_hd__a21boi_2 _18488_ (.A1(_10135_),
    .A2(_03785_),
    .B1_N(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__a21oi_2 _18489_ (.A1(_03709_),
    .A2(\decode.id_ex_imm_reg[29] ),
    .B1(_03787_),
    .Y(_03788_));
 sky130_fd_sc_hd__nor2_2 _18490_ (.A(_03781_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__and2_2 _18491_ (.A(_03781_),
    .B(_03788_),
    .X(_03790_));
 sky130_fd_sc_hd__or2_2 _18492_ (.A(_03789_),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__or3_2 _18493_ (.A(\execute.csr_read_data_out_reg[28] ),
    .B(_03661_),
    .C(_03660_),
    .X(_03792_));
 sky130_fd_sc_hd__o221a_2 _18494_ (.A1(\execute.io_reg_pc[28] ),
    .A2(_03777_),
    .B1(_03666_),
    .B2(io_memory_address[28]),
    .C1(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__o22ai_2 _18495_ (.A1(_03656_),
    .A2(_03793_),
    .B1(\decode.id_ex_rs1_data_reg[28] ),
    .B2(_03689_),
    .Y(_03794_));
 sky130_fd_sc_hd__a211oi_2 _18496_ (.A1(_10127_),
    .A2(_03772_),
    .B1(_03775_),
    .C1(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__nor2_2 _18497_ (.A(_03714_),
    .B(_03724_),
    .Y(_03796_));
 sky130_fd_sc_hd__buf_1 _18498_ (.A(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__or3b_2 _18499_ (.A(_03744_),
    .B(_03797_),
    .C_N(_10127_),
    .X(_03798_));
 sky130_fd_sc_hd__o221a_2 _18500_ (.A1(_03759_),
    .A2(_03793_),
    .B1(\decode.id_ex_rs2_data_reg[28] ),
    .B2(_03747_),
    .C1(_03728_),
    .X(_03799_));
 sky130_fd_sc_hd__a22oi_2 _18501_ (.A1(_03709_),
    .A2(\decode.id_ex_imm_reg[28] ),
    .B1(_03798_),
    .B2(_03799_),
    .Y(_03800_));
 sky130_fd_sc_hd__or2_2 _18502_ (.A(_03795_),
    .B(_03800_),
    .X(_03801_));
 sky130_fd_sc_hd__nand2_2 _18503_ (.A(_03795_),
    .B(_03800_),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_2 _18504_ (.A(_03801_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__o22a_2 _18505_ (.A1(\execute.csr_read_data_out_reg[26] ),
    .A2(_03659_),
    .B1(io_memory_address[26]),
    .B2(_03666_),
    .X(_03804_));
 sky130_fd_sc_hd__o31a_2 _18506_ (.A1(\execute.io_mem_memtoreg[1] ),
    .A2(\execute.io_mem_memtoreg[0] ),
    .A3(\execute.io_reg_pc[26] ),
    .B1(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__o22ai_2 _18507_ (.A1(_03656_),
    .A2(_03805_),
    .B1(\decode.id_ex_rs1_data_reg[26] ),
    .B2(_03689_),
    .Y(_03806_));
 sky130_fd_sc_hd__or3b_2 _18508_ (.A(_03744_),
    .B(_03797_),
    .C_N(_10116_),
    .X(_03807_));
 sky130_fd_sc_hd__o221a_2 _18509_ (.A1(\decode.id_ex_rs2_data_reg[26] ),
    .A2(_03747_),
    .B1(_03805_),
    .B2(_03759_),
    .C1(_03727_),
    .X(_03808_));
 sky130_fd_sc_hd__a22oi_2 _18510_ (.A1(_03709_),
    .A2(\decode.id_ex_imm_reg[26] ),
    .B1(_03807_),
    .B2(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__inv_2 _18511_ (.A(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__a2111o_2 _18512_ (.A1(_10116_),
    .A2(_03772_),
    .B1(_03775_),
    .C1(_03806_),
    .D1(_03810_),
    .X(_03811_));
 sky130_fd_sc_hd__a211oi_2 _18513_ (.A1(_10116_),
    .A2(_03772_),
    .B1(_03775_),
    .C1(_03806_),
    .Y(_03812_));
 sky130_fd_sc_hd__or2_2 _18514_ (.A(_03812_),
    .B(_03809_),
    .X(_03813_));
 sky130_fd_sc_hd__nand2_2 _18515_ (.A(_03811_),
    .B(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__nor3_2 _18516_ (.A(_03768_),
    .B(_03769_),
    .C(_03770_),
    .Y(_03815_));
 sky130_fd_sc_hd__buf_1 _18517_ (.A(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__buf_1 _18518_ (.A(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__o22a_2 _18519_ (.A1(_03659_),
    .A2(\execute.csr_read_data_out_reg[27] ),
    .B1(\execute.io_reg_pc[27] ),
    .B2(_03777_),
    .X(_03818_));
 sky130_fd_sc_hd__o21ai_2 _18520_ (.A1(io_memory_address[27]),
    .A2(_03666_),
    .B1(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__a2bb2o_2 _18521_ (.A1_N(\decode.id_ex_rs1_data_reg[27] ),
    .A2_N(_03689_),
    .B1(_10121_),
    .B2(_03772_),
    .X(_03820_));
 sky130_fd_sc_hd__a211oi_2 _18522_ (.A1(_03817_),
    .A2(_03819_),
    .B1(_03775_),
    .C1(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__a21oi_2 _18523_ (.A1(_03797_),
    .A2(_03819_),
    .B1(_03708_),
    .Y(_03822_));
 sky130_fd_sc_hd__or3b_2 _18524_ (.A(_03744_),
    .B(_03797_),
    .C_N(_10121_),
    .X(_03823_));
 sky130_fd_sc_hd__o211a_2 _18525_ (.A1(\decode.id_ex_rs2_data_reg[27] ),
    .A2(_03747_),
    .B1(_03822_),
    .C1(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__a21oi_2 _18526_ (.A1(_03709_),
    .A2(\decode.id_ex_imm_reg[27] ),
    .B1(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__nor2_2 _18527_ (.A(_03821_),
    .B(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2_2 _18528_ (.A(_03821_),
    .B(_03825_),
    .Y(_03827_));
 sky130_fd_sc_hd__or2b_2 _18529_ (.A(_03826_),
    .B_N(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__buf_1 _18530_ (.A(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__nor2_2 _18531_ (.A(_03814_),
    .B(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__o22a_2 _18532_ (.A1(\execute.csr_read_data_out_reg[25] ),
    .A2(_03659_),
    .B1(io_memory_address[25]),
    .B2(_03666_),
    .X(_03831_));
 sky130_fd_sc_hd__o31a_2 _18533_ (.A1(\execute.io_mem_memtoreg[1] ),
    .A2(\execute.io_mem_memtoreg[0] ),
    .A3(\execute.io_reg_pc[25] ),
    .B1(_03831_),
    .X(_03832_));
 sky130_fd_sc_hd__o21a_2 _18534_ (.A1(\memory.csr_read_data_out_reg[25] ),
    .A2(_09987_),
    .B1(_10110_),
    .X(_03833_));
 sky130_fd_sc_hd__o221a_2 _18535_ (.A1(_03656_),
    .A2(_03832_),
    .B1(_03701_),
    .B2(_03833_),
    .C1(_03670_),
    .X(_03834_));
 sky130_fd_sc_hd__o31a_2 _18536_ (.A1(\decode.id_ex_rs1_data_reg[25] ),
    .A2(_03817_),
    .A3(_03698_),
    .B1(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__o22a_2 _18537_ (.A1(\decode.id_ex_rs2_data_reg[25] ),
    .A2(_03747_),
    .B1(_03833_),
    .B2(_03764_),
    .X(_03836_));
 sky130_fd_sc_hd__o211a_2 _18538_ (.A1(_03759_),
    .A2(_03832_),
    .B1(_03727_),
    .C1(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__a21oi_2 _18539_ (.A1(_03709_),
    .A2(\decode.id_ex_imm_reg[25] ),
    .B1(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__or2_2 _18540_ (.A(_03835_),
    .B(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__or3_2 _18541_ (.A(\execute.csr_read_data_out_reg[24] ),
    .B(_03661_),
    .C(_03660_),
    .X(_03840_));
 sky130_fd_sc_hd__o221a_2 _18542_ (.A1(\execute.io_reg_pc[24] ),
    .A2(_03777_),
    .B1(_03666_),
    .B2(io_memory_address[24]),
    .C1(_03840_),
    .X(_03841_));
 sky130_fd_sc_hd__o22a_2 _18543_ (.A1(\memory.csr_read_data_out_reg[24] ),
    .A2(_09987_),
    .B1(_10104_),
    .B2(_10105_),
    .X(_03842_));
 sky130_fd_sc_hd__o22a_2 _18544_ (.A1(\decode.id_ex_rs1_data_reg[24] ),
    .A2(_03688_),
    .B1(_03842_),
    .B2(_03701_),
    .X(_03843_));
 sky130_fd_sc_hd__o211a_2 _18545_ (.A1(_03656_),
    .A2(_03841_),
    .B1(_03670_),
    .C1(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__o31a_2 _18546_ (.A1(_03715_),
    .A2(_03725_),
    .A3(_03841_),
    .B1(_03727_),
    .X(_03845_));
 sky130_fd_sc_hd__o221a_2 _18547_ (.A1(\decode.id_ex_rs2_data_reg[24] ),
    .A2(_03747_),
    .B1(_03764_),
    .B2(_03842_),
    .C1(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__a21oi_2 _18548_ (.A1(_03709_),
    .A2(\decode.id_ex_imm_reg[24] ),
    .B1(_03846_),
    .Y(_03847_));
 sky130_fd_sc_hd__or2_2 _18549_ (.A(_03844_),
    .B(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__nand2_2 _18550_ (.A(_03844_),
    .B(_03847_),
    .Y(_03849_));
 sky130_fd_sc_hd__and2_2 _18551_ (.A(_03848_),
    .B(_03849_),
    .X(_03850_));
 sky130_fd_sc_hd__buf_1 _18552_ (.A(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__nand2_2 _18553_ (.A(_03835_),
    .B(_03838_),
    .Y(_03852_));
 sky130_fd_sc_hd__and3_2 _18554_ (.A(_03839_),
    .B(_03851_),
    .C(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__xor2_2 _18555_ (.A(_03703_),
    .B(_03766_),
    .X(_03854_));
 sky130_fd_sc_hd__o22a_2 _18556_ (.A1(\execute.csr_read_data_out_reg[30] ),
    .A2(_03659_),
    .B1(io_memory_address[30]),
    .B2(_03666_),
    .X(_03855_));
 sky130_fd_sc_hd__o31a_2 _18557_ (.A1(\execute.io_mem_memtoreg[1] ),
    .A2(\execute.io_mem_memtoreg[0] ),
    .A3(\execute.io_reg_pc[30] ),
    .B1(_03855_),
    .X(_03856_));
 sky130_fd_sc_hd__o21a_2 _18558_ (.A1(\memory.csr_read_data_out_reg[30] ),
    .A2(_09988_),
    .B1(_10140_),
    .X(_03857_));
 sky130_fd_sc_hd__o221a_2 _18559_ (.A1(_03656_),
    .A2(_03856_),
    .B1(_03701_),
    .B2(_03857_),
    .C1(_03670_),
    .X(_03858_));
 sky130_fd_sc_hd__o31a_2 _18560_ (.A1(_03715_),
    .A2(_03725_),
    .A3(_03856_),
    .B1(_03728_),
    .X(_03859_));
 sky130_fd_sc_hd__o22a_2 _18561_ (.A1(\decode.id_ex_rs2_data_reg[30] ),
    .A2(_03747_),
    .B1(_03764_),
    .B2(_03857_),
    .X(_03860_));
 sky130_fd_sc_hd__a22oi_2 _18562_ (.A1(_03709_),
    .A2(\decode.id_ex_imm_reg[30] ),
    .B1(_03859_),
    .B2(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__o211a_2 _18563_ (.A1(\decode.id_ex_rs1_data_reg[30] ),
    .A2(_03689_),
    .B1(_03858_),
    .C1(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__o31a_2 _18564_ (.A1(\decode.id_ex_rs1_data_reg[30] ),
    .A2(_03817_),
    .A3(_03698_),
    .B1(_03858_),
    .X(_03863_));
 sky130_fd_sc_hd__nor2_2 _18565_ (.A(_03863_),
    .B(_03861_),
    .Y(_03864_));
 sky130_fd_sc_hd__nor2_2 _18566_ (.A(_03862_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__and3_2 _18567_ (.A(_03853_),
    .B(_03854_),
    .C(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__or4bb_2 _18568_ (.A(_03791_),
    .B(_03803_),
    .C_N(_03830_),
    .D_N(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__o22a_2 _18569_ (.A1(\memory.csr_read_data_out_reg[23] ),
    .A2(_09987_),
    .B1(_10099_),
    .B2(_10100_),
    .X(_03868_));
 sky130_fd_sc_hd__or3_2 _18570_ (.A(\execute.csr_read_data_out_reg[23] ),
    .B(_03661_),
    .C(_03660_),
    .X(_03869_));
 sky130_fd_sc_hd__o221a_2 _18571_ (.A1(\execute.io_reg_pc[23] ),
    .A2(_03777_),
    .B1(_03665_),
    .B2(io_memory_address[23]),
    .C1(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__o41a_2 _18572_ (.A1(_03768_),
    .A2(_03769_),
    .A3(_03770_),
    .A4(_03870_),
    .B1(_03670_),
    .X(_03871_));
 sky130_fd_sc_hd__o221a_2 _18573_ (.A1(_03868_),
    .A2(_03700_),
    .B1(_03688_),
    .B2(\decode.id_ex_rs1_data_reg[23] ),
    .C1(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__o221ai_2 _18574_ (.A1(_03759_),
    .A2(_03870_),
    .B1(\decode.id_ex_rs2_data_reg[23] ),
    .B2(_03747_),
    .C1(_03727_),
    .Y(_03873_));
 sky130_fd_sc_hd__o2111ai_2 _18575_ (.A1(\csr.io_csr_address[3] ),
    .A2(_09935_),
    .B1(_03733_),
    .C1(_03730_),
    .D1(_03736_),
    .Y(_03874_));
 sky130_fd_sc_hd__nor2_2 _18576_ (.A(_09929_),
    .B(\csr.io_csr_address[2] ),
    .Y(_03875_));
 sky130_fd_sc_hd__and2_2 _18577_ (.A(\decode.io_wb_rd[2] ),
    .B(\csr.io_csr_address[2] ),
    .X(_03876_));
 sky130_fd_sc_hd__o221a_2 _18578_ (.A1(_03710_),
    .A2(_09931_),
    .B1(_03875_),
    .B2(_03876_),
    .C1(_03735_),
    .X(_03877_));
 sky130_fd_sc_hd__o221a_2 _18579_ (.A1(\decode.io_wb_rd[0] ),
    .A2(_03721_),
    .B1(_03755_),
    .B2(_10194_),
    .C1(_03732_),
    .X(_03878_));
 sky130_fd_sc_hd__and4b_2 _18580_ (.A_N(_03874_),
    .B(_03673_),
    .C(_03877_),
    .D(_03878_),
    .X(_03879_));
 sky130_fd_sc_hd__and3_2 _18581_ (.A(_03879_),
    .B(_03759_),
    .C(_10101_),
    .X(_03880_));
 sky130_fd_sc_hd__o2bb2a_2 _18582_ (.A1_N(_03708_),
    .A2_N(\decode.id_ex_imm_reg[23] ),
    .B1(_03873_),
    .B2(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__and2_2 _18583_ (.A(_03872_),
    .B(_03881_),
    .X(_03882_));
 sky130_fd_sc_hd__o21a_2 _18584_ (.A1(\memory.csr_read_data_out_reg[22] ),
    .A2(_09987_),
    .B1(_10095_),
    .X(_03883_));
 sky130_fd_sc_hd__o22a_2 _18585_ (.A1(_03659_),
    .A2(\execute.csr_read_data_out_reg[22] ),
    .B1(\execute.io_reg_pc[22] ),
    .B2(_03777_),
    .X(_03884_));
 sky130_fd_sc_hd__o21ai_2 _18586_ (.A1(io_memory_address[22]),
    .A2(_03666_),
    .B1(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__a21oi_2 _18587_ (.A1(_03817_),
    .A2(_03885_),
    .B1(_03774_),
    .Y(_03886_));
 sky130_fd_sc_hd__o221a_2 _18588_ (.A1(_03688_),
    .A2(\decode.id_ex_rs1_data_reg[22] ),
    .B1(_03700_),
    .B2(_03883_),
    .C1(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__buf_1 _18589_ (.A(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__buf_1 _18590_ (.A(_03706_),
    .X(_03889_));
 sky130_fd_sc_hd__buf_1 _18591_ (.A(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__a21oi_2 _18592_ (.A1(_03797_),
    .A2(_03885_),
    .B1(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__o22a_2 _18593_ (.A1(\decode.id_ex_rs2_data_reg[22] ),
    .A2(_03746_),
    .B1(_03764_),
    .B2(_03883_),
    .X(_03892_));
 sky130_fd_sc_hd__a22oi_2 _18594_ (.A1(_03708_),
    .A2(\decode.id_ex_imm_reg[22] ),
    .B1(_03891_),
    .B2(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__and2_2 _18595_ (.A(_03887_),
    .B(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__or3_2 _18596_ (.A(\execute.io_mem_memtoreg[1] ),
    .B(\execute.io_mem_memtoreg[0] ),
    .C(\execute.io_reg_pc[19] ),
    .X(_03895_));
 sky130_fd_sc_hd__o221a_2 _18597_ (.A1(\execute.csr_read_data_out_reg[19] ),
    .A2(_03659_),
    .B1(io_memory_address[19]),
    .B2(_03665_),
    .C1(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__o221ai_2 _18598_ (.A1(_03759_),
    .A2(_03896_),
    .B1(\decode.id_ex_rs2_data_reg[19] ),
    .B2(_03746_),
    .C1(_03727_),
    .Y(_03897_));
 sky130_fd_sc_hd__a21oi_2 _18599_ (.A1(_10080_),
    .A2(_03785_),
    .B1(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__and2_2 _18600_ (.A(_03707_),
    .B(\decode.id_ex_imm_reg[19] ),
    .X(_03899_));
 sky130_fd_sc_hd__o22a_2 _18601_ (.A1(\memory.csr_read_data_out_reg[19] ),
    .A2(_09986_),
    .B1(_10078_),
    .B2(_10079_),
    .X(_03900_));
 sky130_fd_sc_hd__o41a_2 _18602_ (.A1(_03768_),
    .A2(_03769_),
    .A3(_03770_),
    .A4(_03896_),
    .B1(_03669_),
    .X(_03901_));
 sky130_fd_sc_hd__o221ai_2 _18603_ (.A1(_03900_),
    .A2(_03700_),
    .B1(_03688_),
    .B2(\decode.id_ex_rs1_data_reg[19] ),
    .C1(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__or3_2 _18604_ (.A(_03898_),
    .B(_03899_),
    .C(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__o22a_2 _18605_ (.A1(_03658_),
    .A2(\execute.csr_read_data_out_reg[17] ),
    .B1(\execute.io_reg_pc[17] ),
    .B2(_03776_),
    .X(_03904_));
 sky130_fd_sc_hd__o21ai_2 _18606_ (.A1(io_memory_address[17]),
    .A2(_03665_),
    .B1(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__a221oi_2 _18607_ (.A1(_03797_),
    .A2(_03905_),
    .B1(_03785_),
    .B2(_10068_),
    .C1(_03889_),
    .Y(_03906_));
 sky130_fd_sc_hd__a311o_2 _18608_ (.A1(_03751_),
    .A2(_03752_),
    .A3(_03757_),
    .B1(_03784_),
    .C1(\decode.id_ex_rs2_data_reg[17] ),
    .X(_03907_));
 sky130_fd_sc_hd__buf_1 _18609_ (.A(_03686_),
    .X(_03908_));
 sky130_fd_sc_hd__o2bb2a_2 _18610_ (.A1_N(_10067_),
    .A2_N(_10066_),
    .B1(\memory.csr_read_data_out_reg[17] ),
    .B2(_09986_),
    .X(_03909_));
 sky130_fd_sc_hd__a21oi_2 _18611_ (.A1(_03817_),
    .A2(_03905_),
    .B1(_03774_),
    .Y(_03910_));
 sky130_fd_sc_hd__o221ai_2 _18612_ (.A1(\decode.id_ex_rs1_data_reg[17] ),
    .A2(_03908_),
    .B1(_03909_),
    .B2(_03700_),
    .C1(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__a221o_2 _18613_ (.A1(_03708_),
    .A2(\decode.id_ex_imm_reg[17] ),
    .B1(_03906_),
    .B2(_03907_),
    .C1(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__o2bb2a_2 _18614_ (.A1_N(_10072_),
    .A2_N(_10071_),
    .B1(_09986_),
    .B2(\memory.csr_read_data_out_reg[18] ),
    .X(_03913_));
 sky130_fd_sc_hd__buf_1 _18615_ (.A(_03699_),
    .X(_03914_));
 sky130_fd_sc_hd__o22a_2 _18616_ (.A1(_03659_),
    .A2(\execute.csr_read_data_out_reg[18] ),
    .B1(\execute.io_reg_pc[18] ),
    .B2(_03777_),
    .X(_03915_));
 sky130_fd_sc_hd__o21ai_2 _18617_ (.A1(io_memory_address[18]),
    .A2(_03665_),
    .B1(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__a21oi_2 _18618_ (.A1(_03817_),
    .A2(_03916_),
    .B1(_03774_),
    .Y(_03917_));
 sky130_fd_sc_hd__o221a_2 _18619_ (.A1(\decode.id_ex_rs1_data_reg[18] ),
    .A2(_03908_),
    .B1(_03913_),
    .B2(_03914_),
    .C1(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__a311o_2 _18620_ (.A1(_03751_),
    .A2(_03752_),
    .A3(_03757_),
    .B1(_03784_),
    .C1(\decode.id_ex_rs2_data_reg[18] ),
    .X(_03919_));
 sky130_fd_sc_hd__a21oi_2 _18621_ (.A1(_03797_),
    .A2(_03916_),
    .B1(_03889_),
    .Y(_03920_));
 sky130_fd_sc_hd__nand2_2 _18622_ (.A(_03785_),
    .B(_10073_),
    .Y(_03921_));
 sky130_fd_sc_hd__and2_2 _18623_ (.A(_03889_),
    .B(\decode.id_ex_imm_reg[18] ),
    .X(_03922_));
 sky130_fd_sc_hd__a31oi_2 _18624_ (.A1(_03919_),
    .A2(_03920_),
    .A3(_03921_),
    .B1(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__nand2_2 _18625_ (.A(_03918_),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__o22a_2 _18626_ (.A1(\memory.csr_read_data_out_reg[16] ),
    .A2(_09987_),
    .B1(_10061_),
    .B2(_10062_),
    .X(_03925_));
 sky130_fd_sc_hd__o22a_2 _18627_ (.A1(_03659_),
    .A2(\execute.csr_read_data_out_reg[16] ),
    .B1(\execute.io_reg_pc[16] ),
    .B2(_03777_),
    .X(_03926_));
 sky130_fd_sc_hd__o21ai_2 _18628_ (.A1(io_memory_address[16]),
    .A2(_03665_),
    .B1(_03926_),
    .Y(_03927_));
 sky130_fd_sc_hd__a21oi_2 _18629_ (.A1(_03817_),
    .A2(_03927_),
    .B1(_03774_),
    .Y(_03928_));
 sky130_fd_sc_hd__o221a_2 _18630_ (.A1(_03925_),
    .A2(_03700_),
    .B1(_03688_),
    .B2(\decode.id_ex_rs1_data_reg[16] ),
    .C1(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__nor2_2 _18631_ (.A(\decode.id_ex_rs2_data_reg[16] ),
    .B(_03746_),
    .Y(_03930_));
 sky130_fd_sc_hd__a211o_2 _18632_ (.A1(_03927_),
    .A2(_03797_),
    .B1(_03707_),
    .C1(_03930_),
    .X(_03931_));
 sky130_fd_sc_hd__a21oi_2 _18633_ (.A1(_10063_),
    .A2(_03785_),
    .B1(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__a21oi_2 _18634_ (.A1(_03708_),
    .A2(\decode.id_ex_imm_reg[16] ),
    .B1(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__o221a_2 _18635_ (.A1(_03909_),
    .A2(_03914_),
    .B1(_03908_),
    .B2(\decode.id_ex_rs1_data_reg[17] ),
    .C1(_03910_),
    .X(_03934_));
 sky130_fd_sc_hd__a22oi_2 _18636_ (.A1(_03890_),
    .A2(\decode.id_ex_imm_reg[17] ),
    .B1(_03906_),
    .B2(_03907_),
    .Y(_03935_));
 sky130_fd_sc_hd__o22ai_2 _18637_ (.A1(_03929_),
    .A2(_03933_),
    .B1(_03934_),
    .B2(_03935_),
    .Y(_03936_));
 sky130_fd_sc_hd__o21a_2 _18638_ (.A1(_03898_),
    .A2(_03899_),
    .B1(_03902_),
    .X(_03937_));
 sky130_fd_sc_hd__nor2_2 _18639_ (.A(_03918_),
    .B(_03923_),
    .Y(_03938_));
 sky130_fd_sc_hd__a311o_2 _18640_ (.A1(_03912_),
    .A2(_03924_),
    .A3(_03936_),
    .B1(_03937_),
    .C1(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__o2bb2a_2 _18641_ (.A1_N(_10090_),
    .A2_N(_10089_),
    .B1(\memory.csr_read_data_out_reg[21] ),
    .B2(_10010_),
    .X(_03940_));
 sky130_fd_sc_hd__o22a_2 _18642_ (.A1(_03658_),
    .A2(\execute.csr_read_data_out_reg[21] ),
    .B1(\execute.io_reg_pc[21] ),
    .B2(_03776_),
    .X(_03941_));
 sky130_fd_sc_hd__o21ai_2 _18643_ (.A1(io_memory_address[21]),
    .A2(_03665_),
    .B1(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__a21oi_2 _18644_ (.A1(_03816_),
    .A2(_03942_),
    .B1(_03773_),
    .Y(_03943_));
 sky130_fd_sc_hd__o221a_2 _18645_ (.A1(\decode.id_ex_rs1_data_reg[21] ),
    .A2(_03687_),
    .B1(_03940_),
    .B2(_03914_),
    .C1(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__a21oi_2 _18646_ (.A1(_03797_),
    .A2(_03942_),
    .B1(_03889_),
    .Y(_03945_));
 sky130_fd_sc_hd__o22a_2 _18647_ (.A1(\decode.id_ex_rs2_data_reg[21] ),
    .A2(_03745_),
    .B1(_03940_),
    .B2(_03763_),
    .X(_03946_));
 sky130_fd_sc_hd__a22o_2 _18648_ (.A1(_03707_),
    .A2(\decode.id_ex_imm_reg[21] ),
    .B1(_03945_),
    .B2(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__and2b_2 _18649_ (.A_N(_03944_),
    .B(_03947_),
    .X(_03948_));
 sky130_fd_sc_hd__nand2_2 _18650_ (.A(_10086_),
    .B(_03785_),
    .Y(_03949_));
 sky130_fd_sc_hd__or3_2 _18651_ (.A(\execute.csr_read_data_out_reg[20] ),
    .B(_03661_),
    .C(_03660_),
    .X(_03950_));
 sky130_fd_sc_hd__o221a_2 _18652_ (.A1(\execute.io_reg_pc[20] ),
    .A2(_03776_),
    .B1(_03664_),
    .B2(io_memory_address[20]),
    .C1(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__o31a_2 _18653_ (.A1(_03715_),
    .A2(_03725_),
    .A3(_03951_),
    .B1(_03727_),
    .X(_03952_));
 sky130_fd_sc_hd__o211ai_2 _18654_ (.A1(\decode.id_ex_rs2_data_reg[20] ),
    .A2(_03746_),
    .B1(_03949_),
    .C1(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__nand2_2 _18655_ (.A(_03707_),
    .B(\decode.id_ex_imm_reg[20] ),
    .Y(_03954_));
 sky130_fd_sc_hd__o22ai_2 _18656_ (.A1(_03655_),
    .A2(_03951_),
    .B1(\decode.id_ex_rs1_data_reg[20] ),
    .B2(_03687_),
    .Y(_03955_));
 sky130_fd_sc_hd__a211oi_2 _18657_ (.A1(_10086_),
    .A2(_03771_),
    .B1(_03774_),
    .C1(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__a21oi_2 _18658_ (.A1(_03953_),
    .A2(_03954_),
    .B1(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__a211oi_2 _18659_ (.A1(_03903_),
    .A2(_03939_),
    .B1(_03948_),
    .C1(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__nand2_2 _18660_ (.A(_03953_),
    .B(_03954_),
    .Y(_03959_));
 sky130_fd_sc_hd__a2111o_2 _18661_ (.A1(_10086_),
    .A2(_03772_),
    .B1(_03774_),
    .C1(_03955_),
    .D1(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__o21ai_2 _18662_ (.A1(\decode.id_ex_rs1_data_reg[21] ),
    .A2(_03688_),
    .B1(_03943_),
    .Y(_03961_));
 sky130_fd_sc_hd__a211o_2 _18663_ (.A1(_10091_),
    .A2(_03772_),
    .B1(_03961_),
    .C1(_03947_),
    .X(_03962_));
 sky130_fd_sc_hd__o21ai_2 _18664_ (.A1(_03948_),
    .A2(_03960_),
    .B1(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__or3_2 _18665_ (.A(_03894_),
    .B(_03958_),
    .C(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__o221a_2 _18666_ (.A1(_03888_),
    .A2(_03893_),
    .B1(_03872_),
    .B2(_03881_),
    .C1(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__o22a_2 _18667_ (.A1(\execute.csr_read_data_out_reg[3] ),
    .A2(_03657_),
    .B1(\execute.io_reg_pc[3] ),
    .B2(_03662_),
    .X(_03966_));
 sky130_fd_sc_hd__o21ai_2 _18668_ (.A1(io_memory_address[3]),
    .A2(_03664_),
    .B1(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__and4_2 _18669_ (.A(_09921_),
    .B(_03645_),
    .C(_03641_),
    .D(_03643_),
    .X(_03968_));
 sky130_fd_sc_hd__a41o_2 _18670_ (.A1(_03967_),
    .A2(_03654_),
    .A3(_03968_),
    .A4(_03649_),
    .B1(_03773_),
    .X(_03969_));
 sky130_fd_sc_hd__nor2_2 _18671_ (.A(\decode.id_ex_rs1_data_reg[3] ),
    .B(_03686_),
    .Y(_03970_));
 sky130_fd_sc_hd__a211oi_2 _18672_ (.A1(_09974_),
    .A2(_03771_),
    .B1(_03969_),
    .C1(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__a41o_2 _18673_ (.A1(_03967_),
    .A2(_03757_),
    .A3(_03752_),
    .A4(_03751_),
    .B1(\decode.id_ex_immsrc_reg ),
    .X(_03972_));
 sky130_fd_sc_hd__o211ai_2 _18674_ (.A1(_03714_),
    .A2(_03724_),
    .B1(_09974_),
    .C1(_03879_),
    .Y(_03973_));
 sky130_fd_sc_hd__o21ai_2 _18675_ (.A1(\decode.id_ex_rs2_data_reg[3] ),
    .A2(_03745_),
    .B1(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__o2bb2a_2 _18676_ (.A1_N(_03706_),
    .A2_N(\decode.id_ex_imm_reg[3] ),
    .B1(_03972_),
    .B2(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__nor2_2 _18677_ (.A(_03971_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__o211ai_2 _18678_ (.A1(_03675_),
    .A2(_03685_),
    .B1(\decode.id_ex_rs1_data_reg[0] ),
    .C1(_03655_),
    .Y(_03977_));
 sky130_fd_sc_hd__o2bb2a_2 _18679_ (.A1_N(_09945_),
    .A2_N(_09948_),
    .B1(\memory.csr_read_data_out_reg[0] ),
    .B2(_09942_),
    .X(_03978_));
 sky130_fd_sc_hd__nand3_2 _18680_ (.A(_03655_),
    .B(_03698_),
    .C(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__or2_2 _18681_ (.A(\execute.csr_read_data_out_reg[0] ),
    .B(_03657_),
    .X(_03980_));
 sky130_fd_sc_hd__o221a_2 _18682_ (.A1(_03662_),
    .A2(\execute.io_reg_pc[0] ),
    .B1(io_memory_address[0]),
    .B2(_03663_),
    .C1(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__nand2_2 _18683_ (.A(_03815_),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__a31o_2 _18684_ (.A1(_03977_),
    .A2(_03979_),
    .A3(_03982_),
    .B1(_03773_),
    .X(_03983_));
 sky130_fd_sc_hd__a21oi_2 _18685_ (.A1(_03796_),
    .A2(_03981_),
    .B1(\decode.id_ex_immsrc_reg ),
    .Y(_03984_));
 sky130_fd_sc_hd__o211ai_2 _18686_ (.A1(_03714_),
    .A2(_03724_),
    .B1(\decode.id_ex_rs2_data_reg[0] ),
    .C1(_03744_),
    .Y(_03985_));
 sky130_fd_sc_hd__o211ai_2 _18687_ (.A1(_03715_),
    .A2(_03725_),
    .B1(_03784_),
    .C1(_03978_),
    .Y(_03986_));
 sky130_fd_sc_hd__nor2_2 _18688_ (.A(\decode.id_ex_imm_reg[0] ),
    .B(_03726_),
    .Y(_03987_));
 sky130_fd_sc_hd__a31oi_2 _18689_ (.A1(_03984_),
    .A2(_03985_),
    .A3(_03986_),
    .B1(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__buf_1 _18690_ (.A(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__o211ai_2 _18691_ (.A1(_03714_),
    .A2(_03724_),
    .B1(_03744_),
    .C1(_03598_),
    .Y(_03990_));
 sky130_fd_sc_hd__o211ai_2 _18692_ (.A1(_03714_),
    .A2(_03724_),
    .B1(_09963_),
    .C1(_03784_),
    .Y(_03991_));
 sky130_fd_sc_hd__nand3b_2 _18693_ (.A_N(\execute.csr_read_data_out_reg[1] ),
    .B(\execute.io_mem_memtoreg[0] ),
    .C(\execute.io_mem_memtoreg[1] ),
    .Y(_03992_));
 sky130_fd_sc_hd__o21ba_2 _18694_ (.A1(\execute.io_mem_memtoreg[1] ),
    .A2(\execute.io_mem_memtoreg[0] ),
    .B1_N(io_memory_address[1]),
    .X(_03993_));
 sky130_fd_sc_hd__nand2_2 _18695_ (.A(_03993_),
    .B(_03657_),
    .Y(_03994_));
 sky130_fd_sc_hd__o211ai_2 _18696_ (.A1(_03662_),
    .A2(\execute.io_reg_pc[1] ),
    .B1(_03992_),
    .C1(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__a41oi_2 _18697_ (.A1(_03752_),
    .A2(_03995_),
    .A3(_03757_),
    .A4(_03751_),
    .B1(\decode.id_ex_immsrc_reg ),
    .Y(_03996_));
 sky130_fd_sc_hd__nand3_2 _18698_ (.A(_03990_),
    .B(_03991_),
    .C(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__nand2_2 _18699_ (.A(\decode.id_ex_immsrc_reg ),
    .B(\decode.id_ex_imm_reg[1] ),
    .Y(_03998_));
 sky130_fd_sc_hd__o311a_2 _18700_ (.A1(_03768_),
    .A2(_03769_),
    .A3(_03770_),
    .B1(_09963_),
    .C1(_03698_),
    .X(_03999_));
 sky130_fd_sc_hd__o21bai_2 _18701_ (.A1(_03675_),
    .A2(_03685_),
    .B1_N(\decode.id_ex_rs1_data_reg[1] ),
    .Y(_04000_));
 sky130_fd_sc_hd__a41oi_2 _18702_ (.A1(_03968_),
    .A2(_03995_),
    .A3(_03654_),
    .A4(_03649_),
    .B1(\decode.id_ex_islui_reg ),
    .Y(_04001_));
 sky130_fd_sc_hd__o21ai_2 _18703_ (.A1(_03815_),
    .A2(_04000_),
    .B1(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__o2bb2a_2 _18704_ (.A1_N(_03997_),
    .A2_N(_03998_),
    .B1(_03999_),
    .B2(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__o211a_2 _18705_ (.A1(_03816_),
    .A2(_04000_),
    .B1(_04001_),
    .C1(_03998_),
    .X(_04004_));
 sky130_fd_sc_hd__nand3_2 _18706_ (.A(_09963_),
    .B(_03655_),
    .C(_03698_),
    .Y(_04005_));
 sky130_fd_sc_hd__nand3_2 _18707_ (.A(_04004_),
    .B(_04005_),
    .C(_03997_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand2_2 _18708_ (.A(_03889_),
    .B(\decode.id_ex_imm_reg[3] ),
    .Y(_04007_));
 sky130_fd_sc_hd__o211a_2 _18709_ (.A1(_03972_),
    .A2(_03974_),
    .B1(_04007_),
    .C1(_03971_),
    .X(_04008_));
 sky130_fd_sc_hd__or2_2 _18710_ (.A(_04008_),
    .B(_03976_),
    .X(_04009_));
 sky130_fd_sc_hd__o2bb2a_2 _18711_ (.A1_N(_09967_),
    .A2_N(_09968_),
    .B1(\memory.csr_read_data_out_reg[2] ),
    .B2(_09942_),
    .X(_04010_));
 sky130_fd_sc_hd__o22a_2 _18712_ (.A1(_03657_),
    .A2(\execute.csr_read_data_out_reg[2] ),
    .B1(\execute.io_reg_pc[2] ),
    .B2(_03662_),
    .X(_04011_));
 sky130_fd_sc_hd__o21ai_2 _18713_ (.A1(io_memory_address[2]),
    .A2(_03663_),
    .B1(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__a21oi_2 _18714_ (.A1(_03815_),
    .A2(_04012_),
    .B1(_03773_),
    .Y(_04013_));
 sky130_fd_sc_hd__o221a_2 _18715_ (.A1(_04010_),
    .A2(_03699_),
    .B1(_03686_),
    .B2(\decode.id_ex_rs1_data_reg[2] ),
    .C1(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__a21oi_2 _18716_ (.A1(_03796_),
    .A2(_04012_),
    .B1(\decode.id_ex_immsrc_reg ),
    .Y(_04015_));
 sky130_fd_sc_hd__nand3b_2 _18717_ (.A_N(\decode.id_ex_rs2_data_reg[2] ),
    .B(_03758_),
    .C(_03744_),
    .Y(_04016_));
 sky130_fd_sc_hd__o211ai_2 _18718_ (.A1(_03714_),
    .A2(_03724_),
    .B1(_03784_),
    .C1(_09969_),
    .Y(_04017_));
 sky130_fd_sc_hd__inv_2 _18719_ (.A(\decode.id_ex_imm_reg[2] ),
    .Y(_04018_));
 sky130_fd_sc_hd__nor2_2 _18720_ (.A(_03726_),
    .B(_04018_),
    .Y(_04019_));
 sky130_fd_sc_hd__a31oi_2 _18721_ (.A1(_04015_),
    .A2(_04016_),
    .A3(_04017_),
    .B1(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__buf_1 _18722_ (.A(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__nor2_2 _18723_ (.A(_04014_),
    .B(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__and2_2 _18724_ (.A(_04014_),
    .B(_04020_),
    .X(_04023_));
 sky130_fd_sc_hd__or2_2 _18725_ (.A(_04022_),
    .B(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__nor2_2 _18726_ (.A(_04009_),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__o311a_2 _18727_ (.A1(_03983_),
    .A2(_03989_),
    .A3(_04003_),
    .B1(_04006_),
    .C1(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__a211o_2 _18728_ (.A1(_09974_),
    .A2(_03771_),
    .B1(_03969_),
    .C1(_03970_),
    .X(_04027_));
 sky130_fd_sc_hd__o21ai_2 _18729_ (.A1(_03972_),
    .A2(_03974_),
    .B1(_04007_),
    .Y(_04028_));
 sky130_fd_sc_hd__o21a_2 _18730_ (.A1(_04027_),
    .A2(_04028_),
    .B1(_04022_),
    .X(_04029_));
 sky130_fd_sc_hd__o2bb2a_2 _18731_ (.A1_N(_09982_),
    .A2_N(_09979_),
    .B1(_10010_),
    .B2(\memory.csr_read_data_out_reg[4] ),
    .X(_04030_));
 sky130_fd_sc_hd__o22a_2 _18732_ (.A1(\execute.csr_read_data_out_reg[4] ),
    .A2(_03658_),
    .B1(\execute.io_reg_pc[4] ),
    .B2(_03662_),
    .X(_04031_));
 sky130_fd_sc_hd__o21ai_2 _18733_ (.A1(io_memory_address[4]),
    .A2(_03664_),
    .B1(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__a21oi_2 _18734_ (.A1(_03816_),
    .A2(_04032_),
    .B1(_03773_),
    .Y(_04033_));
 sky130_fd_sc_hd__o221a_2 _18735_ (.A1(\decode.id_ex_rs1_data_reg[4] ),
    .A2(_03687_),
    .B1(_04030_),
    .B2(_03699_),
    .C1(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__a21oi_2 _18736_ (.A1(_03796_),
    .A2(_04032_),
    .B1(_03706_),
    .Y(_04035_));
 sky130_fd_sc_hd__o21ai_2 _18737_ (.A1(\decode.id_ex_rs2_data_reg[4] ),
    .A2(_03745_),
    .B1(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__and3_2 _18738_ (.A(_09983_),
    .B(_03759_),
    .C(_03784_),
    .X(_04037_));
 sky130_fd_sc_hd__o2bb2ai_2 _18739_ (.A1_N(_03889_),
    .A2_N(\decode.id_ex_imm_reg[4] ),
    .B1(_04036_),
    .B2(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__xnor2_2 _18740_ (.A(_04034_),
    .B(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__or3_2 _18741_ (.A(\execute.csr_read_data_out_reg[5] ),
    .B(_03661_),
    .C(_03660_),
    .X(_04040_));
 sky130_fd_sc_hd__o221a_2 _18742_ (.A1(\execute.io_reg_pc[5] ),
    .A2(_03776_),
    .B1(_03664_),
    .B2(io_memory_address[5]),
    .C1(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__o21a_2 _18743_ (.A1(\memory.csr_read_data_out_reg[5] ),
    .A2(_10010_),
    .B1(_09991_),
    .X(_04042_));
 sky130_fd_sc_hd__o22a_2 _18744_ (.A1(\decode.id_ex_rs1_data_reg[5] ),
    .A2(_03686_),
    .B1(_04042_),
    .B2(_03699_),
    .X(_04043_));
 sky130_fd_sc_hd__o211a_2 _18745_ (.A1(_03656_),
    .A2(_04041_),
    .B1(_03669_),
    .C1(_04043_),
    .X(_04044_));
 sky130_fd_sc_hd__buf_1 _18746_ (.A(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__o21ai_2 _18747_ (.A1(_03714_),
    .A2(_03724_),
    .B1(_03784_),
    .Y(_04046_));
 sky130_fd_sc_hd__o31a_2 _18748_ (.A1(_03715_),
    .A2(_03725_),
    .A3(_04041_),
    .B1(_03726_),
    .X(_04047_));
 sky130_fd_sc_hd__o221a_2 _18749_ (.A1(_04042_),
    .A2(_04046_),
    .B1(_03746_),
    .B2(\decode.id_ex_rs2_data_reg[5] ),
    .C1(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__a21oi_2 _18750_ (.A1(_03890_),
    .A2(\decode.id_ex_imm_reg[5] ),
    .B1(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__nor2_2 _18751_ (.A(_04045_),
    .B(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__and2_2 _18752_ (.A(_04044_),
    .B(_04049_),
    .X(_04051_));
 sky130_fd_sc_hd__nor2_2 _18753_ (.A(_04050_),
    .B(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__o311ai_2 _18754_ (.A1(_03976_),
    .A2(_04026_),
    .A3(_04029_),
    .B1(_04039_),
    .C1(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__buf_1 _18755_ (.A(_04034_),
    .X(_04054_));
 sky130_fd_sc_hd__o2bb2a_2 _18756_ (.A1_N(_03706_),
    .A2_N(\decode.id_ex_imm_reg[4] ),
    .B1(_04036_),
    .B2(_04037_),
    .X(_04055_));
 sky130_fd_sc_hd__buf_1 _18757_ (.A(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__or3_2 _18758_ (.A(_04051_),
    .B(_04054_),
    .C(_04056_),
    .X(_04057_));
 sky130_fd_sc_hd__or3_2 _18759_ (.A(\execute.csr_read_data_out_reg[7] ),
    .B(_03661_),
    .C(_03660_),
    .X(_04058_));
 sky130_fd_sc_hd__o221a_2 _18760_ (.A1(\execute.io_reg_pc[7] ),
    .A2(_03777_),
    .B1(_03665_),
    .B2(io_memory_address[7]),
    .C1(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__o22a_2 _18761_ (.A1(\memory.csr_read_data_out_reg[7] ),
    .A2(_09986_),
    .B1(_10002_),
    .B2(_10006_),
    .X(_04060_));
 sky130_fd_sc_hd__o22a_2 _18762_ (.A1(\decode.id_ex_rs1_data_reg[7] ),
    .A2(_03908_),
    .B1(_04060_),
    .B2(_03914_),
    .X(_04061_));
 sky130_fd_sc_hd__o211a_2 _18763_ (.A1(_03656_),
    .A2(_04059_),
    .B1(_03670_),
    .C1(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__o31a_2 _18764_ (.A1(_03715_),
    .A2(_03725_),
    .A3(_04059_),
    .B1(_03727_),
    .X(_04063_));
 sky130_fd_sc_hd__o221a_2 _18765_ (.A1(\decode.id_ex_rs2_data_reg[7] ),
    .A2(_03746_),
    .B1(_03764_),
    .B2(_04060_),
    .C1(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__a21oi_2 _18766_ (.A1(_03708_),
    .A2(\decode.id_ex_imm_reg[7] ),
    .B1(_04064_),
    .Y(_04065_));
 sky130_fd_sc_hd__or3_2 _18767_ (.A(\execute.csr_read_data_out_reg[6] ),
    .B(_03661_),
    .C(_03660_),
    .X(_04066_));
 sky130_fd_sc_hd__o221a_2 _18768_ (.A1(\execute.io_reg_pc[6] ),
    .A2(_03776_),
    .B1(_03664_),
    .B2(io_memory_address[6]),
    .C1(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__o21a_2 _18769_ (.A1(\memory.csr_read_data_out_reg[6] ),
    .A2(_10010_),
    .B1(_09997_),
    .X(_04068_));
 sky130_fd_sc_hd__o22a_2 _18770_ (.A1(\decode.id_ex_rs1_data_reg[6] ),
    .A2(_03687_),
    .B1(_04068_),
    .B2(_03699_),
    .X(_04069_));
 sky130_fd_sc_hd__o211a_2 _18771_ (.A1(_03656_),
    .A2(_04067_),
    .B1(_03670_),
    .C1(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__o31a_2 _18772_ (.A1(_03715_),
    .A2(_03725_),
    .A3(_04067_),
    .B1(_03726_),
    .X(_04071_));
 sky130_fd_sc_hd__o221a_2 _18773_ (.A1(\decode.id_ex_rs2_data_reg[6] ),
    .A2(_03746_),
    .B1(_03764_),
    .B2(_04068_),
    .C1(_04071_),
    .X(_04072_));
 sky130_fd_sc_hd__a21oi_2 _18774_ (.A1(_03890_),
    .A2(\decode.id_ex_imm_reg[6] ),
    .B1(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__or2_2 _18775_ (.A(_04070_),
    .B(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__buf_1 _18776_ (.A(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__o221a_2 _18777_ (.A1(_04045_),
    .A2(_04049_),
    .B1(_04062_),
    .B2(_04065_),
    .C1(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__o21ba_2 _18778_ (.A1(\memory.csr_read_data_out_reg[14] ),
    .A2(_09986_),
    .B1_N(_10051_),
    .X(_04077_));
 sky130_fd_sc_hd__o22a_2 _18779_ (.A1(_03658_),
    .A2(\execute.csr_read_data_out_reg[14] ),
    .B1(\execute.io_reg_pc[14] ),
    .B2(_03776_),
    .X(_04078_));
 sky130_fd_sc_hd__o21ai_2 _18780_ (.A1(io_memory_address[14]),
    .A2(_03665_),
    .B1(_04078_),
    .Y(_04079_));
 sky130_fd_sc_hd__a21oi_2 _18781_ (.A1(_03817_),
    .A2(_04079_),
    .B1(_03774_),
    .Y(_04080_));
 sky130_fd_sc_hd__o221ai_2 _18782_ (.A1(\decode.id_ex_rs1_data_reg[14] ),
    .A2(_03908_),
    .B1(_04077_),
    .B2(_03700_),
    .C1(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__a21oi_2 _18783_ (.A1(_03796_),
    .A2(_04079_),
    .B1(_03889_),
    .Y(_04082_));
 sky130_fd_sc_hd__o221ai_2 _18784_ (.A1(\decode.id_ex_rs2_data_reg[14] ),
    .A2(_03746_),
    .B1(_04077_),
    .B2(_03764_),
    .C1(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__nand2_2 _18785_ (.A(_03707_),
    .B(\decode.id_ex_imm_reg[14] ),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_2 _18786_ (.A(_04083_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__xnor2_2 _18787_ (.A(_04081_),
    .B(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__o2bb2a_2 _18788_ (.A1_N(_10056_),
    .A2_N(_10055_),
    .B1(_10010_),
    .B2(\memory.csr_read_data_out_reg[15] ),
    .X(_04087_));
 sky130_fd_sc_hd__o22a_2 _18789_ (.A1(_03658_),
    .A2(\execute.csr_read_data_out_reg[15] ),
    .B1(\execute.io_reg_pc[15] ),
    .B2(_03776_),
    .X(_04088_));
 sky130_fd_sc_hd__o21ai_2 _18790_ (.A1(io_memory_address[15]),
    .A2(_03664_),
    .B1(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__a21oi_2 _18791_ (.A1(_03816_),
    .A2(_04089_),
    .B1(_03774_),
    .Y(_04090_));
 sky130_fd_sc_hd__o221ai_2 _18792_ (.A1(\decode.id_ex_rs1_data_reg[15] ),
    .A2(_03908_),
    .B1(_04087_),
    .B2(_03914_),
    .C1(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__a21oi_2 _18793_ (.A1(_03796_),
    .A2(_04089_),
    .B1(_03706_),
    .Y(_04092_));
 sky130_fd_sc_hd__o221a_2 _18794_ (.A1(\decode.id_ex_rs2_data_reg[15] ),
    .A2(_03745_),
    .B1(_04087_),
    .B2(_04046_),
    .C1(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__a21oi_2 _18795_ (.A1(_03707_),
    .A2(\decode.id_ex_imm_reg[15] ),
    .B1(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__xor2_2 _18796_ (.A(_04091_),
    .B(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__a31oi_2 _18797_ (.A1(_10045_),
    .A2(_10044_),
    .A3(_09942_),
    .B1(_10046_),
    .Y(_04096_));
 sky130_fd_sc_hd__o22a_2 _18798_ (.A1(\execute.io_reg_pc[13] ),
    .A2(_03776_),
    .B1(io_memory_address[13]),
    .B2(_03664_),
    .X(_04097_));
 sky130_fd_sc_hd__o21ai_2 _18799_ (.A1(\execute.csr_read_data_out_reg[13] ),
    .A2(_03658_),
    .B1(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__a21oi_2 _18800_ (.A1(_04098_),
    .A2(_03816_),
    .B1(_03773_),
    .Y(_04099_));
 sky130_fd_sc_hd__o221ai_2 _18801_ (.A1(_04096_),
    .A2(_03699_),
    .B1(_03687_),
    .B2(\decode.id_ex_rs1_data_reg[13] ),
    .C1(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__a21oi_2 _18802_ (.A1(_04098_),
    .A2(_03796_),
    .B1(_03706_),
    .Y(_04101_));
 sky130_fd_sc_hd__o22a_2 _18803_ (.A1(\decode.id_ex_rs2_data_reg[13] ),
    .A2(_03745_),
    .B1(_04096_),
    .B2(_03763_),
    .X(_04102_));
 sky130_fd_sc_hd__a22oi_2 _18804_ (.A1(_03889_),
    .A2(\decode.id_ex_imm_reg[13] ),
    .B1(_04101_),
    .B2(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__or2_2 _18805_ (.A(_04100_),
    .B(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__o221a_2 _18806_ (.A1(_04096_),
    .A2(_03699_),
    .B1(_03686_),
    .B2(\decode.id_ex_rs1_data_reg[13] ),
    .C1(_04099_),
    .X(_04105_));
 sky130_fd_sc_hd__a221o_2 _18807_ (.A1(_03890_),
    .A2(\decode.id_ex_imm_reg[13] ),
    .B1(_04101_),
    .B2(_04102_),
    .C1(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__nand2_2 _18808_ (.A(_04104_),
    .B(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__o2bb2a_2 _18809_ (.A1_N(_10039_),
    .A2_N(_10040_),
    .B1(\memory.csr_read_data_out_reg[12] ),
    .B2(_09942_),
    .X(_04108_));
 sky130_fd_sc_hd__or3_2 _18810_ (.A(\execute.csr_read_data_out_reg[12] ),
    .B(_03661_),
    .C(_03660_),
    .X(_04109_));
 sky130_fd_sc_hd__o221a_2 _18811_ (.A1(\execute.io_reg_pc[12] ),
    .A2(_03662_),
    .B1(_03663_),
    .B2(io_memory_address[12]),
    .C1(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__o41a_2 _18812_ (.A1(_03768_),
    .A2(_03769_),
    .A3(_03770_),
    .A4(_04110_),
    .B1(_03669_),
    .X(_04111_));
 sky130_fd_sc_hd__o221a_2 _18813_ (.A1(_04108_),
    .A2(_03914_),
    .B1(_03687_),
    .B2(\decode.id_ex_rs1_data_reg[12] ),
    .C1(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__o221a_2 _18814_ (.A1(_03759_),
    .A2(_04110_),
    .B1(\decode.id_ex_rs2_data_reg[12] ),
    .B2(_03745_),
    .C1(_03726_),
    .X(_04113_));
 sky130_fd_sc_hd__a311o_2 _18815_ (.A1(_03751_),
    .A2(_03752_),
    .A3(_03757_),
    .B1(_03744_),
    .C1(_04108_),
    .X(_04114_));
 sky130_fd_sc_hd__a22oi_2 _18816_ (.A1(_03706_),
    .A2(\decode.id_ex_imm_reg[12] ),
    .B1(_04113_),
    .B2(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__nor2_2 _18817_ (.A(_04112_),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__o221ai_2 _18818_ (.A1(_04108_),
    .A2(_03914_),
    .B1(_03908_),
    .B2(\decode.id_ex_rs1_data_reg[12] ),
    .C1(_04111_),
    .Y(_04117_));
 sky130_fd_sc_hd__inv_2 _18819_ (.A(_04115_),
    .Y(_04118_));
 sky130_fd_sc_hd__nor2_2 _18820_ (.A(_04117_),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__nor2_2 _18821_ (.A(_04116_),
    .B(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hd__or4bb_2 _18822_ (.A(_04086_),
    .B(_04095_),
    .C_N(_04107_),
    .D_N(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__inv_2 _18823_ (.A(_10014_),
    .Y(_04122_));
 sky130_fd_sc_hd__o22a_2 _18824_ (.A1(_03659_),
    .A2(\execute.csr_read_data_out_reg[8] ),
    .B1(\execute.io_reg_pc[8] ),
    .B2(_03777_),
    .X(_04123_));
 sky130_fd_sc_hd__o21ai_2 _18825_ (.A1(io_memory_address[8]),
    .A2(_03666_),
    .B1(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__a21oi_2 _18826_ (.A1(_03817_),
    .A2(_04124_),
    .B1(_03774_),
    .Y(_04125_));
 sky130_fd_sc_hd__o221a_2 _18827_ (.A1(_03688_),
    .A2(\decode.id_ex_rs1_data_reg[8] ),
    .B1(_03700_),
    .B2(_04122_),
    .C1(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__a21oi_2 _18828_ (.A1(_03797_),
    .A2(_04124_),
    .B1(_03890_),
    .Y(_04127_));
 sky130_fd_sc_hd__o22a_2 _18829_ (.A1(\decode.id_ex_rs2_data_reg[8] ),
    .A2(_03746_),
    .B1(_03764_),
    .B2(_04122_),
    .X(_04128_));
 sky130_fd_sc_hd__a22oi_2 _18830_ (.A1(_03890_),
    .A2(\decode.id_ex_imm_reg[8] ),
    .B1(_04127_),
    .B2(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__nor2_2 _18831_ (.A(_04126_),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__and2_2 _18832_ (.A(_04126_),
    .B(_04129_),
    .X(_04131_));
 sky130_fd_sc_hd__nor2_2 _18833_ (.A(_04130_),
    .B(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__o22a_2 _18834_ (.A1(\memory.csr_read_data_out_reg[9] ),
    .A2(_10010_),
    .B1(_10022_),
    .B2(_10023_),
    .X(_04133_));
 sky130_fd_sc_hd__o22a_2 _18835_ (.A1(_03658_),
    .A2(\execute.csr_read_data_out_reg[9] ),
    .B1(\execute.io_reg_pc[9] ),
    .B2(_03662_),
    .X(_04134_));
 sky130_fd_sc_hd__o21ai_2 _18836_ (.A1(io_memory_address[9]),
    .A2(_03664_),
    .B1(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__a21oi_2 _18837_ (.A1(_03816_),
    .A2(_04135_),
    .B1(_03773_),
    .Y(_04136_));
 sky130_fd_sc_hd__o221a_2 _18838_ (.A1(_04133_),
    .A2(_03914_),
    .B1(_03687_),
    .B2(\decode.id_ex_rs1_data_reg[9] ),
    .C1(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__or3b_2 _18839_ (.A(_03715_),
    .B(_03725_),
    .C_N(_04135_),
    .X(_04138_));
 sky130_fd_sc_hd__o221ai_2 _18840_ (.A1(\decode.id_ex_rs2_data_reg[9] ),
    .A2(_03745_),
    .B1(_03763_),
    .B2(_04133_),
    .C1(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__nand2_2 _18841_ (.A(_03889_),
    .B(\decode.id_ex_imm_reg[9] ),
    .Y(_04140_));
 sky130_fd_sc_hd__o21a_2 _18842_ (.A1(_03707_),
    .A2(_04139_),
    .B1(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__nor2_2 _18843_ (.A(_04137_),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__o211a_2 _18844_ (.A1(_03890_),
    .A2(_04139_),
    .B1(_04140_),
    .C1(_04137_),
    .X(_04143_));
 sky130_fd_sc_hd__nor2_2 _18845_ (.A(_04142_),
    .B(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__o22a_2 _18846_ (.A1(\memory.csr_read_data_out_reg[11] ),
    .A2(_10010_),
    .B1(_10033_),
    .B2(_10034_),
    .X(_04145_));
 sky130_fd_sc_hd__o22a_2 _18847_ (.A1(_03658_),
    .A2(\execute.csr_read_data_out_reg[11] ),
    .B1(\execute.io_reg_pc[11] ),
    .B2(_03662_),
    .X(_04146_));
 sky130_fd_sc_hd__o21ai_2 _18848_ (.A1(io_memory_address[11]),
    .A2(_03664_),
    .B1(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__a21oi_2 _18849_ (.A1(_03816_),
    .A2(_04147_),
    .B1(_03773_),
    .Y(_04148_));
 sky130_fd_sc_hd__o221a_2 _18850_ (.A1(_04145_),
    .A2(_03699_),
    .B1(_03687_),
    .B2(\decode.id_ex_rs1_data_reg[11] ),
    .C1(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__a21oi_2 _18851_ (.A1(_03796_),
    .A2(_04147_),
    .B1(_03706_),
    .Y(_04150_));
 sky130_fd_sc_hd__o221a_2 _18852_ (.A1(\decode.id_ex_rs2_data_reg[11] ),
    .A2(_03745_),
    .B1(_04145_),
    .B2(_03763_),
    .C1(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__a21oi_2 _18853_ (.A1(_03707_),
    .A2(\decode.id_ex_imm_reg[11] ),
    .B1(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__nand2_2 _18854_ (.A(_04149_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__or2_2 _18855_ (.A(_04149_),
    .B(_04152_),
    .X(_04154_));
 sky130_fd_sc_hd__and2_2 _18856_ (.A(_04153_),
    .B(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__o22a_2 _18857_ (.A1(\memory.csr_read_data_out_reg[10] ),
    .A2(_10010_),
    .B1(_10028_),
    .B2(_10029_),
    .X(_04156_));
 sky130_fd_sc_hd__o22a_2 _18858_ (.A1(_03658_),
    .A2(\execute.csr_read_data_out_reg[10] ),
    .B1(\execute.io_reg_pc[10] ),
    .B2(_03776_),
    .X(_04157_));
 sky130_fd_sc_hd__o21ai_2 _18859_ (.A1(io_memory_address[10]),
    .A2(_03665_),
    .B1(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__a21oi_2 _18860_ (.A1(_03816_),
    .A2(_04158_),
    .B1(_03773_),
    .Y(_04159_));
 sky130_fd_sc_hd__o221ai_2 _18861_ (.A1(\decode.id_ex_rs1_data_reg[10] ),
    .A2(_03908_),
    .B1(_04156_),
    .B2(_03700_),
    .C1(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__a311o_2 _18862_ (.A1(_03751_),
    .A2(_03752_),
    .A3(_03757_),
    .B1(_03744_),
    .C1(_04156_),
    .X(_04161_));
 sky130_fd_sc_hd__nand2_2 _18863_ (.A(_03796_),
    .B(_04158_),
    .Y(_04162_));
 sky130_fd_sc_hd__o311a_2 _18864_ (.A1(\decode.id_ex_rs2_data_reg[10] ),
    .A2(_03796_),
    .A3(_03784_),
    .B1(_04162_),
    .C1(_03727_),
    .X(_04163_));
 sky130_fd_sc_hd__a22oi_2 _18865_ (.A1(_03707_),
    .A2(\decode.id_ex_imm_reg[10] ),
    .B1(_04161_),
    .B2(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__or2_2 _18866_ (.A(_04160_),
    .B(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__o221a_2 _18867_ (.A1(\decode.id_ex_rs1_data_reg[10] ),
    .A2(_03687_),
    .B1(_04156_),
    .B2(_03914_),
    .C1(_04159_),
    .X(_04166_));
 sky130_fd_sc_hd__a221o_2 _18868_ (.A1(_03708_),
    .A2(\decode.id_ex_imm_reg[10] ),
    .B1(_04161_),
    .B2(_04163_),
    .C1(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__nand2_2 _18869_ (.A(_04165_),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__nand4_2 _18870_ (.A(_04132_),
    .B(_04144_),
    .C(_04155_),
    .D(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__or2_2 _18871_ (.A(_04121_),
    .B(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__nor2_2 _18872_ (.A(_04062_),
    .B(_04065_),
    .Y(_04171_));
 sky130_fd_sc_hd__nand2_2 _18873_ (.A(_04070_),
    .B(_04073_),
    .Y(_04172_));
 sky130_fd_sc_hd__and2_2 _18874_ (.A(_04062_),
    .B(_04065_),
    .X(_04173_));
 sky130_fd_sc_hd__o21bai_2 _18875_ (.A1(_04171_),
    .A2(_04172_),
    .B1_N(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__a311o_2 _18876_ (.A1(_04053_),
    .A2(_04057_),
    .A3(_04076_),
    .B1(_04170_),
    .C1(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__o21ai_2 _18877_ (.A1(_04166_),
    .A2(_04164_),
    .B1(_04154_),
    .Y(_04176_));
 sky130_fd_sc_hd__nand2_2 _18878_ (.A(_04137_),
    .B(_04141_),
    .Y(_04177_));
 sky130_fd_sc_hd__o2111a_2 _18879_ (.A1(_04130_),
    .A2(_04142_),
    .B1(_04177_),
    .C1(_04168_),
    .D1(_04155_),
    .X(_04178_));
 sky130_fd_sc_hd__a21oi_2 _18880_ (.A1(_04153_),
    .A2(_04176_),
    .B1(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__o221a_2 _18881_ (.A1(_04087_),
    .A2(_03701_),
    .B1(_03688_),
    .B2(\decode.id_ex_rs1_data_reg[15] ),
    .C1(_04090_),
    .X(_04180_));
 sky130_fd_sc_hd__o221a_2 _18882_ (.A1(_04077_),
    .A2(_03701_),
    .B1(_03689_),
    .B2(\decode.id_ex_rs1_data_reg[14] ),
    .C1(_04080_),
    .X(_04181_));
 sky130_fd_sc_hd__and2_2 _18883_ (.A(_04083_),
    .B(_04084_),
    .X(_04182_));
 sky130_fd_sc_hd__o22a_2 _18884_ (.A1(_04181_),
    .A2(_04182_),
    .B1(_04180_),
    .B2(_04094_),
    .X(_04183_));
 sky130_fd_sc_hd__a21o_2 _18885_ (.A1(_04180_),
    .A2(_04094_),
    .B1(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__o22a_2 _18886_ (.A1(_04112_),
    .A2(_04115_),
    .B1(_04105_),
    .B2(_04103_),
    .X(_04185_));
 sky130_fd_sc_hd__buf_1 _18887_ (.A(_04086_),
    .X(_04186_));
 sky130_fd_sc_hd__a2111o_2 _18888_ (.A1(_04105_),
    .A2(_04103_),
    .B1(_04185_),
    .C1(_04186_),
    .D1(_04095_),
    .X(_04187_));
 sky130_fd_sc_hd__o211a_2 _18889_ (.A1(_04121_),
    .A2(_04179_),
    .B1(_04184_),
    .C1(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__nor2_2 _18890_ (.A(_03888_),
    .B(_03893_),
    .Y(_04189_));
 sky130_fd_sc_hd__nor2_2 _18891_ (.A(_04189_),
    .B(_03894_),
    .Y(_04190_));
 sky130_fd_sc_hd__nand2b_2 _18892_ (.A_N(_03948_),
    .B(_03962_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2b_2 _18893_ (.A_N(_03957_),
    .B(_03960_),
    .Y(_04192_));
 sky130_fd_sc_hd__nor2_2 _18894_ (.A(_04191_),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__nor2_2 _18895_ (.A(_03872_),
    .B(_03881_),
    .Y(_04194_));
 sky130_fd_sc_hd__nor2_2 _18896_ (.A(_04194_),
    .B(_03882_),
    .Y(_04195_));
 sky130_fd_sc_hd__and3_2 _18897_ (.A(_04190_),
    .B(_04193_),
    .C(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__a221oi_2 _18898_ (.A1(_03890_),
    .A2(\decode.id_ex_imm_reg[17] ),
    .B1(_03906_),
    .B2(_03907_),
    .C1(_03934_),
    .Y(_04197_));
 sky130_fd_sc_hd__nor2_2 _18899_ (.A(_03911_),
    .B(_03935_),
    .Y(_04198_));
 sky130_fd_sc_hd__o221ai_2 _18900_ (.A1(\decode.id_ex_rs1_data_reg[18] ),
    .A2(_03908_),
    .B1(_03913_),
    .B2(_03700_),
    .C1(_03917_),
    .Y(_04199_));
 sky130_fd_sc_hd__a31o_2 _18901_ (.A1(_03919_),
    .A2(_03920_),
    .A3(_03921_),
    .B1(_03922_),
    .X(_04200_));
 sky130_fd_sc_hd__nor2_2 _18902_ (.A(_04199_),
    .B(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__nor2_2 _18903_ (.A(_04201_),
    .B(_03938_),
    .Y(_04202_));
 sky130_fd_sc_hd__a21oi_2 _18904_ (.A1(_03890_),
    .A2(\decode.id_ex_imm_reg[19] ),
    .B1(_03898_),
    .Y(_04203_));
 sky130_fd_sc_hd__nand2_2 _18905_ (.A(_04203_),
    .B(_03902_),
    .Y(_04204_));
 sky130_fd_sc_hd__o221a_2 _18906_ (.A1(_03900_),
    .A2(_03914_),
    .B1(_03908_),
    .B2(\decode.id_ex_rs1_data_reg[19] ),
    .C1(_03901_),
    .X(_04205_));
 sky130_fd_sc_hd__o21ai_2 _18907_ (.A1(_03898_),
    .A2(_03899_),
    .B1(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__nand2_2 _18908_ (.A(_04204_),
    .B(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__nor2_2 _18909_ (.A(_03929_),
    .B(_03933_),
    .Y(_04208_));
 sky130_fd_sc_hd__o221ai_2 _18910_ (.A1(\decode.id_ex_rs1_data_reg[16] ),
    .A2(_03688_),
    .B1(_03925_),
    .B2(_03701_),
    .C1(_03928_),
    .Y(_04209_));
 sky130_fd_sc_hd__a211o_2 _18911_ (.A1(_03708_),
    .A2(\decode.id_ex_imm_reg[16] ),
    .B1(_04209_),
    .C1(_03932_),
    .X(_04210_));
 sky130_fd_sc_hd__nor2b_2 _18912_ (.A(_04208_),
    .B_N(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__o2111a_2 _18913_ (.A1(_04197_),
    .A2(_04198_),
    .B1(_04202_),
    .C1(_04207_),
    .D1(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__nand2_2 _18914_ (.A(_04196_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__a211o_2 _18915_ (.A1(_04175_),
    .A2(_04188_),
    .B1(_03867_),
    .C1(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__or2_2 _18916_ (.A(_03863_),
    .B(_03861_),
    .X(_04215_));
 sky130_fd_sc_hd__a211o_2 _18917_ (.A1(_03835_),
    .A2(_03838_),
    .B1(_03844_),
    .C1(_03847_),
    .X(_04216_));
 sky130_fd_sc_hd__o221a_2 _18918_ (.A1(_03835_),
    .A2(_03838_),
    .B1(_03821_),
    .B2(_03825_),
    .C1(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__o21a_2 _18919_ (.A1(_03812_),
    .A2(_03809_),
    .B1(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__a21oi_2 _18920_ (.A1(_03811_),
    .A2(_03827_),
    .B1(_03826_),
    .Y(_04219_));
 sky130_fd_sc_hd__a211o_2 _18921_ (.A1(_03795_),
    .A2(_03800_),
    .B1(_04218_),
    .C1(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__o22a_2 _18922_ (.A1(_03781_),
    .A2(_03788_),
    .B1(_03795_),
    .B2(_03800_),
    .X(_04221_));
 sky130_fd_sc_hd__a211o_2 _18923_ (.A1(_04220_),
    .A2(_04221_),
    .B1(_03790_),
    .C1(_03862_),
    .X(_04222_));
 sky130_fd_sc_hd__and4_2 _18924_ (.A(_04214_),
    .B(_03854_),
    .C(_04215_),
    .D(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__o31a_2 _18925_ (.A1(_03867_),
    .A2(_03882_),
    .A3(_03965_),
    .B1(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__buf_1 _18926_ (.A(_03637_),
    .X(_04225_));
 sky130_fd_sc_hd__and2_2 _18927_ (.A(_04075_),
    .B(_04172_),
    .X(_04226_));
 sky130_fd_sc_hd__nor2_2 _18928_ (.A(_04171_),
    .B(_04173_),
    .Y(_04227_));
 sky130_fd_sc_hd__o2bb2ai_2 _18929_ (.A1_N(_03997_),
    .A2_N(_03998_),
    .B1(_03999_),
    .B2(_04002_),
    .Y(_04228_));
 sky130_fd_sc_hd__nand3_2 _18930_ (.A(_03977_),
    .B(_03979_),
    .C(_03982_),
    .Y(_04229_));
 sky130_fd_sc_hd__a31o_2 _18931_ (.A1(_03984_),
    .A2(_03985_),
    .A3(_03986_),
    .B1(_03987_),
    .X(_04230_));
 sky130_fd_sc_hd__a21o_2 _18932_ (.A1(_03670_),
    .A2(_04229_),
    .B1(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__and3_2 _18933_ (.A(_04006_),
    .B(_04228_),
    .C(_04231_),
    .X(_04232_));
 sky130_fd_sc_hd__buf_1 _18934_ (.A(_03988_),
    .X(_04233_));
 sky130_fd_sc_hd__buf_1 _18935_ (.A(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__a311o_2 _18936_ (.A1(_03977_),
    .A2(_03979_),
    .A3(_03982_),
    .B1(_04234_),
    .C1(_03775_),
    .X(_04235_));
 sky130_fd_sc_hd__and4_2 _18937_ (.A(_04226_),
    .B(_04227_),
    .C(_04232_),
    .D(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__and4_2 _18938_ (.A(_04052_),
    .B(_04039_),
    .C(_04025_),
    .D(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__or4b_2 _18939_ (.A(_03867_),
    .B(_04213_),
    .C(_04170_),
    .D_N(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__o31a_2 _18940_ (.A1(_04225_),
    .A2(_03705_),
    .A3(_03766_),
    .B1(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__or4b_2 _18941_ (.A(_03636_),
    .B(_03767_),
    .C(_04224_),
    .D_N(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__and3b_2 _18942_ (.A_N(_03635_),
    .B(_03634_),
    .C(_03633_),
    .X(_04241_));
 sky130_fd_sc_hd__buf_1 _18943_ (.A(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__buf_1 _18944_ (.A(_04028_),
    .X(_04243_));
 sky130_fd_sc_hd__buf_1 _18945_ (.A(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__buf_1 _18946_ (.A(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__a32o_2 _18947_ (.A1(_03990_),
    .A2(_03991_),
    .A3(_03996_),
    .B1(_03706_),
    .B2(\decode.id_ex_imm_reg[1] ),
    .X(_04246_));
 sky130_fd_sc_hd__buf_1 _18948_ (.A(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__buf_1 _18949_ (.A(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__buf_1 _18950_ (.A(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__mux2_2 _18951_ (.A0(_04209_),
    .A1(_03911_),
    .S(_03989_),
    .X(_04250_));
 sky130_fd_sc_hd__buf_1 _18952_ (.A(_03997_),
    .X(_04251_));
 sky130_fd_sc_hd__buf_1 _18953_ (.A(_03998_),
    .X(_04252_));
 sky130_fd_sc_hd__buf_1 _18954_ (.A(_04233_),
    .X(_04253_));
 sky130_fd_sc_hd__buf_1 _18955_ (.A(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__buf_1 _18956_ (.A(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__a311o_2 _18957_ (.A1(_03986_),
    .A2(_03985_),
    .A3(_03984_),
    .B1(_03987_),
    .C1(_04205_),
    .X(_04256_));
 sky130_fd_sc_hd__o21ai_2 _18958_ (.A1(_03918_),
    .A2(_04255_),
    .B1(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__a21o_2 _18959_ (.A1(_04251_),
    .A2(_04252_),
    .B1(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__o21ai_2 _18960_ (.A1(_04249_),
    .A2(_04250_),
    .B1(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__mux2_2 _18961_ (.A0(_03888_),
    .A1(_03872_),
    .S(_04233_),
    .X(_04260_));
 sky130_fd_sc_hd__buf_1 _18962_ (.A(\decode.id_ex_imm_reg[1] ),
    .X(_04261_));
 sky130_fd_sc_hd__and3_2 _18963_ (.A(_03990_),
    .B(_03991_),
    .C(_03996_),
    .X(_04262_));
 sky130_fd_sc_hd__buf_1 _18964_ (.A(_04262_),
    .X(_04263_));
 sky130_fd_sc_hd__a21oi_2 _18965_ (.A1(_03709_),
    .A2(_04261_),
    .B1(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__a311o_2 _18966_ (.A1(_03986_),
    .A2(_03985_),
    .A3(_03984_),
    .B1(_03987_),
    .C1(_03944_),
    .X(_04265_));
 sky130_fd_sc_hd__o211a_2 _18967_ (.A1(_03956_),
    .A2(_04253_),
    .B1(_04264_),
    .C1(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__a21o_2 _18968_ (.A1(_04260_),
    .A2(_04247_),
    .B1(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__a31o_2 _18969_ (.A1(_04015_),
    .A2(_04016_),
    .A3(_04017_),
    .B1(_04019_),
    .X(_04268_));
 sky130_fd_sc_hd__buf_1 _18970_ (.A(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__buf_1 _18971_ (.A(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__mux2_2 _18972_ (.A0(_04259_),
    .A1(_04267_),
    .S(_04270_),
    .X(_04271_));
 sky130_fd_sc_hd__buf_1 _18973_ (.A(_04021_),
    .X(_04272_));
 sky130_fd_sc_hd__buf_1 _18974_ (.A(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__buf_1 _18975_ (.A(_04230_),
    .X(_04274_));
 sky130_fd_sc_hd__mux2_2 _18976_ (.A0(_03821_),
    .A1(_03812_),
    .S(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__mux2_2 _18977_ (.A0(_03835_),
    .A1(_03844_),
    .S(_04230_),
    .X(_04276_));
 sky130_fd_sc_hd__buf_1 _18978_ (.A(_04264_),
    .X(_04277_));
 sky130_fd_sc_hd__mux2_2 _18979_ (.A0(_04275_),
    .A1(_04276_),
    .S(_04277_),
    .X(_04278_));
 sky130_fd_sc_hd__o221a_2 _18980_ (.A1(\decode.id_ex_rs2_data_reg[2] ),
    .A2(_03745_),
    .B1(_04010_),
    .B2(_04046_),
    .C1(_04015_),
    .X(_04279_));
 sky130_fd_sc_hd__buf_1 _18981_ (.A(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__buf_1 _18982_ (.A(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__buf_1 _18983_ (.A(_04019_),
    .X(_04282_));
 sky130_fd_sc_hd__buf_1 _18984_ (.A(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__mux2_2 _18985_ (.A0(_03795_),
    .A1(_03781_),
    .S(_04253_),
    .X(_04284_));
 sky130_fd_sc_hd__or2_2 _18986_ (.A(_03863_),
    .B(_04254_),
    .X(_04285_));
 sky130_fd_sc_hd__a311o_2 _18987_ (.A1(_03986_),
    .A2(_03985_),
    .A3(_03984_),
    .B1(_03987_),
    .C1(_03703_),
    .X(_04286_));
 sky130_fd_sc_hd__a22o_2 _18988_ (.A1(_04251_),
    .A2(_04252_),
    .B1(_04285_),
    .B2(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__o221a_2 _18989_ (.A1(_04281_),
    .A2(_04283_),
    .B1(_04249_),
    .B2(_04284_),
    .C1(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__buf_1 _18990_ (.A(_03975_),
    .X(_04289_));
 sky130_fd_sc_hd__buf_1 _18991_ (.A(_04289_),
    .X(_04290_));
 sky130_fd_sc_hd__buf_1 _18992_ (.A(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__a211o_2 _18993_ (.A1(_04273_),
    .A2(_04278_),
    .B1(_04288_),
    .C1(_04291_),
    .X(_04292_));
 sky130_fd_sc_hd__o21ai_2 _18994_ (.A1(_04245_),
    .A2(_04271_),
    .B1(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__buf_1 _18995_ (.A(_04038_),
    .X(_04294_));
 sky130_fd_sc_hd__buf_1 _18996_ (.A(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__or3_2 _18997_ (.A(_04255_),
    .B(_03983_),
    .C(_04248_),
    .X(_04296_));
 sky130_fd_sc_hd__buf_1 _18998_ (.A(_03709_),
    .X(_04297_));
 sky130_fd_sc_hd__o22a_2 _18999_ (.A1(\decode.id_ex_rs2_data_reg[4] ),
    .A2(_03747_),
    .B1(_04030_),
    .B2(_03764_),
    .X(_04298_));
 sky130_fd_sc_hd__inv_2 _19000_ (.A(\decode.id_ex_aluop_reg[0] ),
    .Y(_04299_));
 sky130_fd_sc_hd__or4b_2 _19001_ (.A(_04299_),
    .B(\decode.id_ex_aluop_reg[1] ),
    .C(\decode.id_ex_aluop_reg[3] ),
    .D_N(\decode.id_ex_aluop_reg[2] ),
    .X(_04300_));
 sky130_fd_sc_hd__buf_1 _19002_ (.A(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__a221o_2 _19003_ (.A1(_04297_),
    .A2(\decode.id_ex_imm_reg[4] ),
    .B1(_04035_),
    .B2(_04298_),
    .C1(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__buf_1 _19004_ (.A(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__or3_2 _19005_ (.A(_04279_),
    .B(_04019_),
    .C(_04028_),
    .X(_04304_));
 sky130_fd_sc_hd__buf_1 _19006_ (.A(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__nand3b_2 _19007_ (.A_N(_03635_),
    .B(_03634_),
    .C(_03633_),
    .Y(_04306_));
 sky130_fd_sc_hd__buf_1 _19008_ (.A(_04274_),
    .X(_04307_));
 sky130_fd_sc_hd__or4b_2 _19009_ (.A(_03637_),
    .B(_03633_),
    .C(_03635_),
    .D_N(_03634_),
    .X(_04308_));
 sky130_fd_sc_hd__o211ai_2 _19010_ (.A1(_09949_),
    .A2(_04046_),
    .B1(_03985_),
    .C1(_03984_),
    .Y(_04309_));
 sky130_fd_sc_hd__o2111a_2 _19011_ (.A1(\decode.id_ex_imm_reg[0] ),
    .A2(_03726_),
    .B1(_03669_),
    .C1(_04229_),
    .D1(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__or3b_2 _19012_ (.A(\decode.id_ex_aluop_reg[3] ),
    .B(\decode.id_ex_aluop_reg[2] ),
    .C_N(\decode.id_ex_aluop_reg[1] ),
    .X(_04311_));
 sky130_fd_sc_hd__o32a_2 _19013_ (.A1(_03635_),
    .A2(_03634_),
    .A3(_04310_),
    .B1(_04311_),
    .B2(_04299_),
    .X(_04312_));
 sky130_fd_sc_hd__a21o_2 _19014_ (.A1(_03983_),
    .A2(_04307_),
    .B1(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__o31a_2 _19015_ (.A1(_03983_),
    .A2(_04307_),
    .A3(_04308_),
    .B1(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__o311a_2 _19016_ (.A1(_04296_),
    .A2(_04303_),
    .A3(_04305_),
    .B1(_04306_),
    .C1(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__o211a_2 _19017_ (.A1(_03972_),
    .A2(_03974_),
    .B1(_04007_),
    .C1(_04021_),
    .X(_04316_));
 sky130_fd_sc_hd__buf_1 _19018_ (.A(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__o221a_2 _19019_ (.A1(\decode.id_ex_imm_reg[0] ),
    .A2(_03728_),
    .B1(_03999_),
    .B2(_04002_),
    .C1(_04309_),
    .X(_04318_));
 sky130_fd_sc_hd__a211o_2 _19020_ (.A1(_03983_),
    .A2(_04307_),
    .B1(_04249_),
    .C1(_04318_),
    .X(_04319_));
 sky130_fd_sc_hd__buf_1 _19021_ (.A(_04255_),
    .X(_04320_));
 sky130_fd_sc_hd__buf_1 _19022_ (.A(_04014_),
    .X(_04321_));
 sky130_fd_sc_hd__o21ai_2 _19023_ (.A1(_04321_),
    .A2(_04255_),
    .B1(_04248_),
    .Y(_04322_));
 sky130_fd_sc_hd__a21o_2 _19024_ (.A1(_04027_),
    .A2(_04320_),
    .B1(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__buf_1 _19025_ (.A(_04264_),
    .X(_04324_));
 sky130_fd_sc_hd__buf_1 _19026_ (.A(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__mux2_2 _19027_ (.A0(_04045_),
    .A1(_04054_),
    .S(_04307_),
    .X(_04326_));
 sky130_fd_sc_hd__a311o_2 _19028_ (.A1(_03986_),
    .A2(_03985_),
    .A3(_03984_),
    .B1(_03987_),
    .C1(_04062_),
    .X(_04327_));
 sky130_fd_sc_hd__o211a_2 _19029_ (.A1(_04320_),
    .A2(_04070_),
    .B1(_04327_),
    .C1(_04249_),
    .X(_04328_));
 sky130_fd_sc_hd__a21oi_2 _19030_ (.A1(_04325_),
    .A2(_04326_),
    .B1(_04328_),
    .Y(_04329_));
 sky130_fd_sc_hd__o211a_2 _19031_ (.A1(_03972_),
    .A2(_03974_),
    .B1(_04007_),
    .C1(_04268_),
    .X(_04330_));
 sky130_fd_sc_hd__a32o_2 _19032_ (.A1(_04317_),
    .A2(_04319_),
    .A3(_04323_),
    .B1(_04329_),
    .B2(_04330_),
    .X(_04331_));
 sky130_fd_sc_hd__buf_1 _19033_ (.A(_04248_),
    .X(_04332_));
 sky130_fd_sc_hd__mux2_2 _19034_ (.A0(_04126_),
    .A1(_04137_),
    .S(_04255_),
    .X(_04333_));
 sky130_fd_sc_hd__o221ai_2 _19035_ (.A1(\decode.id_ex_rs1_data_reg[11] ),
    .A2(_03689_),
    .B1(_04145_),
    .B2(_03701_),
    .C1(_04148_),
    .Y(_04334_));
 sky130_fd_sc_hd__mux2_2 _19036_ (.A0(_04160_),
    .A1(_04334_),
    .S(_03989_),
    .X(_04335_));
 sky130_fd_sc_hd__nand2_2 _19037_ (.A(_04249_),
    .B(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__o21ai_2 _19038_ (.A1(_04332_),
    .A2(_04333_),
    .B1(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__buf_1 _19039_ (.A(_04324_),
    .X(_04338_));
 sky130_fd_sc_hd__mux2_2 _19040_ (.A0(_04081_),
    .A1(_04091_),
    .S(_03989_),
    .X(_04339_));
 sky130_fd_sc_hd__mux2_2 _19041_ (.A0(_04117_),
    .A1(_04100_),
    .S(_03989_),
    .X(_04340_));
 sky130_fd_sc_hd__a211o_2 _19042_ (.A1(_04297_),
    .A2(_04261_),
    .B1(_04263_),
    .C1(_04340_),
    .X(_04341_));
 sky130_fd_sc_hd__o21ai_2 _19043_ (.A1(_04338_),
    .A2(_04339_),
    .B1(_04341_),
    .Y(_04342_));
 sky130_fd_sc_hd__o21ai_2 _19044_ (.A1(_04281_),
    .A2(_04283_),
    .B1(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__o311a_2 _19045_ (.A1(_04281_),
    .A2(_04337_),
    .A3(_04283_),
    .B1(_04244_),
    .C1(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__buf_1 _19046_ (.A(_04056_),
    .X(_04345_));
 sky130_fd_sc_hd__buf_1 _19047_ (.A(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__o211a_2 _19048_ (.A1(_04331_),
    .A2(_04344_),
    .B1(_04242_),
    .C1(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__a311o_2 _19049_ (.A1(_04242_),
    .A2(_04293_),
    .A3(_04295_),
    .B1(_04315_),
    .C1(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__a21oi_2 _19050_ (.A1(_04240_),
    .A2(_04348_),
    .B1(_03588_),
    .Y(_00548_));
 sky130_fd_sc_hd__buf_1 _19051_ (.A(_04290_),
    .X(_04349_));
 sky130_fd_sc_hd__mux2_2 _19052_ (.A0(_03888_),
    .A1(_03944_),
    .S(_04230_),
    .X(_04350_));
 sky130_fd_sc_hd__mux2_2 _19053_ (.A0(_03872_),
    .A1(_03844_),
    .S(_03989_),
    .X(_04351_));
 sky130_fd_sc_hd__buf_1 _19054_ (.A(_04246_),
    .X(_04352_));
 sky130_fd_sc_hd__mux2_2 _19055_ (.A0(_04350_),
    .A1(_04351_),
    .S(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__mux2_2 _19056_ (.A0(_04205_),
    .A1(_03956_),
    .S(_04233_),
    .X(_04354_));
 sky130_fd_sc_hd__mux2_2 _19057_ (.A0(_03934_),
    .A1(_03918_),
    .S(_03989_),
    .X(_04355_));
 sky130_fd_sc_hd__mux2_2 _19058_ (.A0(_04354_),
    .A1(_04355_),
    .S(_04324_),
    .X(_04356_));
 sky130_fd_sc_hd__mux2_2 _19059_ (.A0(_04353_),
    .A1(_04356_),
    .S(_04272_),
    .X(_04357_));
 sky130_fd_sc_hd__a311o_2 _19060_ (.A1(_03863_),
    .A2(_04251_),
    .A3(_04252_),
    .B1(_04307_),
    .C1(_04272_),
    .X(_04358_));
 sky130_fd_sc_hd__buf_1 _19061_ (.A(_04299_),
    .X(_04359_));
 sky130_fd_sc_hd__nand2_2 _19062_ (.A(_04242_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__a2111o_2 _19063_ (.A1(_04349_),
    .A2(_04357_),
    .B1(_04358_),
    .C1(_04360_),
    .D1(_04346_),
    .X(_04361_));
 sky130_fd_sc_hd__buf_1 _19064_ (.A(_04306_),
    .X(_04362_));
 sky130_fd_sc_hd__mux2_2 _19065_ (.A0(_03821_),
    .A1(_03795_),
    .S(_03988_),
    .X(_04363_));
 sky130_fd_sc_hd__mux2_2 _19066_ (.A0(_03835_),
    .A1(_03812_),
    .S(_03989_),
    .X(_04364_));
 sky130_fd_sc_hd__mux2_2 _19067_ (.A0(_04363_),
    .A1(_04364_),
    .S(_04277_),
    .X(_04365_));
 sky130_fd_sc_hd__a2111oi_2 _19068_ (.A1(_03772_),
    .A2(_10135_),
    .B1(_03775_),
    .C1(_03780_),
    .D1(_03988_),
    .Y(_04366_));
 sky130_fd_sc_hd__a21o_2 _19069_ (.A1(_03863_),
    .A2(_04233_),
    .B1(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__mux2_2 _19070_ (.A0(_04367_),
    .A1(_03704_),
    .S(_04247_),
    .X(_04368_));
 sky130_fd_sc_hd__mux2_2 _19071_ (.A0(_04365_),
    .A1(_04368_),
    .S(_04269_),
    .X(_04369_));
 sky130_fd_sc_hd__mux2_2 _19072_ (.A0(_04369_),
    .A1(_04357_),
    .S(_04291_),
    .X(_04370_));
 sky130_fd_sc_hd__buf_1 _19073_ (.A(_04290_),
    .X(_04371_));
 sky130_fd_sc_hd__mux4_2 _19074_ (.A0(_04062_),
    .A1(_04126_),
    .A2(_04045_),
    .A3(_04070_),
    .S0(_04320_),
    .S1(_04325_),
    .X(_04372_));
 sky130_fd_sc_hd__o211a_2 _19075_ (.A1(\decode.id_ex_rs1_data_reg[1] ),
    .A2(_03686_),
    .B1(_04005_),
    .C1(_04001_),
    .X(_04373_));
 sky130_fd_sc_hd__mux4_2 _19076_ (.A0(_04054_),
    .A1(_03971_),
    .A2(_04321_),
    .A3(_04373_),
    .S0(_04307_),
    .S1(_04338_),
    .X(_04374_));
 sky130_fd_sc_hd__mux2_2 _19077_ (.A0(_04334_),
    .A1(_04117_),
    .S(_04233_),
    .X(_04375_));
 sky130_fd_sc_hd__o221ai_2 _19078_ (.A1(\decode.id_ex_rs1_data_reg[9] ),
    .A2(_03689_),
    .B1(_04133_),
    .B2(_03701_),
    .C1(_04136_),
    .Y(_04376_));
 sky130_fd_sc_hd__mux2_2 _19079_ (.A0(_04376_),
    .A1(_04160_),
    .S(_04254_),
    .X(_04377_));
 sky130_fd_sc_hd__mux2_2 _19080_ (.A0(_04375_),
    .A1(_04377_),
    .S(_04324_),
    .X(_04378_));
 sky130_fd_sc_hd__mux2_2 _19081_ (.A0(_04105_),
    .A1(_04181_),
    .S(_04233_),
    .X(_04379_));
 sky130_fd_sc_hd__nand2_2 _19082_ (.A(_04233_),
    .B(_04209_),
    .Y(_04380_));
 sky130_fd_sc_hd__o21a_2 _19083_ (.A1(_04233_),
    .A2(_04180_),
    .B1(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__mux2_2 _19084_ (.A0(_04379_),
    .A1(_04381_),
    .S(_04352_),
    .X(_04382_));
 sky130_fd_sc_hd__o21ai_2 _19085_ (.A1(_04280_),
    .A2(_04282_),
    .B1(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__o21ai_2 _19086_ (.A1(_04269_),
    .A2(_04378_),
    .B1(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__a22o_2 _19087_ (.A1(_04316_),
    .A2(_04374_),
    .B1(_04384_),
    .B2(_04243_),
    .X(_04385_));
 sky130_fd_sc_hd__a221o_2 _19088_ (.A1(_04297_),
    .A2(\decode.id_ex_imm_reg[4] ),
    .B1(_04035_),
    .B2(_04298_),
    .C1(_04306_),
    .X(_04386_));
 sky130_fd_sc_hd__a311o_2 _19089_ (.A1(_04371_),
    .A2(_04270_),
    .A3(_04372_),
    .B1(_04385_),
    .C1(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__or4b_2 _19090_ (.A(_03635_),
    .B(_03634_),
    .C(_04299_),
    .D_N(_03633_),
    .X(_04388_));
 sky130_fd_sc_hd__nand2_2 _19091_ (.A(_04246_),
    .B(_04373_),
    .Y(_04389_));
 sky130_fd_sc_hd__o221ai_2 _19092_ (.A1(_04325_),
    .A2(_04388_),
    .B1(_04308_),
    .B2(_04389_),
    .C1(_04306_),
    .Y(_04390_));
 sky130_fd_sc_hd__nor3b_2 _19093_ (.A(\decode.id_ex_aluop_reg[1] ),
    .B(\decode.id_ex_aluop_reg[3] ),
    .C_N(\decode.id_ex_aluop_reg[2] ),
    .Y(_04391_));
 sky130_fd_sc_hd__and3_2 _19094_ (.A(_03637_),
    .B(_04056_),
    .C(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__o211a_2 _19095_ (.A1(_04373_),
    .A2(_04255_),
    .B1(_04338_),
    .C1(_04231_),
    .X(_04393_));
 sky130_fd_sc_hd__nor3b_2 _19096_ (.A(_03635_),
    .B(\decode.id_ex_aluop_reg[2] ),
    .C_N(_03633_),
    .Y(_04394_));
 sky130_fd_sc_hd__o2111ai_2 _19097_ (.A1(_03816_),
    .A2(_04000_),
    .B1(_04005_),
    .C1(_04001_),
    .D1(_03998_),
    .Y(_04395_));
 sky130_fd_sc_hd__o21ai_2 _19098_ (.A1(_04263_),
    .A2(_04395_),
    .B1(_04228_),
    .Y(_04396_));
 sky130_fd_sc_hd__a32o_2 _19099_ (.A1(_04392_),
    .A2(_04316_),
    .A3(_04393_),
    .B1(_04394_),
    .B2(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__nand2_2 _19100_ (.A(_04396_),
    .B(_04310_),
    .Y(_04398_));
 sky130_fd_sc_hd__a31o_2 _19101_ (.A1(_03670_),
    .A2(_04229_),
    .A3(_04320_),
    .B1(_04396_),
    .X(_04399_));
 sky130_fd_sc_hd__nor4_2 _19102_ (.A(_03637_),
    .B(\decode.id_ex_aluop_reg[1] ),
    .C(\decode.id_ex_aluop_reg[3] ),
    .D(\decode.id_ex_aluop_reg[2] ),
    .Y(_04400_));
 sky130_fd_sc_hd__or4_2 _19103_ (.A(\decode.id_ex_aluop_reg[1] ),
    .B(\decode.id_ex_aluop_reg[3] ),
    .C(\decode.id_ex_aluop_reg[2] ),
    .D(_04299_),
    .X(_04401_));
 sky130_fd_sc_hd__a31o_2 _19104_ (.A1(_04006_),
    .A2(_04228_),
    .A3(_04231_),
    .B1(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__a31oi_2 _19105_ (.A1(_03983_),
    .A2(_04320_),
    .A3(_04396_),
    .B1(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__a31o_2 _19106_ (.A1(_04398_),
    .A2(_04399_),
    .A3(_04400_),
    .B1(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__or3_2 _19107_ (.A(_04390_),
    .B(_04397_),
    .C(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__o311a_2 _19108_ (.A1(_04346_),
    .A2(_04362_),
    .A3(_04370_),
    .B1(_04387_),
    .C1(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__and3_2 _19109_ (.A(_03594_),
    .B(_04361_),
    .C(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__buf_1 _19110_ (.A(_04407_),
    .X(_00549_));
 sky130_fd_sc_hd__buf_1 _19111_ (.A(_04225_),
    .X(_04408_));
 sky130_fd_sc_hd__buf_1 _19112_ (.A(_04243_),
    .X(_04409_));
 sky130_fd_sc_hd__o211a_2 _19113_ (.A1(_03863_),
    .A2(_04255_),
    .B1(_04338_),
    .C1(_04286_),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_2 _19114_ (.A0(_04275_),
    .A1(_04284_),
    .S(_04352_),
    .X(_04411_));
 sky130_fd_sc_hd__or3_2 _19115_ (.A(_04280_),
    .B(_04282_),
    .C(_04411_),
    .X(_04412_));
 sky130_fd_sc_hd__o21ai_2 _19116_ (.A1(_04273_),
    .A2(_04410_),
    .B1(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__nand2_2 _19117_ (.A(_04409_),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__buf_1 _19118_ (.A(_04242_),
    .X(_04415_));
 sky130_fd_sc_hd__o211a_2 _19119_ (.A1(_03956_),
    .A2(_04254_),
    .B1(_04265_),
    .C1(_04352_),
    .X(_04416_));
 sky130_fd_sc_hd__o21ba_2 _19120_ (.A1(_04248_),
    .A2(_04257_),
    .B1_N(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__a211o_2 _19121_ (.A1(_04297_),
    .A2(_04261_),
    .B1(_04263_),
    .C1(_04260_),
    .X(_04418_));
 sky130_fd_sc_hd__o221a_2 _19122_ (.A1(_04280_),
    .A2(_04282_),
    .B1(_04324_),
    .B2(_04276_),
    .C1(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__o21ba_2 _19123_ (.A1(_04269_),
    .A2(_04417_),
    .B1_N(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__and3_2 _19124_ (.A(_04412_),
    .B(_03704_),
    .C(_04332_),
    .X(_04421_));
 sky130_fd_sc_hd__o2bb2a_2 _19125_ (.A1_N(_04349_),
    .A2_N(_04420_),
    .B1(_04421_),
    .B2(_04414_),
    .X(_04422_));
 sky130_fd_sc_hd__o2111a_2 _19126_ (.A1(_04408_),
    .A2(_04414_),
    .B1(_04295_),
    .C1(_04415_),
    .D1(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__or3b_2 _19127_ (.A(\decode.id_ex_aluop_reg[1] ),
    .B(\decode.id_ex_aluop_reg[3] ),
    .C_N(\decode.id_ex_aluop_reg[2] ),
    .X(_04424_));
 sky130_fd_sc_hd__nor2_2 _19128_ (.A(_03638_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__o21ai_2 _19129_ (.A1(_04321_),
    .A2(_04234_),
    .B1(_04277_),
    .Y(_04426_));
 sky130_fd_sc_hd__o32a_2 _19130_ (.A1(_03983_),
    .A2(_04234_),
    .A3(_04277_),
    .B1(_04318_),
    .B2(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__buf_1 _19131_ (.A(_04392_),
    .X(_04428_));
 sky130_fd_sc_hd__and4b_2 _19132_ (.A_N(_04427_),
    .B(_04428_),
    .C(_04273_),
    .D(_04349_),
    .X(_04429_));
 sky130_fd_sc_hd__mux4_2 _19133_ (.A0(_04045_),
    .A1(_04054_),
    .A2(_03971_),
    .A3(_04321_),
    .S0(_04307_),
    .S1(_04325_),
    .X(_04430_));
 sky130_fd_sc_hd__mux2_2 _19134_ (.A0(_04250_),
    .A1(_04339_),
    .S(_04277_),
    .X(_04431_));
 sky130_fd_sc_hd__mux2_2 _19135_ (.A0(_04335_),
    .A1(_04340_),
    .S(_04247_),
    .X(_04432_));
 sky130_fd_sc_hd__mux2_2 _19136_ (.A0(_04431_),
    .A1(_04432_),
    .S(_04021_),
    .X(_04433_));
 sky130_fd_sc_hd__o211a_2 _19137_ (.A1(_04255_),
    .A2(_04070_),
    .B1(_04251_),
    .C1(_04252_),
    .X(_04434_));
 sky130_fd_sc_hd__a22o_2 _19138_ (.A1(_04249_),
    .A2(_04333_),
    .B1(_04434_),
    .B2(_04327_),
    .X(_04435_));
 sky130_fd_sc_hd__o21ai_2 _19139_ (.A1(_04280_),
    .A2(_04282_),
    .B1(_04289_),
    .Y(_04436_));
 sky130_fd_sc_hd__o2bb2a_2 _19140_ (.A1_N(_04244_),
    .A2_N(_04433_),
    .B1(_04435_),
    .B2(_04436_),
    .X(_04437_));
 sky130_fd_sc_hd__and4b_2 _19141_ (.A_N(_03635_),
    .B(_03634_),
    .C(_04056_),
    .D(_03633_),
    .X(_04438_));
 sky130_fd_sc_hd__buf_1 _19142_ (.A(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__o211a_2 _19143_ (.A1(_04305_),
    .A2(_04430_),
    .B1(_04437_),
    .C1(_04439_),
    .X(_04440_));
 sky130_fd_sc_hd__a311o_2 _19144_ (.A1(_04321_),
    .A2(_04425_),
    .A3(_04270_),
    .B1(_04429_),
    .C1(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__buf_1 _19145_ (.A(_04359_),
    .X(_04442_));
 sky130_fd_sc_hd__buf_1 _19146_ (.A(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__buf_1 _19147_ (.A(_04394_),
    .X(_04444_));
 sky130_fd_sc_hd__buf_1 _19148_ (.A(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__buf_1 _19149_ (.A(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__o21ai_2 _19150_ (.A1(_04443_),
    .A2(_04273_),
    .B1(_04446_),
    .Y(_04447_));
 sky130_fd_sc_hd__nand2_2 _19151_ (.A(_04321_),
    .B(_04021_),
    .Y(_04448_));
 sky130_fd_sc_hd__nand3_2 _19152_ (.A(_04006_),
    .B(_03983_),
    .C(_03988_),
    .Y(_04449_));
 sky130_fd_sc_hd__and4b_2 _19153_ (.A_N(_04022_),
    .B(_04448_),
    .C(_04228_),
    .D(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__a31o_2 _19154_ (.A1(_04006_),
    .A2(_03983_),
    .A3(_04320_),
    .B1(_04003_),
    .X(_04451_));
 sky130_fd_sc_hd__buf_1 _19155_ (.A(_04401_),
    .X(_04452_));
 sky130_fd_sc_hd__a21o_2 _19156_ (.A1(_04024_),
    .A2(_04451_),
    .B1(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__buf_1 _19157_ (.A(_04400_),
    .X(_04454_));
 sky130_fd_sc_hd__a22o_2 _19158_ (.A1(_04332_),
    .A2(_04373_),
    .B1(_04396_),
    .B2(_04310_),
    .X(_04455_));
 sky130_fd_sc_hd__xor2_2 _19159_ (.A(_04024_),
    .B(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__a2bb2o_2 _19160_ (.A1_N(_04450_),
    .A2_N(_04453_),
    .B1(_04454_),
    .B2(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__o22a_2 _19161_ (.A1(_04024_),
    .A2(_04447_),
    .B1(_04446_),
    .B2(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__buf_1 _19162_ (.A(_03594_),
    .X(_04459_));
 sky130_fd_sc_hd__o31a_2 _19163_ (.A1(_04423_),
    .A2(_04441_),
    .A3(_04458_),
    .B1(_04459_),
    .X(_00550_));
 sky130_fd_sc_hd__nor2_2 _19164_ (.A(_04321_),
    .B(_04274_),
    .Y(_04460_));
 sky130_fd_sc_hd__nor2_2 _19165_ (.A(_03971_),
    .B(_04254_),
    .Y(_04461_));
 sky130_fd_sc_hd__o211ai_2 _19166_ (.A1(_04373_),
    .A2(_04255_),
    .B1(_04231_),
    .C1(_04352_),
    .Y(_04462_));
 sky130_fd_sc_hd__o31a_2 _19167_ (.A1(_04248_),
    .A2(_04460_),
    .A3(_04461_),
    .B1(_04462_),
    .X(_04463_));
 sky130_fd_sc_hd__a2111o_2 _19168_ (.A1(_09974_),
    .A2(_03771_),
    .B1(_03970_),
    .C1(_03969_),
    .D1(_04289_),
    .X(_04464_));
 sky130_fd_sc_hd__buf_1 _19169_ (.A(_04308_),
    .X(_04465_));
 sky130_fd_sc_hd__o32a_2 _19170_ (.A1(_04303_),
    .A2(_04305_),
    .A3(_04463_),
    .B1(_04464_),
    .B2(_04465_),
    .X(_04466_));
 sky130_fd_sc_hd__o21ai_2 _19171_ (.A1(_04443_),
    .A2(_04362_),
    .B1(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__and3_2 _19172_ (.A(_03703_),
    .B(_04324_),
    .C(_04274_),
    .X(_04468_));
 sky130_fd_sc_hd__mux2_2 _19173_ (.A0(_04363_),
    .A1(_04367_),
    .S(_04246_),
    .X(_04469_));
 sky130_fd_sc_hd__or3b_2 _19174_ (.A(_04279_),
    .B(_04019_),
    .C_N(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__a21bo_2 _19175_ (.A1(_04269_),
    .A2(_04468_),
    .B1_N(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__mux2_2 _19176_ (.A0(_04364_),
    .A1(_04351_),
    .S(_04277_),
    .X(_04472_));
 sky130_fd_sc_hd__mux2_2 _19177_ (.A0(_04350_),
    .A1(_04354_),
    .S(_04264_),
    .X(_04473_));
 sky130_fd_sc_hd__mux2_2 _19178_ (.A0(_04472_),
    .A1(_04473_),
    .S(_04021_),
    .X(_04474_));
 sky130_fd_sc_hd__or2_2 _19179_ (.A(_04244_),
    .B(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__o21ai_2 _19180_ (.A1(_04349_),
    .A2(_04471_),
    .B1(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__nand2_2 _19181_ (.A(_04295_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__or2_2 _19182_ (.A(_04230_),
    .B(_04126_),
    .X(_04478_));
 sky130_fd_sc_hd__o211a_2 _19183_ (.A1(_04255_),
    .A2(_04062_),
    .B1(_04324_),
    .C1(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__o21ba_2 _19184_ (.A1(_04338_),
    .A2(_04377_),
    .B1_N(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__a21oi_2 _19185_ (.A1(_03997_),
    .A2(_03998_),
    .B1(_04379_),
    .Y(_04481_));
 sky130_fd_sc_hd__a31o_2 _19186_ (.A1(_04251_),
    .A2(_04252_),
    .A3(_04375_),
    .B1(_04481_),
    .X(_04482_));
 sky130_fd_sc_hd__and3_2 _19187_ (.A(_04381_),
    .B(_03998_),
    .C(_03997_),
    .X(_04483_));
 sky130_fd_sc_hd__a21oi_2 _19188_ (.A1(_04247_),
    .A2(_04355_),
    .B1(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__mux2_2 _19189_ (.A0(_04482_),
    .A1(_04484_),
    .S(_04268_),
    .X(_04485_));
 sky130_fd_sc_hd__nor2_2 _19190_ (.A(_04274_),
    .B(_04054_),
    .Y(_04486_));
 sky130_fd_sc_hd__a311o_2 _19191_ (.A1(_03986_),
    .A2(_03985_),
    .A3(_03984_),
    .B1(_03987_),
    .C1(_04070_),
    .X(_04487_));
 sky130_fd_sc_hd__o211ai_2 _19192_ (.A1(_04045_),
    .A2(_04320_),
    .B1(_04487_),
    .C1(_04332_),
    .Y(_04488_));
 sky130_fd_sc_hd__o311a_2 _19193_ (.A1(_04332_),
    .A2(_04486_),
    .A3(_04461_),
    .B1(_04317_),
    .C1(_04488_),
    .X(_04489_));
 sky130_fd_sc_hd__a221o_2 _19194_ (.A1(_04330_),
    .A2(_04480_),
    .B1(_04485_),
    .B2(_04409_),
    .C1(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__nand2_2 _19195_ (.A(_04490_),
    .B(_04346_),
    .Y(_04491_));
 sky130_fd_sc_hd__nor2_2 _19196_ (.A(_03637_),
    .B(_04306_),
    .Y(_04492_));
 sky130_fd_sc_hd__o21ai_2 _19197_ (.A1(_04022_),
    .A2(_04451_),
    .B1(_04448_),
    .Y(_04493_));
 sky130_fd_sc_hd__xnor2_2 _19198_ (.A(_04009_),
    .B(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__nor4_2 _19199_ (.A(_03633_),
    .B(\decode.id_ex_aluop_reg[3] ),
    .C(_03634_),
    .D(_04299_),
    .Y(_04495_));
 sky130_fd_sc_hd__buf_1 _19200_ (.A(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__o21a_2 _19201_ (.A1(_04279_),
    .A2(_04019_),
    .B1(_04321_),
    .X(_04497_));
 sky130_fd_sc_hd__a2bb2oi_2 _19202_ (.A1_N(_04022_),
    .A2_N(_04023_),
    .B1(_04389_),
    .B2(_04398_),
    .Y(_04498_));
 sky130_fd_sc_hd__or4_2 _19203_ (.A(_04008_),
    .B(_03976_),
    .C(_04497_),
    .D(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__o22ai_2 _19204_ (.A1(_04008_),
    .A2(_03976_),
    .B1(_04497_),
    .B2(_04498_),
    .Y(_04500_));
 sky130_fd_sc_hd__and3_2 _19205_ (.A(_04499_),
    .B(_04454_),
    .C(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__a211o_2 _19206_ (.A1(_04494_),
    .A2(_04496_),
    .B1(_04445_),
    .C1(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__buf_1 _19207_ (.A(_03638_),
    .X(_04503_));
 sky130_fd_sc_hd__buf_1 _19208_ (.A(_04311_),
    .X(_04504_));
 sky130_fd_sc_hd__buf_1 _19209_ (.A(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__a211o_2 _19210_ (.A1(_04245_),
    .A2(_04503_),
    .B1(_04505_),
    .C1(_04009_),
    .X(_04506_));
 sky130_fd_sc_hd__a32o_2 _19211_ (.A1(_04477_),
    .A2(_04491_),
    .A3(_04492_),
    .B1(_04502_),
    .B2(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__buf_1 _19212_ (.A(_04345_),
    .X(_04508_));
 sky130_fd_sc_hd__buf_1 _19213_ (.A(_04371_),
    .X(_04509_));
 sky130_fd_sc_hd__o21ai_2 _19214_ (.A1(_04281_),
    .A2(_04283_),
    .B1(_03704_),
    .Y(_04510_));
 sky130_fd_sc_hd__nand2_2 _19215_ (.A(_04470_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__o21a_2 _19216_ (.A1(_04509_),
    .A2(_04511_),
    .B1(_04475_),
    .X(_04512_));
 sky130_fd_sc_hd__o21a_2 _19217_ (.A1(_04508_),
    .A2(_04512_),
    .B1(_04491_),
    .X(_04513_));
 sky130_fd_sc_hd__nand2_2 _19218_ (.A(_03638_),
    .B(_04241_),
    .Y(_04514_));
 sky130_fd_sc_hd__buf_1 _19219_ (.A(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__o221a_2 _19220_ (.A1(_04467_),
    .A2(_04507_),
    .B1(_04513_),
    .B2(_04515_),
    .C1(_04459_),
    .X(_00551_));
 sky130_fd_sc_hd__and2_2 _19221_ (.A(_04038_),
    .B(_04054_),
    .X(_04516_));
 sky130_fd_sc_hd__o211ai_2 _19222_ (.A1(_04321_),
    .A2(_04021_),
    .B1(_04228_),
    .C1(_04449_),
    .Y(_04517_));
 sky130_fd_sc_hd__o211ai_2 _19223_ (.A1(_04027_),
    .A2(_04028_),
    .B1(_04448_),
    .C1(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__nand2_2 _19224_ (.A(_04027_),
    .B(_04028_),
    .Y(_04519_));
 sky130_fd_sc_hd__and3_2 _19225_ (.A(_04518_),
    .B(_04039_),
    .C(_04519_),
    .X(_04520_));
 sky130_fd_sc_hd__a21oi_2 _19226_ (.A1(_04519_),
    .A2(_04518_),
    .B1(_04039_),
    .Y(_04521_));
 sky130_fd_sc_hd__o211ai_2 _19227_ (.A1(_04054_),
    .A2(_04038_),
    .B1(_04394_),
    .C1(_03638_),
    .Y(_04522_));
 sky130_fd_sc_hd__o311a_2 _19228_ (.A1(_03638_),
    .A2(_04504_),
    .A3(_04039_),
    .B1(_04522_),
    .C1(_04308_),
    .X(_04523_));
 sky130_fd_sc_hd__o31a_2 _19229_ (.A1(_04520_),
    .A2(_04452_),
    .A3(_04521_),
    .B1(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__or4_2 _19230_ (.A(_03637_),
    .B(\decode.id_ex_aluop_reg[1] ),
    .C(\decode.id_ex_aluop_reg[3] ),
    .D(\decode.id_ex_aluop_reg[2] ),
    .X(_04525_));
 sky130_fd_sc_hd__buf_1 _19231_ (.A(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__or2_2 _19232_ (.A(_04034_),
    .B(_04055_),
    .X(_04527_));
 sky130_fd_sc_hd__nand2_2 _19233_ (.A(_04054_),
    .B(_04056_),
    .Y(_04528_));
 sky130_fd_sc_hd__a22oi_2 _19234_ (.A1(_04527_),
    .A2(_04528_),
    .B1(_04500_),
    .B2(_04464_),
    .Y(_04529_));
 sky130_fd_sc_hd__and3_2 _19235_ (.A(_04500_),
    .B(_04464_),
    .C(_04039_),
    .X(_04530_));
 sky130_fd_sc_hd__or3_2 _19236_ (.A(_04526_),
    .B(_04529_),
    .C(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__a2bb2o_2 _19237_ (.A1_N(_04516_),
    .A2_N(_04465_),
    .B1(_04524_),
    .B2(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__a211o_2 _19238_ (.A1(_04297_),
    .A2(_04261_),
    .B1(_04263_),
    .C1(_04284_),
    .X(_04533_));
 sky130_fd_sc_hd__nor2_2 _19239_ (.A(_04269_),
    .B(_04289_),
    .Y(_04534_));
 sky130_fd_sc_hd__mux2_2 _19240_ (.A0(_04278_),
    .A1(_04267_),
    .S(_04021_),
    .X(_04535_));
 sky130_fd_sc_hd__a32o_2 _19241_ (.A1(_04287_),
    .A2(_04533_),
    .A3(_04534_),
    .B1(_04535_),
    .B2(_04289_),
    .X(_04536_));
 sky130_fd_sc_hd__buf_1 _19242_ (.A(_04243_),
    .X(_04537_));
 sky130_fd_sc_hd__a31o_2 _19243_ (.A1(_03704_),
    .A2(_04537_),
    .A3(_04270_),
    .B1(_04536_),
    .X(_04538_));
 sky130_fd_sc_hd__and4b_2 _19244_ (.A_N(_03635_),
    .B(_03634_),
    .C(_03637_),
    .D(_03633_),
    .X(_04539_));
 sky130_fd_sc_hd__a22o_2 _19245_ (.A1(_04492_),
    .A2(_04536_),
    .B1(_04538_),
    .B2(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__buf_1 _19246_ (.A(_04272_),
    .X(_04541_));
 sky130_fd_sc_hd__mux2_2 _19247_ (.A0(_04259_),
    .A1(_04342_),
    .S(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__nand2_2 _19248_ (.A(_04542_),
    .B(_04409_),
    .Y(_04543_));
 sky130_fd_sc_hd__o221a_2 _19249_ (.A1(_04337_),
    .A2(_04436_),
    .B1(_04329_),
    .B2(_04305_),
    .C1(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__a2bb2o_2 _19250_ (.A1_N(_04439_),
    .A2_N(_04540_),
    .B1(_04544_),
    .B2(_04346_),
    .X(_04545_));
 sky130_fd_sc_hd__buf_1 _19251_ (.A(_04409_),
    .X(_04546_));
 sky130_fd_sc_hd__mux2_2 _19252_ (.A0(_04054_),
    .A1(_03971_),
    .S(_04233_),
    .X(_04547_));
 sky130_fd_sc_hd__a2bb2o_2 _19253_ (.A1_N(_04322_),
    .A2_N(_04318_),
    .B1(_04338_),
    .B2(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__a41o_2 _19254_ (.A1(_04325_),
    .A2(_04229_),
    .A3(_04307_),
    .A4(_03670_),
    .B1(_04541_),
    .X(_04549_));
 sky130_fd_sc_hd__o31a_2 _19255_ (.A1(_04281_),
    .A2(_04283_),
    .A3(_04548_),
    .B1(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__or4b_2 _19256_ (.A(_04295_),
    .B(_04546_),
    .C(_04301_),
    .D_N(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__a311oi_2 _19257_ (.A1(_04532_),
    .A2(_04545_),
    .A3(_04551_),
    .B1(_10576_),
    .C1(_10910_),
    .Y(_00552_));
 sky130_fd_sc_hd__and2b_2 _19258_ (.A_N(_04049_),
    .B(_04044_),
    .X(_04552_));
 sky130_fd_sc_hd__inv_2 _19259_ (.A(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__mux4_2 _19260_ (.A0(_04045_),
    .A1(_04054_),
    .A2(_03971_),
    .A3(_04321_),
    .S0(_04254_),
    .S1(_04352_),
    .X(_04554_));
 sky130_fd_sc_hd__or3_2 _19261_ (.A(_04280_),
    .B(_04282_),
    .C(_04554_),
    .X(_04555_));
 sky130_fd_sc_hd__o21ai_2 _19262_ (.A1(_04541_),
    .A2(_04393_),
    .B1(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__a21oi_2 _19263_ (.A1(_03638_),
    .A2(_04045_),
    .B1(_04504_),
    .Y(_04557_));
 sky130_fd_sc_hd__and2_2 _19264_ (.A(_04034_),
    .B(_04056_),
    .X(_04558_));
 sky130_fd_sc_hd__a31oi_2 _19265_ (.A1(_04518_),
    .A2(_04039_),
    .A3(_04519_),
    .B1(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__xor2_2 _19266_ (.A(_04052_),
    .B(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__o22a_2 _19267_ (.A1(_04050_),
    .A2(_04051_),
    .B1(_04516_),
    .B2(_04529_),
    .X(_04561_));
 sky130_fd_sc_hd__o41ai_2 _19268_ (.A1(_04050_),
    .A2(_04051_),
    .A3(_04516_),
    .A4(_04529_),
    .B1(_04400_),
    .Y(_04562_));
 sky130_fd_sc_hd__o22a_2 _19269_ (.A1(_04401_),
    .A2(_04560_),
    .B1(_04561_),
    .B2(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__a22o_2 _19270_ (.A1(_04052_),
    .A2(_04557_),
    .B1(_04563_),
    .B2(_04504_),
    .X(_04564_));
 sky130_fd_sc_hd__o311a_2 _19271_ (.A1(_04245_),
    .A2(_04303_),
    .A3(_04556_),
    .B1(_04564_),
    .C1(_04306_),
    .X(_04565_));
 sky130_fd_sc_hd__o21ai_2 _19272_ (.A1(_04465_),
    .A2(_04553_),
    .B1(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__mux2_2 _19273_ (.A0(_04356_),
    .A1(_04382_),
    .S(_04541_),
    .X(_04567_));
 sky130_fd_sc_hd__or3b_2 _19274_ (.A(_04243_),
    .B(_04541_),
    .C_N(_04378_),
    .X(_04568_));
 sky130_fd_sc_hd__o221a_2 _19275_ (.A1(_04305_),
    .A2(_04372_),
    .B1(_04567_),
    .B2(_04291_),
    .C1(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__mux2_2 _19276_ (.A0(_04365_),
    .A1(_04353_),
    .S(_04272_),
    .X(_04570_));
 sky130_fd_sc_hd__or2_2 _19277_ (.A(_04243_),
    .B(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__a21oi_2 _19278_ (.A1(_03863_),
    .A2(_04338_),
    .B1(_04307_),
    .Y(_04572_));
 sky130_fd_sc_hd__or3b_2 _19279_ (.A(_04280_),
    .B(_04282_),
    .C_N(_04368_),
    .X(_04573_));
 sky130_fd_sc_hd__o21ai_2 _19280_ (.A1(_04572_),
    .A2(_04573_),
    .B1(_04244_),
    .Y(_04574_));
 sky130_fd_sc_hd__a31o_2 _19281_ (.A1(_04294_),
    .A2(_04571_),
    .A3(_04574_),
    .B1(_04360_),
    .X(_04575_));
 sky130_fd_sc_hd__nand3_2 _19282_ (.A(_04244_),
    .B(_04510_),
    .C(_04573_),
    .Y(_04576_));
 sky130_fd_sc_hd__a31o_2 _19283_ (.A1(_04294_),
    .A2(_04571_),
    .A3(_04576_),
    .B1(_04514_),
    .X(_04577_));
 sky130_fd_sc_hd__a22o_2 _19284_ (.A1(_04346_),
    .A2(_04569_),
    .B1(_04575_),
    .B2(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__and3_2 _19285_ (.A(_03594_),
    .B(_04566_),
    .C(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__buf_1 _19286_ (.A(_04579_),
    .X(_00553_));
 sky130_fd_sc_hd__nand2_2 _19287_ (.A(_04075_),
    .B(_04172_),
    .Y(_04580_));
 sky130_fd_sc_hd__o21ai_2 _19288_ (.A1(_04443_),
    .A2(_04073_),
    .B1(_04446_),
    .Y(_04581_));
 sky130_fd_sc_hd__o21bai_2 _19289_ (.A1(_04050_),
    .A2(_04559_),
    .B1_N(_04051_),
    .Y(_04582_));
 sky130_fd_sc_hd__xor2_2 _19290_ (.A(_04226_),
    .B(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__o31a_2 _19291_ (.A1(_04552_),
    .A2(_04580_),
    .A3(_04561_),
    .B1(_04454_),
    .X(_04584_));
 sky130_fd_sc_hd__o22ai_2 _19292_ (.A1(_04050_),
    .A2(_04051_),
    .B1(_04516_),
    .B2(_04529_),
    .Y(_04585_));
 sky130_fd_sc_hd__a22o_2 _19293_ (.A1(_04075_),
    .A2(_04172_),
    .B1(_04585_),
    .B2(_04553_),
    .X(_04586_));
 sky130_fd_sc_hd__a221o_2 _19294_ (.A1(_04496_),
    .A2(_04583_),
    .B1(_04584_),
    .B2(_04586_),
    .C1(_04445_),
    .X(_04587_));
 sky130_fd_sc_hd__o21a_2 _19295_ (.A1(_04580_),
    .A2(_04581_),
    .B1(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__buf_1 _19296_ (.A(_04391_),
    .X(_04589_));
 sky130_fd_sc_hd__and2b_2 _19297_ (.A_N(_04073_),
    .B(_04070_),
    .X(_04590_));
 sky130_fd_sc_hd__mux2_2 _19298_ (.A0(_04045_),
    .A1(_04070_),
    .S(_04274_),
    .X(_04591_));
 sky130_fd_sc_hd__mux2_2 _19299_ (.A0(_04591_),
    .A1(_04547_),
    .S(_04247_),
    .X(_04592_));
 sky130_fd_sc_hd__o21ai_2 _19300_ (.A1(_04279_),
    .A2(_04019_),
    .B1(_04427_),
    .Y(_04593_));
 sky130_fd_sc_hd__o31a_2 _19301_ (.A1(_04280_),
    .A2(_04282_),
    .A3(_04592_),
    .B1(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__and4_2 _19302_ (.A(_03637_),
    .B(_04056_),
    .C(_04289_),
    .D(_04391_),
    .X(_04595_));
 sky130_fd_sc_hd__a32o_2 _19303_ (.A1(_04443_),
    .A2(_04589_),
    .A3(_04590_),
    .B1(_04594_),
    .B2(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__o211a_2 _19304_ (.A1(_04324_),
    .A2(_04276_),
    .B1(_04021_),
    .C1(_04418_),
    .X(_04597_));
 sky130_fd_sc_hd__a21o_2 _19305_ (.A1(_04269_),
    .A2(_04411_),
    .B1(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__o221a_2 _19306_ (.A1(_04270_),
    .A2(_04332_),
    .B1(_04244_),
    .B2(_04598_),
    .C1(_03705_),
    .X(_04599_));
 sky130_fd_sc_hd__a22o_2 _19307_ (.A1(_04410_),
    .A2(_04534_),
    .B1(_04598_),
    .B2(_04290_),
    .X(_04600_));
 sky130_fd_sc_hd__a211o_2 _19308_ (.A1(_04503_),
    .A2(_04599_),
    .B1(_04600_),
    .C1(_04346_),
    .X(_04601_));
 sky130_fd_sc_hd__mux2_2 _19309_ (.A0(_04417_),
    .A1(_04431_),
    .S(_04272_),
    .X(_04602_));
 sky130_fd_sc_hd__o22ai_2 _19310_ (.A1(_04436_),
    .A2(_04432_),
    .B1(_04371_),
    .B2(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__a211o_2 _19311_ (.A1(_04435_),
    .A2(_04317_),
    .B1(_04294_),
    .C1(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__and3_2 _19312_ (.A(_04601_),
    .B(_04604_),
    .C(_04415_),
    .X(_04605_));
 sky130_fd_sc_hd__o31a_2 _19313_ (.A1(_04588_),
    .A2(_04596_),
    .A3(_04605_),
    .B1(_04459_),
    .X(_00554_));
 sky130_fd_sc_hd__o21ai_2 _19314_ (.A1(_04279_),
    .A2(_04019_),
    .B1(_04473_),
    .Y(_04606_));
 sky130_fd_sc_hd__o31a_2 _19315_ (.A1(_04280_),
    .A2(_04019_),
    .A3(_04484_),
    .B1(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__a22o_2 _19316_ (.A1(_04330_),
    .A2(_04482_),
    .B1(_04607_),
    .B2(_04243_),
    .X(_04608_));
 sky130_fd_sc_hd__a31o_2 _19317_ (.A1(_04290_),
    .A2(_04273_),
    .A3(_04480_),
    .B1(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__nand2_2 _19318_ (.A(_04609_),
    .B(_04345_),
    .Y(_04610_));
 sky130_fd_sc_hd__a22oi_2 _19319_ (.A1(_04075_),
    .A2(_04172_),
    .B1(_04585_),
    .B2(_04553_),
    .Y(_04611_));
 sky130_fd_sc_hd__o22ai_2 _19320_ (.A1(_04171_),
    .A2(_04173_),
    .B1(_04611_),
    .B2(_04590_),
    .Y(_04612_));
 sky130_fd_sc_hd__or4_2 _19321_ (.A(_04171_),
    .B(_04173_),
    .C(_04611_),
    .D(_04590_),
    .X(_04613_));
 sky130_fd_sc_hd__a21bo_2 _19322_ (.A1(_04582_),
    .A2(_04075_),
    .B1_N(_04172_),
    .X(_04614_));
 sky130_fd_sc_hd__xnor2_2 _19323_ (.A(_04227_),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__o21ai_2 _19324_ (.A1(_04452_),
    .A2(_04615_),
    .B1(_04505_),
    .Y(_04616_));
 sky130_fd_sc_hd__a31oi_2 _19325_ (.A1(_04454_),
    .A2(_04612_),
    .A3(_04613_),
    .B1(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__buf_1 _19326_ (.A(_04442_),
    .X(_04618_));
 sky130_fd_sc_hd__o211a_2 _19327_ (.A1(_04065_),
    .A2(_04618_),
    .B1(_04445_),
    .C1(_04227_),
    .X(_04619_));
 sky130_fd_sc_hd__buf_1 _19328_ (.A(_04424_),
    .X(_04620_));
 sky130_fd_sc_hd__or2b_2 _19329_ (.A(_04065_),
    .B_N(_04062_),
    .X(_04621_));
 sky130_fd_sc_hd__or3_2 _19330_ (.A(_04408_),
    .B(_04620_),
    .C(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__o21ai_2 _19331_ (.A1(_04045_),
    .A2(_04234_),
    .B1(_04247_),
    .Y(_04623_));
 sky130_fd_sc_hd__o21ai_2 _19332_ (.A1(_04234_),
    .A2(_04062_),
    .B1(_04487_),
    .Y(_04624_));
 sky130_fd_sc_hd__o221a_2 _19333_ (.A1(_04623_),
    .A2(_04486_),
    .B1(_04249_),
    .B2(_04624_),
    .C1(_04541_),
    .X(_04625_));
 sky130_fd_sc_hd__a21o_2 _19334_ (.A1(_04270_),
    .A2(_04463_),
    .B1(_04625_),
    .X(_04626_));
 sky130_fd_sc_hd__mux2_2 _19335_ (.A0(_04469_),
    .A1(_04472_),
    .S(_04021_),
    .X(_04627_));
 sky130_fd_sc_hd__o211a_2 _19336_ (.A1(_03972_),
    .A2(_03974_),
    .B1(_04007_),
    .C1(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__a31o_2 _19337_ (.A1(_04244_),
    .A2(_04273_),
    .A3(_04468_),
    .B1(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__o2111ai_2 _19338_ (.A1(_04345_),
    .A2(_04629_),
    .B1(_04242_),
    .C1(_04442_),
    .D1(_04610_),
    .Y(_04630_));
 sky130_fd_sc_hd__o311a_2 _19339_ (.A1(_04546_),
    .A2(_04303_),
    .A3(_04626_),
    .B1(_04630_),
    .C1(_04515_),
    .X(_04631_));
 sky130_fd_sc_hd__o211ai_2 _19340_ (.A1(_04617_),
    .A2(_04619_),
    .B1(_04622_),
    .C1(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__a21o_2 _19341_ (.A1(_03704_),
    .A2(_04537_),
    .B1(_04345_),
    .X(_04633_));
 sky130_fd_sc_hd__or4_2 _19342_ (.A(_04443_),
    .B(_04362_),
    .C(_04633_),
    .D(_04628_),
    .X(_04634_));
 sky130_fd_sc_hd__o2111a_2 _19343_ (.A1(_04515_),
    .A2(_04610_),
    .B1(_04632_),
    .C1(_04634_),
    .D1(_03595_),
    .X(_00555_));
 sky130_fd_sc_hd__or2_2 _19344_ (.A(_04130_),
    .B(_04131_),
    .X(_04635_));
 sky130_fd_sc_hd__o21ai_2 _19345_ (.A1(_04618_),
    .A2(_04129_),
    .B1(_04446_),
    .Y(_04636_));
 sky130_fd_sc_hd__a41oi_2 _19346_ (.A1(_04582_),
    .A2(_04172_),
    .A3(_04075_),
    .A4(_04227_),
    .B1(_04174_),
    .Y(_04637_));
 sky130_fd_sc_hd__a21oi_2 _19347_ (.A1(_04637_),
    .A2(_04635_),
    .B1(_04452_),
    .Y(_04638_));
 sky130_fd_sc_hd__or3_2 _19348_ (.A(_04130_),
    .B(_04131_),
    .C(_04637_),
    .X(_04639_));
 sky130_fd_sc_hd__nand2_2 _19349_ (.A(_04612_),
    .B(_04621_),
    .Y(_04640_));
 sky130_fd_sc_hd__o31a_2 _19350_ (.A1(_04130_),
    .A2(_04131_),
    .A3(_04640_),
    .B1(_04454_),
    .X(_04641_));
 sky130_fd_sc_hd__a2bb2o_2 _19351_ (.A1_N(_04130_),
    .A2_N(_04131_),
    .B1(_04612_),
    .B2(_04621_),
    .X(_04642_));
 sky130_fd_sc_hd__a22o_2 _19352_ (.A1(_04638_),
    .A2(_04639_),
    .B1(_04641_),
    .B2(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__o22a_2 _19353_ (.A1(_04635_),
    .A2(_04636_),
    .B1(_04446_),
    .B2(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__nand2b_2 _19354_ (.A_N(_04129_),
    .B(_04126_),
    .Y(_04645_));
 sky130_fd_sc_hd__a311o_2 _19355_ (.A1(_04017_),
    .A2(_04015_),
    .A3(_04016_),
    .B1(_04282_),
    .C1(_04289_),
    .X(_04646_));
 sky130_fd_sc_hd__o21a_2 _19356_ (.A1(_04254_),
    .A2(_04126_),
    .B1(_04327_),
    .X(_04647_));
 sky130_fd_sc_hd__mux2_2 _19357_ (.A0(_04647_),
    .A1(_04591_),
    .S(_04248_),
    .X(_04648_));
 sky130_fd_sc_hd__mux2_2 _19358_ (.A0(_04648_),
    .A1(_04548_),
    .S(_04270_),
    .X(_04649_));
 sky130_fd_sc_hd__a2bb2o_2 _19359_ (.A1_N(_04296_),
    .A2_N(_04646_),
    .B1(_04649_),
    .B2(_04349_),
    .X(_04650_));
 sky130_fd_sc_hd__a2bb2o_2 _19360_ (.A1_N(_04465_),
    .A2_N(_04645_),
    .B1(_04428_),
    .B2(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__a311o_2 _19361_ (.A1(_04245_),
    .A2(_03705_),
    .A3(_04503_),
    .B1(_04345_),
    .C1(_04362_),
    .X(_04652_));
 sky130_fd_sc_hd__a21oi_2 _19362_ (.A1(_04273_),
    .A2(_04278_),
    .B1(_04288_),
    .Y(_04653_));
 sky130_fd_sc_hd__nor2_2 _19363_ (.A(_04546_),
    .B(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__o21ai_2 _19364_ (.A1(_04270_),
    .A2(_04337_),
    .B1(_04343_),
    .Y(_04655_));
 sky130_fd_sc_hd__o211a_2 _19365_ (.A1(_03972_),
    .A2(_03974_),
    .B1(_04007_),
    .C1(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__a211o_2 _19366_ (.A1(_04271_),
    .A2(_04546_),
    .B1(_04295_),
    .C1(_04362_),
    .X(_04657_));
 sky130_fd_sc_hd__o22a_2 _19367_ (.A1(_04652_),
    .A2(_04654_),
    .B1(_04656_),
    .B2(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__o311a_2 _19368_ (.A1(_04415_),
    .A2(_04644_),
    .A3(_04651_),
    .B1(_04658_),
    .C1(_03595_),
    .X(_00556_));
 sky130_fd_sc_hd__a211o_2 _19369_ (.A1(_04612_),
    .A2(_04621_),
    .B1(_04132_),
    .C1(_04144_),
    .X(_04659_));
 sky130_fd_sc_hd__o211ai_2 _19370_ (.A1(_04144_),
    .A2(_04645_),
    .B1(_04454_),
    .C1(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__a31oi_2 _19371_ (.A1(_04144_),
    .A2(_04642_),
    .A3(_04645_),
    .B1(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__o21ai_2 _19372_ (.A1(_04142_),
    .A2(_04143_),
    .B1(_04639_),
    .Y(_04662_));
 sky130_fd_sc_hd__or4_2 _19373_ (.A(_04635_),
    .B(_04142_),
    .C(_04143_),
    .D(_04637_),
    .X(_04663_));
 sky130_fd_sc_hd__nand2_2 _19374_ (.A(_04126_),
    .B(_04129_),
    .Y(_04664_));
 sky130_fd_sc_hd__o31a_2 _19375_ (.A1(_04143_),
    .A2(_04664_),
    .A3(_04142_),
    .B1(_04496_),
    .X(_04665_));
 sky130_fd_sc_hd__o211a_2 _19376_ (.A1(_04131_),
    .A2(_04662_),
    .B1(_04663_),
    .C1(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__buf_1 _19377_ (.A(_04311_),
    .X(_04667_));
 sky130_fd_sc_hd__a2111o_2 _19378_ (.A1(_04503_),
    .A2(_04137_),
    .B1(_04667_),
    .C1(_04143_),
    .D1(_04142_),
    .X(_04668_));
 sky130_fd_sc_hd__o31a_2 _19379_ (.A1(_04446_),
    .A2(_04661_),
    .A3(_04666_),
    .B1(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__or2_2 _19380_ (.A(_04376_),
    .B(_04141_),
    .X(_04670_));
 sky130_fd_sc_hd__o21a_2 _19381_ (.A1(_04253_),
    .A2(_04137_),
    .B1(_04478_),
    .X(_04671_));
 sky130_fd_sc_hd__o211a_2 _19382_ (.A1(_04254_),
    .A2(_04062_),
    .B1(_04487_),
    .C1(_04352_),
    .X(_04672_));
 sky130_fd_sc_hd__a31o_2 _19383_ (.A1(_04251_),
    .A2(_04252_),
    .A3(_04671_),
    .B1(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__mux2_2 _19384_ (.A0(_04673_),
    .A1(_04554_),
    .S(_04269_),
    .X(_04674_));
 sky130_fd_sc_hd__a22o_2 _19385_ (.A1(_04393_),
    .A2(_04534_),
    .B1(_04674_),
    .B2(_04371_),
    .X(_04675_));
 sky130_fd_sc_hd__a2bb2o_2 _19386_ (.A1_N(_04465_),
    .A2_N(_04670_),
    .B1(_04428_),
    .B2(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__mux2_2 _19387_ (.A0(_04357_),
    .A1(_04384_),
    .S(_04349_),
    .X(_04677_));
 sky130_fd_sc_hd__a211o_2 _19388_ (.A1(_04509_),
    .A2(_04369_),
    .B1(_04515_),
    .C1(_04633_),
    .X(_04678_));
 sky130_fd_sc_hd__and3_2 _19389_ (.A(_04291_),
    .B(_04369_),
    .C(_04358_),
    .X(_04679_));
 sky130_fd_sc_hd__or4_2 _19390_ (.A(_03639_),
    .B(_04345_),
    .C(_04306_),
    .D(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__o211a_2 _19391_ (.A1(_04386_),
    .A2(_04677_),
    .B1(_04678_),
    .C1(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__o311a_2 _19392_ (.A1(_04415_),
    .A2(_04669_),
    .A3(_04676_),
    .B1(_04681_),
    .C1(_03595_),
    .X(_00557_));
 sky130_fd_sc_hd__o21a_2 _19393_ (.A1(_04359_),
    .A2(_04160_),
    .B1(_04444_),
    .X(_04682_));
 sky130_fd_sc_hd__o21a_2 _19394_ (.A1(_04664_),
    .A2(_04142_),
    .B1(_04177_),
    .X(_04683_));
 sky130_fd_sc_hd__a22oi_2 _19395_ (.A1(_04165_),
    .A2(_04167_),
    .B1(_04663_),
    .B2(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__a41o_2 _19396_ (.A1(_04683_),
    .A2(_04663_),
    .A3(_04167_),
    .A4(_04165_),
    .B1(_04401_),
    .X(_04685_));
 sky130_fd_sc_hd__o211ai_2 _19397_ (.A1(_04645_),
    .A2(_04144_),
    .B1(_04670_),
    .C1(_04659_),
    .Y(_04686_));
 sky130_fd_sc_hd__xor2_2 _19398_ (.A(_04168_),
    .B(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__o22a_2 _19399_ (.A1(_04684_),
    .A2(_04685_),
    .B1(_04526_),
    .B2(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__a22o_2 _19400_ (.A1(_04168_),
    .A2(_04682_),
    .B1(_04688_),
    .B2(_04505_),
    .X(_04689_));
 sky130_fd_sc_hd__mux2_2 _19401_ (.A0(_04166_),
    .A1(_04137_),
    .S(_04234_),
    .X(_04690_));
 sky130_fd_sc_hd__mux2_2 _19402_ (.A0(_04647_),
    .A1(_04690_),
    .S(_04324_),
    .X(_04691_));
 sky130_fd_sc_hd__mux2_2 _19403_ (.A0(_04691_),
    .A1(_04592_),
    .S(_04269_),
    .X(_04692_));
 sky130_fd_sc_hd__o2bb2a_2 _19404_ (.A1_N(_04291_),
    .A2_N(_04692_),
    .B1(_04646_),
    .B2(_04427_),
    .X(_04693_));
 sky130_fd_sc_hd__o32a_2 _19405_ (.A1(_03639_),
    .A2(_04165_),
    .A3(_04620_),
    .B1(_04303_),
    .B2(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__or2_2 _19406_ (.A(_04243_),
    .B(_04433_),
    .X(_04695_));
 sky130_fd_sc_hd__o211a_2 _19407_ (.A1(_04291_),
    .A2(_04420_),
    .B1(_04695_),
    .C1(_04345_),
    .X(_04696_));
 sky130_fd_sc_hd__o21a_2 _19408_ (.A1(_04409_),
    .A2(_04413_),
    .B1(_04038_),
    .X(_04697_));
 sky130_fd_sc_hd__o31a_2 _19409_ (.A1(_04503_),
    .A2(_04696_),
    .A3(_04697_),
    .B1(_04242_),
    .X(_04698_));
 sky130_fd_sc_hd__a31o_2 _19410_ (.A1(_04360_),
    .A2(_04689_),
    .A3(_04694_),
    .B1(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__o211a_2 _19411_ (.A1(_04273_),
    .A2(_04410_),
    .B1(_04290_),
    .C1(_04412_),
    .X(_04700_));
 sky130_fd_sc_hd__a211o_2 _19412_ (.A1(_04371_),
    .A2(_04421_),
    .B1(_04633_),
    .C1(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__or4b_2 _19413_ (.A(_04443_),
    .B(_04362_),
    .C(_04696_),
    .D_N(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__a21oi_2 _19414_ (.A1(_04699_),
    .A2(_04702_),
    .B1(_03587_),
    .Y(_00558_));
 sky130_fd_sc_hd__nor2_2 _19415_ (.A(_04334_),
    .B(_04152_),
    .Y(_04703_));
 sky130_fd_sc_hd__mux2_2 _19416_ (.A0(_04149_),
    .A1(_04166_),
    .S(_03989_),
    .X(_04704_));
 sky130_fd_sc_hd__mux2_2 _19417_ (.A0(_04671_),
    .A1(_04704_),
    .S(_04277_),
    .X(_04705_));
 sky130_fd_sc_hd__o221a_2 _19418_ (.A1(_04623_),
    .A2(_04486_),
    .B1(_04247_),
    .B2(_04624_),
    .C1(_04268_),
    .X(_04706_));
 sky130_fd_sc_hd__o21ba_2 _19419_ (.A1(_04268_),
    .A2(_04705_),
    .B1_N(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__a2bb2o_2 _19420_ (.A1_N(_04646_),
    .A2_N(_04463_),
    .B1(_04289_),
    .B2(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__a32o_2 _19421_ (.A1(_04359_),
    .A2(_04703_),
    .A3(_04391_),
    .B1(_04708_),
    .B2(_04392_),
    .X(_04709_));
 sky130_fd_sc_hd__a21o_2 _19422_ (.A1(_04471_),
    .A2(_04289_),
    .B1(_04056_),
    .X(_04710_));
 sky130_fd_sc_hd__nor2_2 _19423_ (.A(_04028_),
    .B(_04485_),
    .Y(_04711_));
 sky130_fd_sc_hd__a211o_2 _19424_ (.A1(_04474_),
    .A2(_04243_),
    .B1(_04038_),
    .C1(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__and3_2 _19425_ (.A(_04710_),
    .B(_04241_),
    .C(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__o21a_2 _19426_ (.A1(_04359_),
    .A2(_04152_),
    .B1(_04394_),
    .X(_04714_));
 sky130_fd_sc_hd__inv_2 _19427_ (.A(_04155_),
    .Y(_04715_));
 sky130_fd_sc_hd__a21oi_2 _19428_ (.A1(_04166_),
    .A2(_04164_),
    .B1(_04684_),
    .Y(_04716_));
 sky130_fd_sc_hd__or2_2 _19429_ (.A(_04715_),
    .B(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__a221o_2 _19430_ (.A1(_04153_),
    .A2(_04154_),
    .B1(_04166_),
    .B2(_04164_),
    .C1(_04684_),
    .X(_04718_));
 sky130_fd_sc_hd__o22a_2 _19431_ (.A1(_04130_),
    .A2(_04131_),
    .B1(_04142_),
    .B2(_04143_),
    .X(_04719_));
 sky130_fd_sc_hd__o221ai_2 _19432_ (.A1(_04376_),
    .A2(_04141_),
    .B1(_04645_),
    .B2(_04144_),
    .C1(_04165_),
    .Y(_04720_));
 sky130_fd_sc_hd__a21oi_2 _19433_ (.A1(_04640_),
    .A2(_04719_),
    .B1(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__a21oi_2 _19434_ (.A1(_04160_),
    .A2(_04164_),
    .B1(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__a211o_2 _19435_ (.A1(_04160_),
    .A2(_04164_),
    .B1(_04155_),
    .C1(_04721_),
    .X(_04723_));
 sky130_fd_sc_hd__o211a_2 _19436_ (.A1(_04715_),
    .A2(_04722_),
    .B1(_04400_),
    .C1(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__a31o_2 _19437_ (.A1(_04495_),
    .A2(_04717_),
    .A3(_04718_),
    .B1(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__o2bb2a_2 _19438_ (.A1_N(_04155_),
    .A2_N(_04714_),
    .B1(_04444_),
    .B2(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__or4_2 _19439_ (.A(_04539_),
    .B(_04709_),
    .C(_04713_),
    .D(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__and3b_2 _19440_ (.A_N(_10909_),
    .B(_03636_),
    .C(_09954_),
    .X(_04728_));
 sky130_fd_sc_hd__buf_1 _19441_ (.A(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__a211o_2 _19442_ (.A1(_04511_),
    .A2(_04509_),
    .B1(_04515_),
    .C1(_04633_),
    .X(_04730_));
 sky130_fd_sc_hd__or3_2 _19443_ (.A(_04618_),
    .B(_04306_),
    .C(_04712_),
    .X(_04731_));
 sky130_fd_sc_hd__and4_2 _19444_ (.A(_04727_),
    .B(_04729_),
    .C(_04730_),
    .D(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__buf_1 _19445_ (.A(_04732_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_2 _19446_ (.A0(_04112_),
    .A1(_04149_),
    .S(_04234_),
    .X(_04733_));
 sky130_fd_sc_hd__mux2_2 _19447_ (.A0(_04733_),
    .A1(_04690_),
    .S(_04248_),
    .X(_04734_));
 sky130_fd_sc_hd__mux2_2 _19448_ (.A0(_04648_),
    .A1(_04734_),
    .S(_04541_),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_2 _19449_ (.A0(_04735_),
    .A1(_04550_),
    .S(_04409_),
    .X(_04736_));
 sky130_fd_sc_hd__and4_2 _19450_ (.A(_04736_),
    .B(_04589_),
    .C(_04346_),
    .D(_04408_),
    .X(_04737_));
 sky130_fd_sc_hd__o21ai_2 _19451_ (.A1(_04664_),
    .A2(_04142_),
    .B1(_04177_),
    .Y(_04738_));
 sky130_fd_sc_hd__a22o_2 _19452_ (.A1(_04149_),
    .A2(_04152_),
    .B1(_04166_),
    .B2(_04164_),
    .X(_04739_));
 sky130_fd_sc_hd__a32o_2 _19453_ (.A1(_04155_),
    .A2(_04168_),
    .A3(_04738_),
    .B1(_04739_),
    .B2(_04154_),
    .X(_04740_));
 sky130_fd_sc_hd__o21bai_2 _19454_ (.A1(_04169_),
    .A2(_04637_),
    .B1_N(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__and2_2 _19455_ (.A(_04741_),
    .B(_04120_),
    .X(_04742_));
 sky130_fd_sc_hd__nor2_2 _19456_ (.A(_04120_),
    .B(_04741_),
    .Y(_04743_));
 sky130_fd_sc_hd__a22o_2 _19457_ (.A1(_04334_),
    .A2(_04152_),
    .B1(_04160_),
    .B2(_04164_),
    .X(_04744_));
 sky130_fd_sc_hd__o22ai_2 _19458_ (.A1(_04334_),
    .A2(_04152_),
    .B1(_04744_),
    .B2(_04721_),
    .Y(_04745_));
 sky130_fd_sc_hd__xor2_2 _19459_ (.A(_04120_),
    .B(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__o32a_2 _19460_ (.A1(_04452_),
    .A2(_04742_),
    .A3(_04743_),
    .B1(_04526_),
    .B2(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__o211a_2 _19461_ (.A1(_04115_),
    .A2(_04442_),
    .B1(_04444_),
    .C1(_04120_),
    .X(_04748_));
 sky130_fd_sc_hd__a21oi_2 _19462_ (.A1(_04747_),
    .A2(_04505_),
    .B1(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__a31o_2 _19463_ (.A1(_04112_),
    .A2(_04118_),
    .A3(_04425_),
    .B1(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__o211a_2 _19464_ (.A1(_04332_),
    .A2(_04284_),
    .B1(_04317_),
    .C1(_04287_),
    .X(_04751_));
 sky130_fd_sc_hd__a31o_2 _19465_ (.A1(_04408_),
    .A2(_03705_),
    .A3(_04305_),
    .B1(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__or2_2 _19466_ (.A(_04291_),
    .B(_04535_),
    .X(_04753_));
 sky130_fd_sc_hd__o211a_2 _19467_ (.A1(_04245_),
    .A2(_04542_),
    .B1(_04346_),
    .C1(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__a211o_2 _19468_ (.A1(_04295_),
    .A2(_04752_),
    .B1(_04362_),
    .C1(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__o311a_2 _19469_ (.A1(_04415_),
    .A2(_04737_),
    .A3(_04750_),
    .B1(_04755_),
    .C1(_04729_),
    .X(_00560_));
 sky130_fd_sc_hd__inv_2 _19470_ (.A(_04120_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand2_2 _19471_ (.A(_04745_),
    .B(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__nand2_2 _19472_ (.A(_04118_),
    .B(_04112_),
    .Y(_04758_));
 sky130_fd_sc_hd__a41o_2 _19473_ (.A1(_04104_),
    .A2(_04112_),
    .A3(_04118_),
    .A4(_04106_),
    .B1(_04525_),
    .X(_04759_));
 sky130_fd_sc_hd__a31o_2 _19474_ (.A1(_04107_),
    .A2(_04757_),
    .A3(_04758_),
    .B1(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__o21bai_2 _19475_ (.A1(_04107_),
    .A2(_04757_),
    .B1_N(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__or3_2 _19476_ (.A(_04119_),
    .B(_04107_),
    .C(_04742_),
    .X(_04762_));
 sky130_fd_sc_hd__o21ai_2 _19477_ (.A1(_04119_),
    .A2(_04742_),
    .B1(_04107_),
    .Y(_04763_));
 sky130_fd_sc_hd__nand3_2 _19478_ (.A(_04762_),
    .B(_04763_),
    .C(_04496_),
    .Y(_04764_));
 sky130_fd_sc_hd__a211o_2 _19479_ (.A1(_04103_),
    .A2(_04100_),
    .B1(_04359_),
    .C1(_04504_),
    .X(_04765_));
 sky130_fd_sc_hd__o311a_2 _19480_ (.A1(_04504_),
    .A2(_04225_),
    .A3(_04107_),
    .B1(_04465_),
    .C1(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__a32o_2 _19481_ (.A1(_04761_),
    .A2(_04764_),
    .A3(_04766_),
    .B1(_04104_),
    .B2(_04425_),
    .X(_04767_));
 sky130_fd_sc_hd__mux2_2 _19482_ (.A0(_04112_),
    .A1(_04105_),
    .S(_04274_),
    .X(_04768_));
 sky130_fd_sc_hd__mux2_2 _19483_ (.A0(_04768_),
    .A1(_04704_),
    .S(_04352_),
    .X(_04769_));
 sky130_fd_sc_hd__mux2_2 _19484_ (.A0(_04673_),
    .A1(_04769_),
    .S(_04541_),
    .X(_04770_));
 sky130_fd_sc_hd__nand2_2 _19485_ (.A(_04409_),
    .B(_04556_),
    .Y(_04771_));
 sky130_fd_sc_hd__o21ai_2 _19486_ (.A1(_04409_),
    .A2(_04770_),
    .B1(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__or4_2 _19487_ (.A(_04618_),
    .B(_04294_),
    .C(_04620_),
    .D(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__mux2_2 _19488_ (.A0(_04570_),
    .A1(_04567_),
    .S(_04371_),
    .X(_04774_));
 sky130_fd_sc_hd__o2bb2a_2 _19489_ (.A1_N(_04304_),
    .A2_N(_03704_),
    .B1(_04537_),
    .B2(_04573_),
    .X(_04775_));
 sky130_fd_sc_hd__or3_2 _19490_ (.A(_04537_),
    .B(_04572_),
    .C(_04573_),
    .X(_04776_));
 sky130_fd_sc_hd__a22o_2 _19491_ (.A1(_04539_),
    .A2(_04775_),
    .B1(_04776_),
    .B2(_04492_),
    .X(_04777_));
 sky130_fd_sc_hd__a2bb2o_2 _19492_ (.A1_N(_04386_),
    .A2_N(_04774_),
    .B1(_04777_),
    .B2(_04295_),
    .X(_04778_));
 sky130_fd_sc_hd__or4b_2 _19493_ (.A(reset),
    .B(_10908_),
    .C(_10758_),
    .D_N(_03636_),
    .X(_04779_));
 sky130_fd_sc_hd__a311oi_2 _19494_ (.A1(_04362_),
    .A2(_04767_),
    .A3(_04773_),
    .B1(_04778_),
    .C1(_04779_),
    .Y(_00561_));
 sky130_fd_sc_hd__a211o_2 _19495_ (.A1(_04085_),
    .A2(_04225_),
    .B1(_04504_),
    .C1(_04186_),
    .X(_04780_));
 sky130_fd_sc_hd__o32a_2 _19496_ (.A1(_04117_),
    .A2(_04115_),
    .A3(_04107_),
    .B1(_04103_),
    .B2(_04100_),
    .X(_04781_));
 sky130_fd_sc_hd__o21ai_2 _19497_ (.A1(_04107_),
    .A2(_04757_),
    .B1(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__nand2_2 _19498_ (.A(_04186_),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__or2_2 _19499_ (.A(_04186_),
    .B(_04782_),
    .X(_04784_));
 sky130_fd_sc_hd__a221o_2 _19500_ (.A1(_03708_),
    .A2(\decode.id_ex_imm_reg[13] ),
    .B1(_04101_),
    .B2(_04102_),
    .C1(_04100_),
    .X(_04785_));
 sky130_fd_sc_hd__a21o_2 _19501_ (.A1(_04785_),
    .A2(_04763_),
    .B1(_04186_),
    .X(_04786_));
 sky130_fd_sc_hd__nand3_2 _19502_ (.A(_04186_),
    .B(_04785_),
    .C(_04763_),
    .Y(_04787_));
 sky130_fd_sc_hd__a31o_2 _19503_ (.A1(_04786_),
    .A2(_04787_),
    .A3(_04495_),
    .B1(_04444_),
    .X(_04788_));
 sky130_fd_sc_hd__a31o_2 _19504_ (.A1(_04454_),
    .A2(_04783_),
    .A3(_04784_),
    .B1(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__mux2_2 _19505_ (.A0(_04181_),
    .A1(_04105_),
    .S(_04253_),
    .X(_04790_));
 sky130_fd_sc_hd__mux2_2 _19506_ (.A0(_04733_),
    .A1(_04790_),
    .S(_04324_),
    .X(_04791_));
 sky130_fd_sc_hd__mux2_2 _19507_ (.A0(_04691_),
    .A1(_04791_),
    .S(_04272_),
    .X(_04792_));
 sky130_fd_sc_hd__or2_2 _19508_ (.A(_04289_),
    .B(_04594_),
    .X(_04793_));
 sky130_fd_sc_hd__o21ai_2 _19509_ (.A1(_04537_),
    .A2(_04792_),
    .B1(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__a21oi_2 _19510_ (.A1(_04083_),
    .A2(_04084_),
    .B1(_04081_),
    .Y(_04795_));
 sky130_fd_sc_hd__a2bb2o_2 _19511_ (.A1_N(_04302_),
    .A2_N(_04794_),
    .B1(_04795_),
    .B2(_04425_),
    .X(_04796_));
 sky130_fd_sc_hd__a211o_2 _19512_ (.A1(_04780_),
    .A2(_04789_),
    .B1(_04796_),
    .C1(_04242_),
    .X(_04797_));
 sky130_fd_sc_hd__o211a_2 _19513_ (.A1(_04270_),
    .A2(_04332_),
    .B1(_03704_),
    .C1(_04291_),
    .X(_04798_));
 sky130_fd_sc_hd__and3_2 _19514_ (.A(_04290_),
    .B(_04273_),
    .C(_04410_),
    .X(_04799_));
 sky130_fd_sc_hd__or4_2 _19515_ (.A(_04514_),
    .B(_04798_),
    .C(_04633_),
    .D(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__nand2_2 _19516_ (.A(_04602_),
    .B(_04291_),
    .Y(_04801_));
 sky130_fd_sc_hd__o211a_2 _19517_ (.A1(_04291_),
    .A2(_04598_),
    .B1(_04345_),
    .C1(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__a221o_2 _19518_ (.A1(_04386_),
    .A2(_04360_),
    .B1(_04799_),
    .B2(_04294_),
    .C1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__and4_2 _19519_ (.A(_04729_),
    .B(_04797_),
    .C(_04800_),
    .D(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__buf_1 _19520_ (.A(_04804_),
    .X(_00562_));
 sky130_fd_sc_hd__buf_1 _19521_ (.A(_04346_),
    .X(_04805_));
 sky130_fd_sc_hd__or3_2 _19522_ (.A(_04359_),
    .B(_04306_),
    .C(_03704_),
    .X(_04806_));
 sky130_fd_sc_hd__and3_2 _19523_ (.A(_04349_),
    .B(_04273_),
    .C(_04468_),
    .X(_04807_));
 sky130_fd_sc_hd__nor2_2 _19524_ (.A(_04245_),
    .B(_04607_),
    .Y(_04808_));
 sky130_fd_sc_hd__a211o_2 _19525_ (.A1(_04245_),
    .A2(_04627_),
    .B1(_04294_),
    .C1(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__o311a_2 _19526_ (.A1(_04408_),
    .A2(_04508_),
    .A3(_04807_),
    .B1(_04415_),
    .C1(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__or2_2 _19527_ (.A(_04091_),
    .B(_04094_),
    .X(_04811_));
 sky130_fd_sc_hd__mux2_2 _19528_ (.A0(_04180_),
    .A1(_04181_),
    .S(_03989_),
    .X(_04812_));
 sky130_fd_sc_hd__a21o_2 _19529_ (.A1(_04251_),
    .A2(_04252_),
    .B1(_04768_),
    .X(_04813_));
 sky130_fd_sc_hd__o21ai_2 _19530_ (.A1(_04249_),
    .A2(_04812_),
    .B1(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__o21ai_2 _19531_ (.A1(_04281_),
    .A2(_04283_),
    .B1(_04705_),
    .Y(_04815_));
 sky130_fd_sc_hd__o31a_2 _19532_ (.A1(_04281_),
    .A2(_04283_),
    .A3(_04814_),
    .B1(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__mux2_2 _19533_ (.A0(_04626_),
    .A1(_04816_),
    .S(_04349_),
    .X(_04817_));
 sky130_fd_sc_hd__a21oi_2 _19534_ (.A1(_04186_),
    .A2(_04782_),
    .B1(_04795_),
    .Y(_04818_));
 sky130_fd_sc_hd__o21ai_2 _19535_ (.A1(_04081_),
    .A2(_04085_),
    .B1(_04786_),
    .Y(_04819_));
 sky130_fd_sc_hd__a221oi_2 _19536_ (.A1(_04454_),
    .A2(_04818_),
    .B1(_04819_),
    .B2(_04496_),
    .C1(_04445_),
    .Y(_04820_));
 sky130_fd_sc_hd__a21oi_2 _19537_ (.A1(_03638_),
    .A2(_04444_),
    .B1(_04095_),
    .Y(_04821_));
 sky130_fd_sc_hd__o221a_2 _19538_ (.A1(_04818_),
    .A2(_04526_),
    .B1(_04452_),
    .B2(_04819_),
    .C1(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__and4_2 _19539_ (.A(_04225_),
    .B(_04094_),
    .C(_04444_),
    .D(_04091_),
    .X(_04823_));
 sky130_fd_sc_hd__a211o_2 _19540_ (.A1(_04095_),
    .A2(_04820_),
    .B1(_04822_),
    .C1(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__o221ai_2 _19541_ (.A1(_04811_),
    .A2(_04465_),
    .B1(_04817_),
    .B2(_04303_),
    .C1(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__o221a_2 _19542_ (.A1(_04805_),
    .A2(_04806_),
    .B1(_04810_),
    .B2(_04825_),
    .C1(_04729_),
    .X(_00563_));
 sky130_fd_sc_hd__nand2_2 _19543_ (.A(_04408_),
    .B(_03929_),
    .Y(_04826_));
 sky130_fd_sc_hd__nand2_2 _19544_ (.A(_04095_),
    .B(_04186_),
    .Y(_04827_));
 sky130_fd_sc_hd__and4b_2 _19545_ (.A_N(_04827_),
    .B(_04106_),
    .C(_04104_),
    .D(_04756_),
    .X(_04828_));
 sky130_fd_sc_hd__nand2_2 _19546_ (.A(_04745_),
    .B(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__a221o_2 _19547_ (.A1(_04083_),
    .A2(_04084_),
    .B1(_04094_),
    .B2(_04091_),
    .C1(_04081_),
    .X(_04830_));
 sky130_fd_sc_hd__o211a_2 _19548_ (.A1(_04827_),
    .A2(_04781_),
    .B1(_04811_),
    .C1(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__a21oi_2 _19549_ (.A1(_04829_),
    .A2(_04831_),
    .B1(_04211_),
    .Y(_04832_));
 sky130_fd_sc_hd__a31o_2 _19550_ (.A1(_04829_),
    .A2(_04831_),
    .A3(_04211_),
    .B1(_04526_),
    .X(_04833_));
 sky130_fd_sc_hd__nor2_2 _19551_ (.A(_04186_),
    .B(_04095_),
    .Y(_04834_));
 sky130_fd_sc_hd__nand4_2 _19552_ (.A(_04740_),
    .B(_04120_),
    .C(_04834_),
    .D(_04107_),
    .Y(_04835_));
 sky130_fd_sc_hd__o21ai_2 _19553_ (.A1(_04105_),
    .A2(_04103_),
    .B1(_04119_),
    .Y(_04836_));
 sky130_fd_sc_hd__a211oi_2 _19554_ (.A1(_04785_),
    .A2(_04836_),
    .B1(_04186_),
    .C1(_04095_),
    .Y(_04837_));
 sky130_fd_sc_hd__o211a_2 _19555_ (.A1(_04180_),
    .A2(_04094_),
    .B1(_04181_),
    .C1(_04182_),
    .X(_04838_));
 sky130_fd_sc_hd__a211oi_2 _19556_ (.A1(_04180_),
    .A2(_04094_),
    .B1(_04837_),
    .C1(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__o211ai_2 _19557_ (.A1(_04637_),
    .A2(_04170_),
    .B1(_04835_),
    .C1(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hd__a21oi_2 _19558_ (.A1(_04840_),
    .A2(_04211_),
    .B1(_04452_),
    .Y(_04841_));
 sky130_fd_sc_hd__o21ai_2 _19559_ (.A1(_04211_),
    .A2(_04840_),
    .B1(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__o211a_2 _19560_ (.A1(_04832_),
    .A2(_04833_),
    .B1(_04842_),
    .C1(_04505_),
    .X(_04843_));
 sky130_fd_sc_hd__a31o_2 _19561_ (.A1(_04211_),
    .A2(_04446_),
    .A3(_04826_),
    .B1(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__or4_2 _19562_ (.A(_04408_),
    .B(_04209_),
    .C(_04620_),
    .D(_03933_),
    .X(_04845_));
 sky130_fd_sc_hd__or4b_2 _19563_ (.A(_04038_),
    .B(_04371_),
    .C(_04301_),
    .D_N(_04649_),
    .X(_04846_));
 sky130_fd_sc_hd__mux2_2 _19564_ (.A0(_03929_),
    .A1(_04180_),
    .S(_04253_),
    .X(_04847_));
 sky130_fd_sc_hd__and3_2 _19565_ (.A(_04847_),
    .B(_04252_),
    .C(_04251_),
    .X(_04848_));
 sky130_fd_sc_hd__a21oi_2 _19566_ (.A1(_04332_),
    .A2(_04790_),
    .B1(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__o21ai_2 _19567_ (.A1(_04281_),
    .A2(_04283_),
    .B1(_04734_),
    .Y(_04850_));
 sky130_fd_sc_hd__o31a_2 _19568_ (.A1(_04281_),
    .A2(_04283_),
    .A3(_04849_),
    .B1(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__or4_2 _19569_ (.A(_04056_),
    .B(_04296_),
    .C(_04301_),
    .D(_04305_),
    .X(_04852_));
 sky130_fd_sc_hd__o311a_2 _19570_ (.A1(_04409_),
    .A2(_04302_),
    .A3(_04851_),
    .B1(_04852_),
    .C1(_04515_),
    .X(_04853_));
 sky130_fd_sc_hd__o311a_2 _19571_ (.A1(_04408_),
    .A2(_04293_),
    .A3(_04386_),
    .B1(_04846_),
    .C1(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__o311a_2 _19572_ (.A1(_04442_),
    .A2(_03705_),
    .A3(_04306_),
    .B1(_03636_),
    .C1(_03593_),
    .X(_04855_));
 sky130_fd_sc_hd__o21ai_2 _19573_ (.A1(_04618_),
    .A2(_04386_),
    .B1(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__o31a_2 _19574_ (.A1(_04295_),
    .A2(_04293_),
    .A3(_04779_),
    .B1(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__a31oi_2 _19575_ (.A1(_04844_),
    .A2(_04845_),
    .A3(_04854_),
    .B1(_04857_),
    .Y(_00564_));
 sky130_fd_sc_hd__a21o_2 _19576_ (.A1(_04198_),
    .A2(_04359_),
    .B1(_04504_),
    .X(_04858_));
 sky130_fd_sc_hd__o22a_2 _19577_ (.A1(_03639_),
    .A2(_04620_),
    .B1(_04197_),
    .B2(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__nor2_2 _19578_ (.A(_04197_),
    .B(_04198_),
    .Y(_04860_));
 sky130_fd_sc_hd__inv_2 _19579_ (.A(_04211_),
    .Y(_04861_));
 sky130_fd_sc_hd__or3b_2 _19580_ (.A(_04861_),
    .B(_04860_),
    .C_N(_04840_),
    .X(_04862_));
 sky130_fd_sc_hd__o211ai_2 _19581_ (.A1(_04197_),
    .A2(_04198_),
    .B1(_03929_),
    .C1(_03933_),
    .Y(_04863_));
 sky130_fd_sc_hd__nor2_2 _19582_ (.A(_04209_),
    .B(_03933_),
    .Y(_04864_));
 sky130_fd_sc_hd__or3_2 _19583_ (.A(_04209_),
    .B(_03933_),
    .C(_04197_),
    .X(_04865_));
 sky130_fd_sc_hd__a21boi_2 _19584_ (.A1(_04745_),
    .A2(_04828_),
    .B1_N(_04831_),
    .Y(_04866_));
 sky130_fd_sc_hd__or4_2 _19585_ (.A(_04211_),
    .B(_04197_),
    .C(_04198_),
    .D(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__o211a_2 _19586_ (.A1(_04198_),
    .A2(_04865_),
    .B1(_04400_),
    .C1(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__o31a_2 _19587_ (.A1(_04860_),
    .A2(_04832_),
    .A3(_04864_),
    .B1(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__a31oi_2 _19588_ (.A1(_04496_),
    .A2(_04862_),
    .A3(_04863_),
    .B1(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__a31o_2 _19589_ (.A1(_04210_),
    .A2(_04860_),
    .A3(_04841_),
    .B1(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__o2bb2a_2 _19590_ (.A1_N(_04859_),
    .A2_N(_04871_),
    .B1(_04465_),
    .B2(_04198_),
    .X(_04872_));
 sky130_fd_sc_hd__o21a_2 _19591_ (.A1(_04349_),
    .A2(_04358_),
    .B1(_04370_),
    .X(_04873_));
 sky130_fd_sc_hd__and3_2 _19592_ (.A(_04873_),
    .B(_04492_),
    .C(_04508_),
    .X(_04874_));
 sky130_fd_sc_hd__o21a_2 _19593_ (.A1(_03934_),
    .A2(_04253_),
    .B1(_04380_),
    .X(_04875_));
 sky130_fd_sc_hd__mux2_2 _19594_ (.A0(_04812_),
    .A1(_04875_),
    .S(_04277_),
    .X(_04876_));
 sky130_fd_sc_hd__mux2_2 _19595_ (.A0(_04769_),
    .A1(_04876_),
    .S(_04272_),
    .X(_04877_));
 sky130_fd_sc_hd__and3_2 _19596_ (.A(_04038_),
    .B(_04391_),
    .C(_03637_),
    .X(_04878_));
 sky130_fd_sc_hd__buf_1 _19597_ (.A(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__a31o_2 _19598_ (.A1(_04317_),
    .A2(_04393_),
    .A3(_04879_),
    .B1(_04539_),
    .X(_04880_));
 sky130_fd_sc_hd__a31o_2 _19599_ (.A1(_04674_),
    .A2(_04546_),
    .A3(_04428_),
    .B1(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__a31o_2 _19600_ (.A1(_04509_),
    .A2(_04428_),
    .A3(_04877_),
    .B1(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__o311a_2 _19601_ (.A1(_04442_),
    .A2(_04294_),
    .A3(_04362_),
    .B1(_04806_),
    .C1(_04728_),
    .X(_04883_));
 sky130_fd_sc_hd__a31o_2 _19602_ (.A1(_04805_),
    .A2(_04370_),
    .A3(_04729_),
    .B1(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__o31a_2 _19603_ (.A1(_04872_),
    .A2(_04874_),
    .A3(_04882_),
    .B1(_04884_),
    .X(_00565_));
 sky130_fd_sc_hd__o21a_2 _19604_ (.A1(_03911_),
    .A2(_03935_),
    .B1(_04865_),
    .X(_04885_));
 sky130_fd_sc_hd__a31o_2 _19605_ (.A1(_04867_),
    .A2(_04885_),
    .A3(_04202_),
    .B1(_04526_),
    .X(_04886_));
 sky130_fd_sc_hd__o2bb2a_2 _19606_ (.A1_N(_04885_),
    .A2_N(_04867_),
    .B1(_03938_),
    .B2(_04201_),
    .X(_04887_));
 sky130_fd_sc_hd__o2111a_2 _19607_ (.A1(_04201_),
    .A2(_03938_),
    .B1(_04862_),
    .C1(_04863_),
    .D1(_03912_),
    .X(_04888_));
 sky130_fd_sc_hd__a311o_2 _19608_ (.A1(_03912_),
    .A2(_04862_),
    .A3(_04863_),
    .B1(_04201_),
    .C1(_03938_),
    .X(_04889_));
 sky130_fd_sc_hd__or3b_2 _19609_ (.A(_04888_),
    .B(_04452_),
    .C_N(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__o211a_2 _19610_ (.A1(_04886_),
    .A2(_04887_),
    .B1(_04505_),
    .C1(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__o211a_2 _19611_ (.A1(_03923_),
    .A2(_04443_),
    .B1(_04446_),
    .C1(_04202_),
    .X(_04892_));
 sky130_fd_sc_hd__nor2_2 _19612_ (.A(_04891_),
    .B(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hd__o211a_2 _19613_ (.A1(_03972_),
    .A2(_03974_),
    .B1(_04007_),
    .C1(_04420_),
    .X(_04894_));
 sky130_fd_sc_hd__and4b_2 _19614_ (.A_N(_04894_),
    .B(_04414_),
    .C(_04508_),
    .D(_04242_),
    .X(_04895_));
 sky130_fd_sc_hd__mux2_2 _19615_ (.A0(_03918_),
    .A1(_03934_),
    .S(_04253_),
    .X(_04896_));
 sky130_fd_sc_hd__mux2_2 _19616_ (.A0(_04847_),
    .A1(_04896_),
    .S(_04277_),
    .X(_04897_));
 sky130_fd_sc_hd__mux2_2 _19617_ (.A0(_04791_),
    .A1(_04897_),
    .S(_04272_),
    .X(_04898_));
 sky130_fd_sc_hd__nor2_2 _19618_ (.A(_04199_),
    .B(_03923_),
    .Y(_04899_));
 sky130_fd_sc_hd__and4b_2 _19619_ (.A_N(_04427_),
    .B(_04879_),
    .C(_04290_),
    .D(_04541_),
    .X(_04900_));
 sky130_fd_sc_hd__a221o_2 _19620_ (.A1(_04225_),
    .A2(_04242_),
    .B1(_04425_),
    .B2(_04899_),
    .C1(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__a31o_2 _19621_ (.A1(_04509_),
    .A2(_04428_),
    .A3(_04898_),
    .B1(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__a31o_2 _19622_ (.A1(_04546_),
    .A2(_04428_),
    .A3(_04692_),
    .B1(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__a31o_2 _19623_ (.A1(_04805_),
    .A2(_04422_),
    .A3(_04729_),
    .B1(_04883_),
    .X(_04904_));
 sky130_fd_sc_hd__o31a_2 _19624_ (.A1(_04893_),
    .A2(_04895_),
    .A3(_04903_),
    .B1(_04904_),
    .X(_00566_));
 sky130_fd_sc_hd__and3_2 _19625_ (.A(_03594_),
    .B(_04345_),
    .C(_03636_),
    .X(_04905_));
 sky130_fd_sc_hd__a21oi_2 _19626_ (.A1(_04512_),
    .A2(_04905_),
    .B1(_04883_),
    .Y(_04906_));
 sky130_fd_sc_hd__and4_2 _19627_ (.A(_04503_),
    .B(_04203_),
    .C(_04445_),
    .D(_03902_),
    .X(_04907_));
 sky130_fd_sc_hd__a21oi_2 _19628_ (.A1(_04204_),
    .A2(_04206_),
    .B1(_03638_),
    .Y(_04908_));
 sky130_fd_sc_hd__o22ai_2 _19629_ (.A1(_03638_),
    .A2(_04207_),
    .B1(_04887_),
    .B2(_04899_),
    .Y(_04909_));
 sky130_fd_sc_hd__o31ai_2 _19630_ (.A1(_04887_),
    .A2(_04899_),
    .A3(_04908_),
    .B1(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__and2_2 _19631_ (.A(_04204_),
    .B(_04206_),
    .X(_04911_));
 sky130_fd_sc_hd__and3_2 _19632_ (.A(_03912_),
    .B(_04862_),
    .C(_04863_),
    .X(_04912_));
 sky130_fd_sc_hd__o21ai_2 _19633_ (.A1(_03938_),
    .A2(_04912_),
    .B1(_03924_),
    .Y(_04913_));
 sky130_fd_sc_hd__and3_2 _19634_ (.A(_03924_),
    .B(_04889_),
    .C(_04207_),
    .X(_04914_));
 sky130_fd_sc_hd__a211oi_2 _19635_ (.A1(_04911_),
    .A2(_04913_),
    .B1(_04401_),
    .C1(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__nor4_2 _19636_ (.A(_03633_),
    .B(_03635_),
    .C(_03634_),
    .D(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__o2bb2a_2 _19637_ (.A1_N(_04910_),
    .A2_N(_04916_),
    .B1(_04908_),
    .B2(_04667_),
    .X(_04917_));
 sky130_fd_sc_hd__mux2_2 _19638_ (.A0(_04205_),
    .A1(_03918_),
    .S(_04253_),
    .X(_04918_));
 sky130_fd_sc_hd__mux2_2 _19639_ (.A0(_04918_),
    .A1(_04875_),
    .S(_04247_),
    .X(_04919_));
 sky130_fd_sc_hd__or3b_2 _19640_ (.A(_04280_),
    .B(_04282_),
    .C_N(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__o21a_2 _19641_ (.A1(_04541_),
    .A2(_04814_),
    .B1(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__o32a_2 _19642_ (.A1(_04244_),
    .A2(_04302_),
    .A3(_04921_),
    .B1(_04308_),
    .B2(_04206_),
    .X(_04922_));
 sky130_fd_sc_hd__or4b_2 _19643_ (.A(_04038_),
    .B(_04290_),
    .C(_04301_),
    .D_N(_04707_),
    .X(_04923_));
 sky130_fd_sc_hd__or3_2 _19644_ (.A(_04299_),
    .B(_04424_),
    .C(_04056_),
    .X(_04924_));
 sky130_fd_sc_hd__or4_2 _19645_ (.A(_04537_),
    .B(_04270_),
    .C(_04924_),
    .D(_04463_),
    .X(_04925_));
 sky130_fd_sc_hd__and4_2 _19646_ (.A(_04922_),
    .B(_04923_),
    .C(_04925_),
    .D(_04515_),
    .X(_04926_));
 sky130_fd_sc_hd__o221a_2 _19647_ (.A1(_04386_),
    .A2(_04476_),
    .B1(_04907_),
    .B2(_04917_),
    .C1(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__nor2_2 _19648_ (.A(_04906_),
    .B(_04927_),
    .Y(_00567_));
 sky130_fd_sc_hd__o2111ai_2 _19649_ (.A1(_04201_),
    .A2(_03938_),
    .B1(_04911_),
    .C1(_04860_),
    .D1(_04861_),
    .Y(_04928_));
 sky130_fd_sc_hd__a21oi_2 _19650_ (.A1(_04829_),
    .A2(_04831_),
    .B1(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__o31ai_2 _19651_ (.A1(_04202_),
    .A2(_04207_),
    .A3(_04885_),
    .B1(_04206_),
    .Y(_04930_));
 sky130_fd_sc_hd__a31o_2 _19652_ (.A1(_03918_),
    .A2(_04200_),
    .A3(_04204_),
    .B1(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__o21bai_2 _19653_ (.A1(_04866_),
    .A2(_04928_),
    .B1_N(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__a21oi_2 _19654_ (.A1(_04932_),
    .A2(_04192_),
    .B1(_04526_),
    .Y(_04933_));
 sky130_fd_sc_hd__o31a_2 _19655_ (.A1(_04192_),
    .A2(_04929_),
    .A3(_04931_),
    .B1(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__a211o_2 _19656_ (.A1(_04204_),
    .A2(_04206_),
    .B1(_04201_),
    .C1(_03938_),
    .X(_04935_));
 sky130_fd_sc_hd__o31a_2 _19657_ (.A1(_04199_),
    .A2(_04200_),
    .A3(_03937_),
    .B1(_03903_),
    .X(_04936_));
 sky130_fd_sc_hd__o21ai_2 _19658_ (.A1(_04935_),
    .A2(_04912_),
    .B1(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__nand3b_2 _19659_ (.A_N(_03957_),
    .B(_03960_),
    .C(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__o211ai_2 _19660_ (.A1(_04935_),
    .A2(_04912_),
    .B1(_04936_),
    .C1(_04192_),
    .Y(_04939_));
 sky130_fd_sc_hd__and3_2 _19661_ (.A(_04938_),
    .B(_04939_),
    .C(_04496_),
    .X(_04940_));
 sky130_fd_sc_hd__a211o_2 _19662_ (.A1(_03959_),
    .A2(_03639_),
    .B1(_04667_),
    .C1(_04192_),
    .X(_04941_));
 sky130_fd_sc_hd__o31a_2 _19663_ (.A1(_04446_),
    .A2(_04934_),
    .A3(_04940_),
    .B1(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__and3_2 _19664_ (.A(_03959_),
    .B(_04425_),
    .C(_03956_),
    .X(_04943_));
 sky130_fd_sc_hd__o21a_2 _19665_ (.A1(_03956_),
    .A2(_04234_),
    .B1(_04256_),
    .X(_04944_));
 sky130_fd_sc_hd__mux2_2 _19666_ (.A0(_04944_),
    .A1(_04896_),
    .S(_04248_),
    .X(_04945_));
 sky130_fd_sc_hd__a211o_2 _19667_ (.A1(_04790_),
    .A2(_04249_),
    .B1(_04272_),
    .C1(_04848_),
    .X(_04946_));
 sky130_fd_sc_hd__o31a_2 _19668_ (.A1(_04281_),
    .A2(_04283_),
    .A3(_04945_),
    .B1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__a32o_2 _19669_ (.A1(_04509_),
    .A2(_04550_),
    .A3(_04879_),
    .B1(_04947_),
    .B2(_04595_),
    .X(_04948_));
 sky130_fd_sc_hd__buf_1 _19670_ (.A(_04539_),
    .X(_04949_));
 sky130_fd_sc_hd__a31o_2 _19671_ (.A1(_04735_),
    .A2(_04245_),
    .A3(_04428_),
    .B1(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__a31o_2 _19672_ (.A1(_04508_),
    .A2(_04492_),
    .A3(_04536_),
    .B1(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__a31o_2 _19673_ (.A1(_04805_),
    .A2(_04538_),
    .A3(_04728_),
    .B1(_04883_),
    .X(_04952_));
 sky130_fd_sc_hd__o41a_2 _19674_ (.A1(_04942_),
    .A2(_04943_),
    .A3(_04948_),
    .A4(_04951_),
    .B1(_04952_),
    .X(_00568_));
 sky130_fd_sc_hd__a31oi_2 _19675_ (.A1(_04574_),
    .A2(_04439_),
    .A3(_04571_),
    .B1(_04949_),
    .Y(_04953_));
 sky130_fd_sc_hd__a21o_2 _19676_ (.A1(_03947_),
    .A2(_03944_),
    .B1(_04503_),
    .X(_04954_));
 sky130_fd_sc_hd__a21o_2 _19677_ (.A1(_03960_),
    .A2(_04938_),
    .B1(_04191_),
    .X(_04955_));
 sky130_fd_sc_hd__nand3_2 _19678_ (.A(_04191_),
    .B(_03960_),
    .C(_04938_),
    .Y(_04956_));
 sky130_fd_sc_hd__and3_2 _19679_ (.A(_04932_),
    .B(_04192_),
    .C(_04191_),
    .X(_04957_));
 sky130_fd_sc_hd__a221oi_2 _19680_ (.A1(_03956_),
    .A2(_03959_),
    .B1(_04932_),
    .B2(_04192_),
    .C1(_04191_),
    .Y(_04958_));
 sky130_fd_sc_hd__a311o_2 _19681_ (.A1(_04191_),
    .A2(_03956_),
    .A3(_03959_),
    .B1(_04525_),
    .C1(_04958_),
    .X(_04959_));
 sky130_fd_sc_hd__nor2_2 _19682_ (.A(_04957_),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__a311o_2 _19683_ (.A1(_04496_),
    .A2(_04955_),
    .A3(_04956_),
    .B1(_04960_),
    .C1(_04445_),
    .X(_04961_));
 sky130_fd_sc_hd__a211o_2 _19684_ (.A1(_03947_),
    .A2(_03639_),
    .B1(_04667_),
    .C1(_04191_),
    .X(_04962_));
 sky130_fd_sc_hd__a22o_2 _19685_ (.A1(_04589_),
    .A2(_04954_),
    .B1(_04961_),
    .B2(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__mux2_2 _19686_ (.A0(_03944_),
    .A1(_03956_),
    .S(_04253_),
    .X(_04964_));
 sky130_fd_sc_hd__mux2_2 _19687_ (.A0(_04964_),
    .A1(_04918_),
    .S(_04247_),
    .X(_04965_));
 sky130_fd_sc_hd__mux2_2 _19688_ (.A0(_04965_),
    .A1(_04876_),
    .S(_04268_),
    .X(_04966_));
 sky130_fd_sc_hd__o21ai_2 _19689_ (.A1(_04546_),
    .A2(_04556_),
    .B1(_04879_),
    .Y(_04967_));
 sky130_fd_sc_hd__or4_2 _19690_ (.A(_04294_),
    .B(_04371_),
    .C(_04301_),
    .D(_04770_),
    .X(_04968_));
 sky130_fd_sc_hd__o311a_2 _19691_ (.A1(_04546_),
    .A2(_04966_),
    .A3(_04303_),
    .B1(_04967_),
    .C1(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__nand2_2 _19692_ (.A(_04963_),
    .B(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__and3_2 _19693_ (.A(_04905_),
    .B(_04576_),
    .C(_04571_),
    .X(_04971_));
 sky130_fd_sc_hd__o2bb2a_2 _19694_ (.A1_N(_04953_),
    .A2_N(_04970_),
    .B1(_04971_),
    .B2(_04883_),
    .X(_00569_));
 sky130_fd_sc_hd__a32o_2 _19695_ (.A1(_04191_),
    .A2(_03956_),
    .A3(_03959_),
    .B1(_03947_),
    .B2(_03944_),
    .X(_04972_));
 sky130_fd_sc_hd__o22a_2 _19696_ (.A1(_04189_),
    .A2(_03894_),
    .B1(_04972_),
    .B2(_04957_),
    .X(_04973_));
 sky130_fd_sc_hd__or2_2 _19697_ (.A(_04189_),
    .B(_03894_),
    .X(_04974_));
 sky130_fd_sc_hd__o31ai_2 _19698_ (.A1(_04974_),
    .A2(_04972_),
    .A3(_04957_),
    .B1(_04454_),
    .Y(_04975_));
 sky130_fd_sc_hd__nor2_2 _19699_ (.A(_04973_),
    .B(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__a21oi_2 _19700_ (.A1(_04937_),
    .A2(_04193_),
    .B1(_03963_),
    .Y(_04977_));
 sky130_fd_sc_hd__a21oi_2 _19701_ (.A1(_04977_),
    .A2(_04974_),
    .B1(_04452_),
    .Y(_04978_));
 sky130_fd_sc_hd__o31a_2 _19702_ (.A1(_04189_),
    .A2(_03894_),
    .A3(_04977_),
    .B1(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__a2111o_2 _19703_ (.A1(_04503_),
    .A2(_03888_),
    .B1(_04189_),
    .C1(_04505_),
    .D1(_03894_),
    .X(_04980_));
 sky130_fd_sc_hd__o31a_2 _19704_ (.A1(_04446_),
    .A2(_04976_),
    .A3(_04979_),
    .B1(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__and2b_2 _19705_ (.A_N(_03893_),
    .B(_03888_),
    .X(_04982_));
 sky130_fd_sc_hd__o211a_2 _19706_ (.A1(_03888_),
    .A2(_04234_),
    .B1(_04277_),
    .C1(_04265_),
    .X(_04983_));
 sky130_fd_sc_hd__a21o_2 _19707_ (.A1(_04944_),
    .A2(_04352_),
    .B1(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__mux2_2 _19708_ (.A0(_04984_),
    .A1(_04897_),
    .S(_04268_),
    .X(_04985_));
 sky130_fd_sc_hd__a32o_2 _19709_ (.A1(_04290_),
    .A2(_04594_),
    .A3(_04879_),
    .B1(_04985_),
    .B2(_04595_),
    .X(_04986_));
 sky130_fd_sc_hd__a31o_2 _19710_ (.A1(_04600_),
    .A2(_04359_),
    .A3(_04439_),
    .B1(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__a311o_2 _19711_ (.A1(_04618_),
    .A2(_04391_),
    .A3(_04982_),
    .B1(_04949_),
    .C1(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__a31o_2 _19712_ (.A1(_04546_),
    .A2(_04428_),
    .A3(_04792_),
    .B1(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__o211a_2 _19713_ (.A1(_04599_),
    .A2(_04600_),
    .B1(_04728_),
    .C1(_04805_),
    .X(_04990_));
 sky130_fd_sc_hd__o22a_2 _19714_ (.A1(_04981_),
    .A2(_04989_),
    .B1(_04883_),
    .B2(_04990_),
    .X(_00570_));
 sky130_fd_sc_hd__o221ai_2 _19715_ (.A1(_03868_),
    .A2(_03701_),
    .B1(_03689_),
    .B2(\decode.id_ex_rs1_data_reg[23] ),
    .C1(_03871_),
    .Y(_04991_));
 sky130_fd_sc_hd__or2_2 _19716_ (.A(_04991_),
    .B(_03881_),
    .X(_04992_));
 sky130_fd_sc_hd__nand2_2 _19717_ (.A(_03881_),
    .B(_04991_),
    .Y(_04993_));
 sky130_fd_sc_hd__or2_2 _19718_ (.A(_04973_),
    .B(_04982_),
    .X(_04994_));
 sky130_fd_sc_hd__or2_2 _19719_ (.A(_04194_),
    .B(_03882_),
    .X(_04995_));
 sky130_fd_sc_hd__o21ai_2 _19720_ (.A1(_04995_),
    .A2(_04994_),
    .B1(_04454_),
    .Y(_04996_));
 sky130_fd_sc_hd__a31o_2 _19721_ (.A1(_04992_),
    .A2(_04993_),
    .A3(_04994_),
    .B1(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__nor2_2 _19722_ (.A(_04974_),
    .B(_04977_),
    .Y(_04998_));
 sky130_fd_sc_hd__a21oi_2 _19723_ (.A1(_03888_),
    .A2(_03893_),
    .B1(_04998_),
    .Y(_04999_));
 sky130_fd_sc_hd__o31a_2 _19724_ (.A1(_03894_),
    .A2(_04195_),
    .A3(_04998_),
    .B1(_04496_),
    .X(_05000_));
 sky130_fd_sc_hd__o21ai_2 _19725_ (.A1(_04995_),
    .A2(_04999_),
    .B1(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__o211ai_2 _19726_ (.A1(_04408_),
    .A2(_04992_),
    .B1(_04993_),
    .C1(_04445_),
    .Y(_05002_));
 sky130_fd_sc_hd__o31a_2 _19727_ (.A1(_03639_),
    .A2(_04991_),
    .A3(_03881_),
    .B1(_04589_),
    .X(_05003_));
 sky130_fd_sc_hd__a41o_2 _19728_ (.A1(_04465_),
    .A2(_04997_),
    .A3(_05001_),
    .A4(_05002_),
    .B1(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__or3b_2 _19729_ (.A(_04295_),
    .B(_04362_),
    .C_N(_04629_),
    .X(_05005_));
 sky130_fd_sc_hd__mux2_2 _19730_ (.A0(_03888_),
    .A1(_03872_),
    .S(_04274_),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_2 _19731_ (.A0(_05006_),
    .A1(_04964_),
    .S(_04352_),
    .X(_05007_));
 sky130_fd_sc_hd__mux2_2 _19732_ (.A0(_05007_),
    .A1(_04919_),
    .S(_04269_),
    .X(_05008_));
 sky130_fd_sc_hd__or4b_2 _19733_ (.A(_04038_),
    .B(_04537_),
    .C(_04301_),
    .D_N(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__o31a_2 _19734_ (.A1(_04349_),
    .A2(_04303_),
    .A3(_04816_),
    .B1(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__o311a_2 _19735_ (.A1(_04546_),
    .A2(_04626_),
    .A3(_04924_),
    .B1(_04515_),
    .C1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__o32a_2 _19736_ (.A1(_04618_),
    .A2(_04245_),
    .A3(_04386_),
    .B1(_04515_),
    .B2(_03705_),
    .X(_05012_));
 sky130_fd_sc_hd__o221ai_2 _19737_ (.A1(_04805_),
    .A2(_04806_),
    .B1(_05012_),
    .B2(_04628_),
    .C1(_04729_),
    .Y(_05013_));
 sky130_fd_sc_hd__a31oi_2 _19738_ (.A1(_05004_),
    .A2(_05005_),
    .A3(_05011_),
    .B1(_05013_),
    .Y(_00571_));
 sky130_fd_sc_hd__and4_2 _19739_ (.A(_04974_),
    .B(_04995_),
    .C(_04191_),
    .D(_04192_),
    .X(_05014_));
 sky130_fd_sc_hd__inv_2 _19740_ (.A(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__o21bai_2 _19741_ (.A1(_04931_),
    .A2(_04929_),
    .B1_N(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__a21bo_2 _19742_ (.A1(_04982_),
    .A2(_04993_),
    .B1_N(_04992_),
    .X(_05017_));
 sky130_fd_sc_hd__a31oi_2 _19743_ (.A1(_04974_),
    .A2(_04972_),
    .A3(_04995_),
    .B1(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__a21oi_2 _19744_ (.A1(_05016_),
    .A2(_05018_),
    .B1(_03851_),
    .Y(_05019_));
 sky130_fd_sc_hd__a31o_2 _19745_ (.A1(_05016_),
    .A2(_05018_),
    .A3(_03851_),
    .B1(_04525_),
    .X(_05020_));
 sky130_fd_sc_hd__o21ba_2 _19746_ (.A1(_03894_),
    .A2(_03882_),
    .B1_N(_04194_),
    .X(_05021_));
 sky130_fd_sc_hd__o21ai_2 _19747_ (.A1(_03924_),
    .A2(_03937_),
    .B1(_03903_),
    .Y(_05022_));
 sky130_fd_sc_hd__a21oi_2 _19748_ (.A1(_03912_),
    .A2(_04863_),
    .B1(_04935_),
    .Y(_05023_));
 sky130_fd_sc_hd__o2111a_2 _19749_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_04190_),
    .C1(_04195_),
    .D1(_04193_),
    .X(_05024_));
 sky130_fd_sc_hd__a311o_2 _19750_ (.A1(_04190_),
    .A2(_04195_),
    .A3(_03963_),
    .B1(_05021_),
    .C1(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__a31o_2 _19751_ (.A1(_04840_),
    .A2(_04212_),
    .A3(_04196_),
    .B1(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__o21ai_2 _19752_ (.A1(_03851_),
    .A2(_05026_),
    .B1(_04495_),
    .Y(_05027_));
 sky130_fd_sc_hd__a21o_2 _19753_ (.A1(_03851_),
    .A2(_05026_),
    .B1(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__o211a_2 _19754_ (.A1(_05019_),
    .A2(_05020_),
    .B1(_05028_),
    .C1(_04667_),
    .X(_05029_));
 sky130_fd_sc_hd__o211a_2 _19755_ (.A1(_03847_),
    .A2(_04442_),
    .B1(_04444_),
    .C1(_03851_),
    .X(_05030_));
 sky130_fd_sc_hd__and2b_2 _19756_ (.A_N(_03847_),
    .B(_03844_),
    .X(_05031_));
 sky130_fd_sc_hd__o21ai_2 _19757_ (.A1(_04503_),
    .A2(_05031_),
    .B1(_04589_),
    .Y(_05032_));
 sky130_fd_sc_hd__o21ai_2 _19758_ (.A1(_05029_),
    .A2(_05030_),
    .B1(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__mux2_2 _19759_ (.A0(_03872_),
    .A1(_03844_),
    .S(_04307_),
    .X(_05034_));
 sky130_fd_sc_hd__o211a_2 _19760_ (.A1(_03888_),
    .A2(_04320_),
    .B1(_04265_),
    .C1(_04249_),
    .X(_05035_));
 sky130_fd_sc_hd__a21oi_2 _19761_ (.A1(_04325_),
    .A2(_05034_),
    .B1(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__o22ai_2 _19762_ (.A1(_04305_),
    .A2(_05036_),
    .B1(_04371_),
    .B2(_04851_),
    .Y(_05037_));
 sky130_fd_sc_hd__a211o_2 _19763_ (.A1(_04330_),
    .A2(_04945_),
    .B1(_05037_),
    .C1(_04303_),
    .X(_05038_));
 sky130_fd_sc_hd__o311a_2 _19764_ (.A1(_04508_),
    .A2(_04301_),
    .A3(_04650_),
    .B1(_05033_),
    .C1(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__and3_2 _19765_ (.A(_04508_),
    .B(_04415_),
    .C(_04654_),
    .X(_05040_));
 sky130_fd_sc_hd__o311a_2 _19766_ (.A1(_04442_),
    .A2(_04245_),
    .A3(_04386_),
    .B1(_04806_),
    .C1(_04728_),
    .X(_05041_));
 sky130_fd_sc_hd__a31o_2 _19767_ (.A1(_04805_),
    .A2(_04654_),
    .A3(_04729_),
    .B1(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__o31a_2 _19768_ (.A1(_04949_),
    .A2(_05039_),
    .A3(_05040_),
    .B1(_05042_),
    .X(_00572_));
 sky130_fd_sc_hd__and3_2 _19769_ (.A(_04509_),
    .B(_04369_),
    .C(_04905_),
    .X(_05043_));
 sky130_fd_sc_hd__a31o_2 _19770_ (.A1(_04442_),
    .A2(_03852_),
    .A3(_03839_),
    .B1(_04667_),
    .X(_05044_));
 sky130_fd_sc_hd__nand2_2 _19771_ (.A(_03852_),
    .B(_03839_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand2_2 _19772_ (.A(_05026_),
    .B(_03851_),
    .Y(_05046_));
 sky130_fd_sc_hd__and3_2 _19773_ (.A(_03849_),
    .B(_05045_),
    .C(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__nand2_2 _19774_ (.A(_05026_),
    .B(_03853_),
    .Y(_05048_));
 sky130_fd_sc_hd__or2_2 _19775_ (.A(_03849_),
    .B(_05045_),
    .X(_05049_));
 sky130_fd_sc_hd__and4b_2 _19776_ (.A_N(_05047_),
    .B(_04495_),
    .C(_05048_),
    .D(_05049_),
    .X(_05050_));
 sky130_fd_sc_hd__a21o_2 _19777_ (.A1(_03852_),
    .A2(_03839_),
    .B1(_03851_),
    .X(_05051_));
 sky130_fd_sc_hd__a21oi_2 _19778_ (.A1(_05016_),
    .A2(_05018_),
    .B1(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__a211oi_2 _19779_ (.A1(_05045_),
    .A2(_05031_),
    .B1(_04525_),
    .C1(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__or4_2 _19780_ (.A(_05045_),
    .B(_04495_),
    .C(_05019_),
    .D(_05031_),
    .X(_05054_));
 sky130_fd_sc_hd__o221ai_2 _19781_ (.A1(_04225_),
    .A2(_04667_),
    .B1(_05050_),
    .B2(_05053_),
    .C1(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__buf_1 _19782_ (.A(_04297_),
    .X(_05056_));
 sky130_fd_sc_hd__a211o_2 _19783_ (.A1(_05056_),
    .A2(\decode.id_ex_imm_reg[25] ),
    .B1(_04388_),
    .C1(_03837_),
    .X(_05057_));
 sky130_fd_sc_hd__o2bb2ai_2 _19784_ (.A1_N(_05044_),
    .A2_N(_05055_),
    .B1(_03835_),
    .B2(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__nand2_2 _19785_ (.A(_04620_),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__and2b_2 _19786_ (.A_N(_03838_),
    .B(_03835_),
    .X(_05060_));
 sky130_fd_sc_hd__mux2_2 _19787_ (.A0(_03835_),
    .A1(_03844_),
    .S(_04234_),
    .X(_05061_));
 sky130_fd_sc_hd__a211o_2 _19788_ (.A1(_04297_),
    .A2(_04261_),
    .B1(_04263_),
    .C1(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__o211a_2 _19789_ (.A1(_04325_),
    .A2(_05006_),
    .B1(_04317_),
    .C1(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__a221o_2 _19790_ (.A1(_04330_),
    .A2(_04965_),
    .B1(_04877_),
    .B2(_04537_),
    .C1(_04302_),
    .X(_05064_));
 sky130_fd_sc_hd__o32a_2 _19791_ (.A1(_04225_),
    .A2(_04424_),
    .A3(_05060_),
    .B1(_05063_),
    .B2(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__o211a_2 _19792_ (.A1(_04675_),
    .A2(_04924_),
    .B1(_04360_),
    .C1(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__a221oi_2 _19793_ (.A1(_04439_),
    .A2(_04679_),
    .B1(_05059_),
    .B2(_05066_),
    .C1(_04949_),
    .Y(_05067_));
 sky130_fd_sc_hd__o21bai_2 _19794_ (.A1(_05041_),
    .A2(_05043_),
    .B1_N(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__inv_2 _19795_ (.A(_05068_),
    .Y(_00573_));
 sky130_fd_sc_hd__a2111o_2 _19796_ (.A1(_03772_),
    .A2(_10116_),
    .B1(_03775_),
    .C1(_03806_),
    .D1(_03809_),
    .X(_05069_));
 sky130_fd_sc_hd__mux2_2 _19797_ (.A0(_03835_),
    .A1(_03812_),
    .S(_04274_),
    .X(_05070_));
 sky130_fd_sc_hd__a211o_2 _19798_ (.A1(_04297_),
    .A2(_04261_),
    .B1(_04263_),
    .C1(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__o21ai_2 _19799_ (.A1(_04325_),
    .A2(_05034_),
    .B1(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__a2bb2o_2 _19800_ (.A1_N(_04304_),
    .A2_N(_05072_),
    .B1(_04537_),
    .B2(_04898_),
    .X(_05073_));
 sky130_fd_sc_hd__a211oi_2 _19801_ (.A1(_04330_),
    .A2(_04984_),
    .B1(_05073_),
    .C1(_04302_),
    .Y(_05074_));
 sky130_fd_sc_hd__a311o_2 _19802_ (.A1(_04618_),
    .A2(_05069_),
    .A3(_04589_),
    .B1(_04492_),
    .C1(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__a21o_2 _19803_ (.A1(_05045_),
    .A2(_05031_),
    .B1(_05060_),
    .X(_05076_));
 sky130_fd_sc_hd__o31a_2 _19804_ (.A1(_03814_),
    .A2(_05076_),
    .A3(_05052_),
    .B1(_04400_),
    .X(_05077_));
 sky130_fd_sc_hd__o21ai_2 _19805_ (.A1(_05076_),
    .A2(_05052_),
    .B1(_03814_),
    .Y(_05078_));
 sky130_fd_sc_hd__a31o_2 _19806_ (.A1(_03852_),
    .A2(_05048_),
    .A3(_05049_),
    .B1(_03814_),
    .X(_05079_));
 sky130_fd_sc_hd__o2111ai_2 _19807_ (.A1(_05045_),
    .A2(_05046_),
    .B1(_05049_),
    .C1(_03814_),
    .D1(_03852_),
    .Y(_05080_));
 sky130_fd_sc_hd__and3_2 _19808_ (.A(_05079_),
    .B(_04495_),
    .C(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__a211o_2 _19809_ (.A1(_05077_),
    .A2(_05078_),
    .B1(_04445_),
    .C1(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__a211o_2 _19810_ (.A1(_03810_),
    .A2(_03639_),
    .B1(_04667_),
    .C1(_03814_),
    .X(_05083_));
 sky130_fd_sc_hd__a21oi_2 _19811_ (.A1(_05082_),
    .A2(_05083_),
    .B1(_04589_),
    .Y(_05084_));
 sky130_fd_sc_hd__a211oi_2 _19812_ (.A1(_04693_),
    .A2(_04879_),
    .B1(_05075_),
    .C1(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__and3_2 _19813_ (.A(_04508_),
    .B(_04415_),
    .C(_04700_),
    .X(_05086_));
 sky130_fd_sc_hd__a41o_2 _19814_ (.A1(_03705_),
    .A2(_04509_),
    .A3(_04332_),
    .A4(_04412_),
    .B1(_04700_),
    .X(_05087_));
 sky130_fd_sc_hd__a31o_2 _19815_ (.A1(_04805_),
    .A2(_05087_),
    .A3(_04729_),
    .B1(_05041_),
    .X(_05088_));
 sky130_fd_sc_hd__o31a_2 _19816_ (.A1(_04949_),
    .A2(_05085_),
    .A3(_05086_),
    .B1(_05088_),
    .X(_00574_));
 sky130_fd_sc_hd__a31o_2 _19817_ (.A1(_04471_),
    .A2(_04439_),
    .A3(_04509_),
    .B1(_04949_),
    .X(_05089_));
 sky130_fd_sc_hd__a2111o_2 _19818_ (.A1(_03819_),
    .A2(_03817_),
    .B1(_03775_),
    .C1(_03820_),
    .D1(_03825_),
    .X(_05090_));
 sky130_fd_sc_hd__mux2_2 _19819_ (.A0(_03821_),
    .A1(_03812_),
    .S(_04254_),
    .X(_05091_));
 sky130_fd_sc_hd__a211o_2 _19820_ (.A1(_04297_),
    .A2(_04261_),
    .B1(_04263_),
    .C1(_05091_),
    .X(_05092_));
 sky130_fd_sc_hd__o21ai_2 _19821_ (.A1(_04338_),
    .A2(_05061_),
    .B1(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__o2bb2a_2 _19822_ (.A1_N(_04330_),
    .A2_N(_05007_),
    .B1(_04304_),
    .B2(_05093_),
    .X(_05094_));
 sky130_fd_sc_hd__o211a_2 _19823_ (.A1(_04921_),
    .A2(_04371_),
    .B1(_04392_),
    .C1(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__a31o_2 _19824_ (.A1(_04618_),
    .A2(_04589_),
    .A3(_05090_),
    .B1(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__nor2_2 _19825_ (.A(_04708_),
    .B(_04924_),
    .Y(_05097_));
 sky130_fd_sc_hd__inv_2 _19826_ (.A(_03825_),
    .Y(_05098_));
 sky130_fd_sc_hd__a211o_2 _19827_ (.A1(_05098_),
    .A2(_03639_),
    .B1(_04667_),
    .C1(_03829_),
    .X(_05099_));
 sky130_fd_sc_hd__nand2_2 _19828_ (.A(_03814_),
    .B(_03829_),
    .Y(_05100_));
 sky130_fd_sc_hd__o21bai_2 _19829_ (.A1(_05076_),
    .A2(_05052_),
    .B1_N(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__nand3_2 _19830_ (.A(_03829_),
    .B(_03812_),
    .C(_03810_),
    .Y(_05102_));
 sky130_fd_sc_hd__and3_2 _19831_ (.A(_05101_),
    .B(_05102_),
    .C(_04400_),
    .X(_05103_));
 sky130_fd_sc_hd__nand3b_2 _19832_ (.A_N(_03829_),
    .B(_05078_),
    .C(_05069_),
    .Y(_05104_));
 sky130_fd_sc_hd__a21oi_2 _19833_ (.A1(_03811_),
    .A2(_05079_),
    .B1(_03829_),
    .Y(_05105_));
 sky130_fd_sc_hd__and3_2 _19834_ (.A(_03811_),
    .B(_03829_),
    .C(_05079_),
    .X(_05106_));
 sky130_fd_sc_hd__o31a_2 _19835_ (.A1(_05105_),
    .A2(_04401_),
    .A3(_05106_),
    .B1(_04504_),
    .X(_05107_));
 sky130_fd_sc_hd__a21bo_2 _19836_ (.A1(_05103_),
    .A2(_05104_),
    .B1_N(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__a21oi_2 _19837_ (.A1(_05099_),
    .A2(_05108_),
    .B1(_04589_),
    .Y(_05109_));
 sky130_fd_sc_hd__nor4_2 _19838_ (.A(_04492_),
    .B(_05096_),
    .C(_05097_),
    .D(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__and3_2 _19839_ (.A(_04509_),
    .B(_04905_),
    .C(_04511_),
    .X(_05111_));
 sky130_fd_sc_hd__o22a_2 _19840_ (.A1(_05089_),
    .A2(_05110_),
    .B1(_05111_),
    .B2(_05041_),
    .X(_00575_));
 sky130_fd_sc_hd__a21o_2 _19841_ (.A1(_03705_),
    .A2(_04305_),
    .B1(_04751_),
    .X(_05112_));
 sky130_fd_sc_hd__and3_2 _19842_ (.A(_04508_),
    .B(_04728_),
    .C(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__a31o_2 _19843_ (.A1(_04805_),
    .A2(_04415_),
    .A3(_04751_),
    .B1(_04949_),
    .X(_05114_));
 sky130_fd_sc_hd__mux2_2 _19844_ (.A0(_03821_),
    .A1(_03795_),
    .S(_04274_),
    .X(_05115_));
 sky130_fd_sc_hd__a211o_2 _19845_ (.A1(_05056_),
    .A2(_04261_),
    .B1(_04263_),
    .C1(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__o211a_2 _19846_ (.A1(_04325_),
    .A2(_05070_),
    .B1(_04317_),
    .C1(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__a2bb2o_2 _19847_ (.A1_N(_04436_),
    .A2_N(_05036_),
    .B1(_04409_),
    .B2(_04947_),
    .X(_05118_));
 sky130_fd_sc_hd__o31a_2 _19848_ (.A1(_04303_),
    .A2(_05117_),
    .A3(_05118_),
    .B1(_04360_),
    .X(_05119_));
 sky130_fd_sc_hd__a2111o_2 _19849_ (.A1(_03772_),
    .A2(_10127_),
    .B1(_03775_),
    .C1(_03794_),
    .D1(_03800_),
    .X(_05120_));
 sky130_fd_sc_hd__a211oi_2 _19850_ (.A1(_03639_),
    .A2(_03795_),
    .B1(_03803_),
    .C1(_04667_),
    .Y(_05121_));
 sky130_fd_sc_hd__a32oi_2 _19851_ (.A1(_03829_),
    .A2(_03812_),
    .A3(_03810_),
    .B1(_05098_),
    .B2(_03821_),
    .Y(_05122_));
 sky130_fd_sc_hd__nand2_2 _19852_ (.A(_05101_),
    .B(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__a21oi_2 _19853_ (.A1(_03803_),
    .A2(_05123_),
    .B1(_04526_),
    .Y(_05124_));
 sky130_fd_sc_hd__nand4_2 _19854_ (.A(_05122_),
    .B(_05101_),
    .C(_03802_),
    .D(_03801_),
    .Y(_05125_));
 sky130_fd_sc_hd__o211ai_2 _19855_ (.A1(_05045_),
    .A2(_05046_),
    .B1(_05049_),
    .C1(_03852_),
    .Y(_05126_));
 sky130_fd_sc_hd__a21oi_2 _19856_ (.A1(_05126_),
    .A2(_03830_),
    .B1(_04219_),
    .Y(_05127_));
 sky130_fd_sc_hd__or2_2 _19857_ (.A(_03803_),
    .B(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__a221o_2 _19858_ (.A1(_03801_),
    .A2(_03802_),
    .B1(_05126_),
    .B2(_03830_),
    .C1(_04219_),
    .X(_05129_));
 sky130_fd_sc_hd__a31o_2 _19859_ (.A1(_05128_),
    .A2(_04495_),
    .A3(_05129_),
    .B1(_04444_),
    .X(_05130_));
 sky130_fd_sc_hd__a21oi_2 _19860_ (.A1(_05124_),
    .A2(_05125_),
    .B1(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__o221ai_2 _19861_ (.A1(_04620_),
    .A2(_05120_),
    .B1(_05121_),
    .B2(_05131_),
    .C1(_04301_),
    .Y(_05132_));
 sky130_fd_sc_hd__o311a_2 _19862_ (.A1(_04508_),
    .A2(_04301_),
    .A3(_04736_),
    .B1(_05119_),
    .C1(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__o22a_2 _19863_ (.A1(_04883_),
    .A2(_05113_),
    .B1(_05114_),
    .B2(_05133_),
    .X(_00576_));
 sky130_fd_sc_hd__or3_2 _19864_ (.A(_04295_),
    .B(_04775_),
    .C(_04779_),
    .X(_05134_));
 sky130_fd_sc_hd__o21ai_2 _19865_ (.A1(_04338_),
    .A2(_05006_),
    .B1(_05062_),
    .Y(_05135_));
 sky130_fd_sc_hd__o2bb2a_2 _19866_ (.A1_N(_04243_),
    .A2_N(_04966_),
    .B1(_05135_),
    .B2(_04436_),
    .X(_05136_));
 sky130_fd_sc_hd__a21oi_2 _19867_ (.A1(_03795_),
    .A2(_04320_),
    .B1(_04366_),
    .Y(_05137_));
 sky130_fd_sc_hd__a21oi_2 _19868_ (.A1(_04251_),
    .A2(_04252_),
    .B1(_05091_),
    .Y(_05138_));
 sky130_fd_sc_hd__a311o_2 _19869_ (.A1(_04251_),
    .A2(_04252_),
    .A3(_05137_),
    .B1(_04304_),
    .C1(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__a31o_2 _19870_ (.A1(_04392_),
    .A2(_05136_),
    .A3(_05139_),
    .B1(_04492_),
    .X(_05140_));
 sky130_fd_sc_hd__a41o_2 _19871_ (.A1(_04503_),
    .A2(_04772_),
    .A3(_04294_),
    .A4(_04391_),
    .B1(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__a21o_2 _19872_ (.A1(_04297_),
    .A2(\decode.id_ex_imm_reg[29] ),
    .B1(_03787_),
    .X(_05142_));
 sky130_fd_sc_hd__a21o_2 _19873_ (.A1(_05142_),
    .A2(_03781_),
    .B1(_04225_),
    .X(_05143_));
 sky130_fd_sc_hd__or3b_2 _19874_ (.A(_03789_),
    .B(_03790_),
    .C_N(_05120_),
    .X(_05144_));
 sky130_fd_sc_hd__a21oi_2 _19875_ (.A1(_03803_),
    .A2(_05123_),
    .B1(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__o21ba_2 _19876_ (.A1(_03789_),
    .A2(_03790_),
    .B1_N(_05120_),
    .X(_05146_));
 sky130_fd_sc_hd__or2_2 _19877_ (.A(_04525_),
    .B(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__a31o_2 _19878_ (.A1(_03791_),
    .A2(_03803_),
    .A3(_05123_),
    .B1(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__o221a_2 _19879_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03803_),
    .B2(_05127_),
    .C1(_03802_),
    .X(_05149_));
 sky130_fd_sc_hd__a21oi_2 _19880_ (.A1(_03802_),
    .A2(_05128_),
    .B1(_03791_),
    .Y(_05150_));
 sky130_fd_sc_hd__o31a_2 _19881_ (.A1(_05149_),
    .A2(_04401_),
    .A3(_05150_),
    .B1(_04504_),
    .X(_05151_));
 sky130_fd_sc_hd__o21ai_2 _19882_ (.A1(_05145_),
    .A2(_05148_),
    .B1(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__o21ai_2 _19883_ (.A1(_04359_),
    .A2(_03788_),
    .B1(_04444_),
    .Y(_05153_));
 sky130_fd_sc_hd__o31a_2 _19884_ (.A1(_03789_),
    .A2(_03790_),
    .A3(_05153_),
    .B1(_04465_),
    .X(_05154_));
 sky130_fd_sc_hd__a22oi_2 _19885_ (.A1(_04589_),
    .A2(_05143_),
    .B1(_05152_),
    .B2(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__o221a_2 _19886_ (.A1(_04386_),
    .A2(_04776_),
    .B1(_05141_),
    .B2(_05155_),
    .C1(_04515_),
    .X(_05156_));
 sky130_fd_sc_hd__a21oi_2 _19887_ (.A1(_04856_),
    .A2(_05134_),
    .B1(_05156_),
    .Y(_00577_));
 sky130_fd_sc_hd__o211a_2 _19888_ (.A1(_04799_),
    .A2(_04798_),
    .B1(_04805_),
    .C1(_04729_),
    .X(_05157_));
 sky130_fd_sc_hd__o211ai_2 _19889_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03803_),
    .C1(_05123_),
    .Y(_05158_));
 sky130_fd_sc_hd__a21oi_2 _19890_ (.A1(_03781_),
    .A2(_05142_),
    .B1(_05146_),
    .Y(_05159_));
 sky130_fd_sc_hd__a31oi_2 _19891_ (.A1(_05158_),
    .A2(_05159_),
    .A3(_03865_),
    .B1(_04526_),
    .Y(_05160_));
 sky130_fd_sc_hd__o2bb2ai_2 _19892_ (.A1_N(_05159_),
    .A2_N(_05158_),
    .B1(_03864_),
    .B2(_03862_),
    .Y(_05161_));
 sky130_fd_sc_hd__a21oi_2 _19893_ (.A1(_03802_),
    .A2(_05128_),
    .B1(_03789_),
    .Y(_05162_));
 sky130_fd_sc_hd__a211oi_2 _19894_ (.A1(_03781_),
    .A2(_03788_),
    .B1(_03865_),
    .C1(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__o21a_2 _19895_ (.A1(_03790_),
    .A2(_05162_),
    .B1(_03865_),
    .X(_05164_));
 sky130_fd_sc_hd__o31ai_2 _19896_ (.A1(_04452_),
    .A2(_05163_),
    .A3(_05164_),
    .B1(_04505_),
    .Y(_05165_));
 sky130_fd_sc_hd__a21oi_2 _19897_ (.A1(_05160_),
    .A2(_05161_),
    .B1(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__o211a_2 _19898_ (.A1(_03861_),
    .A2(_04618_),
    .B1(_04445_),
    .C1(_03865_),
    .X(_05167_));
 sky130_fd_sc_hd__o21ai_2 _19899_ (.A1(_05166_),
    .A2(_05167_),
    .B1(_04620_),
    .Y(_05168_));
 sky130_fd_sc_hd__or2b_2 _19900_ (.A(_03861_),
    .B_N(_03863_),
    .X(_05169_));
 sky130_fd_sc_hd__mux2_2 _19901_ (.A0(_03863_),
    .A1(_03781_),
    .S(_04254_),
    .X(_05170_));
 sky130_fd_sc_hd__mux2_2 _19902_ (.A0(_05170_),
    .A1(_05115_),
    .S(_04248_),
    .X(_05171_));
 sky130_fd_sc_hd__a22oi_2 _19903_ (.A1(_04317_),
    .A2(_05171_),
    .B1(_04985_),
    .B2(_04537_),
    .Y(_05172_));
 sky130_fd_sc_hd__o211a_2 _19904_ (.A1(_04436_),
    .A2(_05072_),
    .B1(_05172_),
    .C1(_04392_),
    .X(_05173_));
 sky130_fd_sc_hd__a221o_2 _19905_ (.A1(_04425_),
    .A2(_05169_),
    .B1(_04794_),
    .B2(_04879_),
    .C1(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__a21oi_2 _19906_ (.A1(_04443_),
    .A2(_04415_),
    .B1(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__a31o_2 _19907_ (.A1(_04317_),
    .A2(_04439_),
    .A3(_04410_),
    .B1(_04949_),
    .X(_05176_));
 sky130_fd_sc_hd__a21o_2 _19908_ (.A1(_05168_),
    .A2(_05175_),
    .B1(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__o21ai_2 _19909_ (.A1(_05041_),
    .A2(_05157_),
    .B1(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__inv_2 _19910_ (.A(_05178_),
    .Y(_00578_));
 sky130_fd_sc_hd__a21oi_2 _19911_ (.A1(_03704_),
    .A2(_04338_),
    .B1(_04320_),
    .Y(_05179_));
 sky130_fd_sc_hd__o22a_2 _19912_ (.A1(_04325_),
    .A2(_05137_),
    .B1(_05179_),
    .B2(_04572_),
    .X(_05180_));
 sky130_fd_sc_hd__o2bb2a_2 _19913_ (.A1_N(_04244_),
    .A2_N(_05008_),
    .B1(_05180_),
    .B2(_04305_),
    .X(_05181_));
 sky130_fd_sc_hd__o211a_2 _19914_ (.A1(_05093_),
    .A2(_04436_),
    .B1(_04428_),
    .C1(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__a221o_2 _19915_ (.A1(_04443_),
    .A2(_04242_),
    .B1(_04817_),
    .B2(_04879_),
    .C1(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__nand2_2 _19916_ (.A(_03854_),
    .B(_05169_),
    .Y(_05184_));
 sky130_fd_sc_hd__inv_2 _19917_ (.A(_03862_),
    .Y(_05185_));
 sky130_fd_sc_hd__a22oi_2 _19918_ (.A1(_05185_),
    .A2(_04215_),
    .B1(_05158_),
    .B2(_05159_),
    .Y(_05186_));
 sky130_fd_sc_hd__o21bai_2 _19919_ (.A1(_05184_),
    .A2(_05186_),
    .B1_N(_04526_),
    .Y(_05187_));
 sky130_fd_sc_hd__a21oi_2 _19920_ (.A1(_05161_),
    .A2(_05169_),
    .B1(_03854_),
    .Y(_05188_));
 sky130_fd_sc_hd__o21a_2 _19921_ (.A1(_03862_),
    .A2(_05164_),
    .B1(_03854_),
    .X(_05189_));
 sky130_fd_sc_hd__o31ai_2 _19922_ (.A1(_03854_),
    .A2(_03862_),
    .A3(_05164_),
    .B1(_04496_),
    .Y(_05190_));
 sky130_fd_sc_hd__o21ai_2 _19923_ (.A1(_05189_),
    .A2(_05190_),
    .B1(_04505_),
    .Y(_05191_));
 sky130_fd_sc_hd__o21bai_2 _19924_ (.A1(_05187_),
    .A2(_05188_),
    .B1_N(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__o21ai_2 _19925_ (.A1(_04442_),
    .A2(_03766_),
    .B1(_03854_),
    .Y(_05193_));
 sky130_fd_sc_hd__o22a_2 _19926_ (.A1(_04620_),
    .A2(_04408_),
    .B1(_04505_),
    .B2(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__or4b_2 _19927_ (.A(_04225_),
    .B(_03766_),
    .C(_04424_),
    .D_N(_03705_),
    .X(_05195_));
 sky130_fd_sc_hd__o21ai_2 _19928_ (.A1(_04443_),
    .A2(_04620_),
    .B1(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__a21oi_2 _19929_ (.A1(_05192_),
    .A2(_05194_),
    .B1(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__a31o_2 _19930_ (.A1(_04317_),
    .A2(_04439_),
    .A3(_04468_),
    .B1(_04949_),
    .X(_05198_));
 sky130_fd_sc_hd__o21bai_2 _19931_ (.A1(_05183_),
    .A2(_05197_),
    .B1_N(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__nand2_2 _19932_ (.A(_05199_),
    .B(_04855_),
    .Y(_05200_));
 sky130_fd_sc_hd__inv_2 _19933_ (.A(_05200_),
    .Y(_00579_));
 sky130_fd_sc_hd__nor2_2 _19934_ (.A(_03588_),
    .B(_04238_),
    .Y(_00580_));
 sky130_fd_sc_hd__buf_1 _19935_ (.A(_09955_),
    .X(_05201_));
 sky130_fd_sc_hd__and3b_2 _19936_ (.A_N(_03581_),
    .B(_05201_),
    .C(\decode.id_ex_memtoreg_reg[0] ),
    .X(_05202_));
 sky130_fd_sc_hd__buf_1 _19937_ (.A(_05202_),
    .X(_00581_));
 sky130_fd_sc_hd__and3b_2 _19938_ (.A_N(_03581_),
    .B(_05201_),
    .C(\decode.id_ex_memtoreg_reg[1] ),
    .X(_05203_));
 sky130_fd_sc_hd__buf_1 _19939_ (.A(_05203_),
    .X(_00582_));
 sky130_fd_sc_hd__and3b_2 _19940_ (.A_N(_03581_),
    .B(_05201_),
    .C(\decode.id_ex_regwrite_reg ),
    .X(_05204_));
 sky130_fd_sc_hd__buf_1 _19941_ (.A(_05204_),
    .X(_00583_));
 sky130_fd_sc_hd__and3b_2 _19942_ (.A_N(_03581_),
    .B(_05201_),
    .C(\decode.id_ex_memwrite_reg ),
    .X(_05205_));
 sky130_fd_sc_hd__buf_1 _19943_ (.A(_05205_),
    .X(_00584_));
 sky130_fd_sc_hd__buf_1 _19944_ (.A(\decode.id_ex_memread_reg ),
    .X(_05206_));
 sky130_fd_sc_hd__and2_2 _19945_ (.A(_05206_),
    .B(_03627_),
    .X(_05207_));
 sky130_fd_sc_hd__buf_1 _19946_ (.A(_05207_),
    .X(_00585_));
 sky130_fd_sc_hd__and3b_2 _19947_ (.A_N(_03581_),
    .B(_05201_),
    .C(\decode.id_ex_isjump_reg ),
    .X(_05208_));
 sky130_fd_sc_hd__buf_1 _19948_ (.A(_05208_),
    .X(_00586_));
 sky130_fd_sc_hd__and3b_2 _19949_ (.A_N(_03581_),
    .B(_05201_),
    .C(\decode.id_ex_isbranch_reg ),
    .X(_05209_));
 sky130_fd_sc_hd__buf_1 _19950_ (.A(_05209_),
    .X(_00587_));
 sky130_fd_sc_hd__and2_2 _19951_ (.A(\decode.id_ex_pc_reg[0] ),
    .B(_03627_),
    .X(_05210_));
 sky130_fd_sc_hd__buf_1 _19952_ (.A(_05210_),
    .X(_00588_));
 sky130_fd_sc_hd__and2_2 _19953_ (.A(\decode.id_ex_pc_reg[1] ),
    .B(_03627_),
    .X(_05211_));
 sky130_fd_sc_hd__buf_1 _19954_ (.A(_05211_),
    .X(_00589_));
 sky130_fd_sc_hd__nor2_2 _19955_ (.A(_10711_),
    .B(_03599_),
    .Y(_00590_));
 sky130_fd_sc_hd__nor2_2 _19956_ (.A(_10748_),
    .B(_03599_),
    .Y(_00591_));
 sky130_fd_sc_hd__nor2_2 _19957_ (.A(_10690_),
    .B(_03599_),
    .Y(_00592_));
 sky130_fd_sc_hd__nor2_2 _19958_ (.A(_10705_),
    .B(_03599_),
    .Y(_00593_));
 sky130_fd_sc_hd__and2_2 _19959_ (.A(_10678_),
    .B(_03627_),
    .X(_05212_));
 sky130_fd_sc_hd__buf_1 _19960_ (.A(_05212_),
    .X(_00594_));
 sky130_fd_sc_hd__nor2_2 _19961_ (.A(_10731_),
    .B(_03599_),
    .Y(_00595_));
 sky130_fd_sc_hd__nor2_2 _19962_ (.A(_10680_),
    .B(_03599_),
    .Y(_00596_));
 sky130_fd_sc_hd__nor2_2 _19963_ (.A(_10707_),
    .B(_03599_),
    .Y(_00597_));
 sky130_fd_sc_hd__nor2_2 _19964_ (.A(_10721_),
    .B(_03599_),
    .Y(_00598_));
 sky130_fd_sc_hd__and2_2 _19965_ (.A(_10689_),
    .B(_03627_),
    .X(_05213_));
 sky130_fd_sc_hd__buf_1 _19966_ (.A(_05213_),
    .X(_00599_));
 sky130_fd_sc_hd__buf_1 _19967_ (.A(_03594_),
    .X(_05214_));
 sky130_fd_sc_hd__and2_2 _19968_ (.A(_10694_),
    .B(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__buf_1 _19969_ (.A(_05215_),
    .X(_00600_));
 sky130_fd_sc_hd__and2_2 _19970_ (.A(_10710_),
    .B(_05214_),
    .X(_05216_));
 sky130_fd_sc_hd__buf_1 _19971_ (.A(_05216_),
    .X(_00601_));
 sky130_fd_sc_hd__nor2_2 _19972_ (.A(_10702_),
    .B(_03599_),
    .Y(_00602_));
 sky130_fd_sc_hd__buf_1 _19973_ (.A(_03588_),
    .X(_05217_));
 sky130_fd_sc_hd__nor2_2 _19974_ (.A(_10682_),
    .B(_05217_),
    .Y(_00603_));
 sky130_fd_sc_hd__nor2_2 _19975_ (.A(_10675_),
    .B(_05217_),
    .Y(_00604_));
 sky130_fd_sc_hd__nor2_2 _19976_ (.A(_10736_),
    .B(_05217_),
    .Y(_00605_));
 sky130_fd_sc_hd__nor2_2 _19977_ (.A(_10713_),
    .B(_05217_),
    .Y(_00606_));
 sky130_fd_sc_hd__nor2_2 _19978_ (.A(_10692_),
    .B(_05217_),
    .Y(_00607_));
 sky130_fd_sc_hd__nor2_2 _19979_ (.A(_10716_),
    .B(_05217_),
    .Y(_00608_));
 sky130_fd_sc_hd__and2_2 _19980_ (.A(_10798_),
    .B(_05214_),
    .X(_05218_));
 sky130_fd_sc_hd__buf_1 _19981_ (.A(_05218_),
    .X(_00609_));
 sky130_fd_sc_hd__nor2_2 _19982_ (.A(_10677_),
    .B(_05217_),
    .Y(_00610_));
 sky130_fd_sc_hd__nor2_2 _19983_ (.A(_10732_),
    .B(_05217_),
    .Y(_00611_));
 sky130_fd_sc_hd__nor2_2 _19984_ (.A(_10693_),
    .B(_05217_),
    .Y(_00612_));
 sky130_fd_sc_hd__nor2_2 _19985_ (.A(_10725_),
    .B(_05217_),
    .Y(_00613_));
 sky130_fd_sc_hd__buf_1 _19986_ (.A(_03588_),
    .X(_05219_));
 sky130_fd_sc_hd__nor2_2 _19987_ (.A(_10720_),
    .B(_05219_),
    .Y(_00614_));
 sky130_fd_sc_hd__and2_2 _19988_ (.A(_10854_),
    .B(_05214_),
    .X(_05220_));
 sky130_fd_sc_hd__buf_1 _19989_ (.A(_05220_),
    .X(_00615_));
 sky130_fd_sc_hd__nor2_2 _19990_ (.A(_10743_),
    .B(_05219_),
    .Y(_00616_));
 sky130_fd_sc_hd__and2_2 _19991_ (.A(_10697_),
    .B(_05214_),
    .X(_05221_));
 sky130_fd_sc_hd__buf_1 _19992_ (.A(_05221_),
    .X(_00617_));
 sky130_fd_sc_hd__nor2_2 _19993_ (.A(_10684_),
    .B(_05219_),
    .Y(_00618_));
 sky130_fd_sc_hd__nor2_2 _19994_ (.A(_10733_),
    .B(_05219_),
    .Y(_00619_));
 sky130_fd_sc_hd__buf_1 _19995_ (.A(\decode.id_ex_pcsel_reg ),
    .X(_05222_));
 sky130_fd_sc_hd__nor2_2 _19996_ (.A(\decode.id_ex_imm_reg[0] ),
    .B(\decode.id_ex_pc_reg[0] ),
    .Y(_05223_));
 sky130_fd_sc_hd__and2_2 _19997_ (.A(\decode.id_ex_imm_reg[0] ),
    .B(\decode.id_ex_pc_reg[0] ),
    .X(_05224_));
 sky130_fd_sc_hd__nor2_2 _19998_ (.A(_05223_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__nor2_2 _19999_ (.A(_05222_),
    .B(_03587_),
    .Y(_05226_));
 sky130_fd_sc_hd__buf_1 _20000_ (.A(_05226_),
    .X(_05227_));
 sky130_fd_sc_hd__o22a_2 _20001_ (.A1(_05222_),
    .A2(_05225_),
    .B1(_05227_),
    .B2(_00548_),
    .X(_00620_));
 sky130_fd_sc_hd__buf_1 _20002_ (.A(_05226_),
    .X(_05228_));
 sky130_fd_sc_hd__xnor2_2 _20003_ (.A(_04261_),
    .B(\decode.id_ex_pc_reg[1] ),
    .Y(_05229_));
 sky130_fd_sc_hd__xnor2_2 _20004_ (.A(_05224_),
    .B(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__buf_1 _20005_ (.A(_05222_),
    .X(_05231_));
 sky130_fd_sc_hd__o22a_2 _20006_ (.A1(_00549_),
    .A2(_05228_),
    .B1(_05230_),
    .B2(_05231_),
    .X(_00621_));
 sky130_fd_sc_hd__nor2_2 _20007_ (.A(_04018_),
    .B(_10711_),
    .Y(_05232_));
 sky130_fd_sc_hd__nor2_2 _20008_ (.A(\decode.id_ex_imm_reg[2] ),
    .B(_10834_),
    .Y(_05233_));
 sky130_fd_sc_hd__a22o_2 _20009_ (.A1(\decode.id_ex_imm_reg[0] ),
    .A2(\decode.id_ex_pc_reg[0] ),
    .B1(\decode.id_ex_pc_reg[1] ),
    .B2(\decode.id_ex_imm_reg[1] ),
    .X(_05234_));
 sky130_fd_sc_hd__o21a_2 _20010_ (.A1(_04261_),
    .A2(\decode.id_ex_pc_reg[1] ),
    .B1(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__o21ai_2 _20011_ (.A1(_05232_),
    .A2(_05233_),
    .B1(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__or3_2 _20012_ (.A(_05232_),
    .B(_05233_),
    .C(_05235_),
    .X(_05237_));
 sky130_fd_sc_hd__nand2_2 _20013_ (.A(_05236_),
    .B(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__buf_1 _20014_ (.A(_05222_),
    .X(_05239_));
 sky130_fd_sc_hd__o22a_2 _20015_ (.A1(_05238_),
    .A2(_05239_),
    .B1(_00550_),
    .B2(_05227_),
    .X(_00622_));
 sky130_fd_sc_hd__or2_2 _20016_ (.A(\decode.id_ex_imm_reg[3] ),
    .B(_10747_),
    .X(_05240_));
 sky130_fd_sc_hd__nand2_2 _20017_ (.A(\decode.id_ex_imm_reg[3] ),
    .B(\decode.id_ex_pc_reg[3] ),
    .Y(_05241_));
 sky130_fd_sc_hd__nand2_2 _20018_ (.A(_05240_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__o221ai_2 _20019_ (.A1(\decode.id_ex_imm_reg[1] ),
    .A2(\decode.id_ex_pc_reg[1] ),
    .B1(_10834_),
    .B2(\decode.id_ex_imm_reg[2] ),
    .C1(_05234_),
    .Y(_05243_));
 sky130_fd_sc_hd__o21a_2 _20020_ (.A1(_04018_),
    .A2(_10711_),
    .B1(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__xor2_2 _20021_ (.A(_05242_),
    .B(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__o22a_2 _20022_ (.A1(_05245_),
    .A2(_05239_),
    .B1(_00551_),
    .B2(_05227_),
    .X(_00623_));
 sky130_fd_sc_hd__buf_1 _20023_ (.A(_10758_),
    .X(_05246_));
 sky130_fd_sc_hd__or4_2 _20024_ (.A(_10575_),
    .B(_05222_),
    .C(_05246_),
    .D(_10908_),
    .X(_05247_));
 sky130_fd_sc_hd__nor2_2 _20025_ (.A(\decode.id_ex_imm_reg[4] ),
    .B(\decode.id_ex_pc_reg[4] ),
    .Y(_05248_));
 sky130_fd_sc_hd__nand2_2 _20026_ (.A(\decode.id_ex_imm_reg[4] ),
    .B(\decode.id_ex_pc_reg[4] ),
    .Y(_05249_));
 sky130_fd_sc_hd__and2b_2 _20027_ (.A_N(_05248_),
    .B(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__o211ai_2 _20028_ (.A1(_04018_),
    .A2(_10711_),
    .B1(_05241_),
    .C1(_05243_),
    .Y(_05251_));
 sky130_fd_sc_hd__o21ai_2 _20029_ (.A1(\decode.id_ex_imm_reg[3] ),
    .A2(_10747_),
    .B1(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__xor2_2 _20030_ (.A(_05250_),
    .B(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__o2bb2ai_2 _20031_ (.A1_N(_05231_),
    .A2_N(_00552_),
    .B1(_05247_),
    .B2(_05253_),
    .Y(_00624_));
 sky130_fd_sc_hd__or2_2 _20032_ (.A(\decode.id_ex_imm_reg[5] ),
    .B(_10704_),
    .X(_05254_));
 sky130_fd_sc_hd__nand2_2 _20033_ (.A(\decode.id_ex_imm_reg[5] ),
    .B(\decode.id_ex_pc_reg[5] ),
    .Y(_05255_));
 sky130_fd_sc_hd__o21ai_2 _20034_ (.A1(_05248_),
    .A2(_05252_),
    .B1(_05249_),
    .Y(_05256_));
 sky130_fd_sc_hd__a21oi_2 _20035_ (.A1(_05254_),
    .A2(_05255_),
    .B1(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__and3_2 _20036_ (.A(_05254_),
    .B(_05255_),
    .C(_05256_),
    .X(_05258_));
 sky130_fd_sc_hd__nor2_2 _20037_ (.A(_05257_),
    .B(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__o22a_2 _20038_ (.A1(_00553_),
    .A2(_05228_),
    .B1(_05259_),
    .B2(_05231_),
    .X(_00625_));
 sky130_fd_sc_hd__nor2_2 _20039_ (.A(\decode.id_ex_imm_reg[6] ),
    .B(_10678_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand2_2 _20040_ (.A(\decode.id_ex_imm_reg[6] ),
    .B(\decode.id_ex_pc_reg[6] ),
    .Y(_05261_));
 sky130_fd_sc_hd__and2b_2 _20041_ (.A_N(_05260_),
    .B(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__o211ai_2 _20042_ (.A1(\decode.id_ex_imm_reg[3] ),
    .A2(_10747_),
    .B1(_05250_),
    .C1(_05251_),
    .Y(_05263_));
 sky130_fd_sc_hd__nand3_2 _20043_ (.A(_05249_),
    .B(_05263_),
    .C(_05255_),
    .Y(_05264_));
 sky130_fd_sc_hd__o21ai_2 _20044_ (.A1(\decode.id_ex_imm_reg[5] ),
    .A2(_10704_),
    .B1(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__xor2_2 _20045_ (.A(_05262_),
    .B(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__inv_2 _20046_ (.A(_05222_),
    .Y(_05267_));
 sky130_fd_sc_hd__a2bb2oi_2 _20047_ (.A1_N(_00554_),
    .A2_N(_05227_),
    .B1(_05266_),
    .B2(_05267_),
    .Y(_00626_));
 sky130_fd_sc_hd__o211ai_2 _20048_ (.A1(\decode.id_ex_imm_reg[5] ),
    .A2(_10704_),
    .B1(_05262_),
    .C1(_05264_),
    .Y(_05268_));
 sky130_fd_sc_hd__nor2_2 _20049_ (.A(\decode.id_ex_imm_reg[7] ),
    .B(_10730_),
    .Y(_05269_));
 sky130_fd_sc_hd__and2_2 _20050_ (.A(\decode.id_ex_imm_reg[7] ),
    .B(\decode.id_ex_pc_reg[7] ),
    .X(_05270_));
 sky130_fd_sc_hd__nor2_2 _20051_ (.A(_05269_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__a21boi_2 _20052_ (.A1(_05261_),
    .A2(_05268_),
    .B1_N(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__o221a_2 _20053_ (.A1(_05269_),
    .A2(_05270_),
    .B1(_05260_),
    .B2(_05265_),
    .C1(_05261_),
    .X(_05273_));
 sky130_fd_sc_hd__nor2_2 _20054_ (.A(_05272_),
    .B(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__o22a_2 _20055_ (.A1(_00555_),
    .A2(_05228_),
    .B1(_05274_),
    .B2(_05231_),
    .X(_00627_));
 sky130_fd_sc_hd__a21oi_2 _20056_ (.A1(\decode.id_ex_imm_reg[7] ),
    .A2(_10730_),
    .B1(_05272_),
    .Y(_05275_));
 sky130_fd_sc_hd__xnor2_2 _20057_ (.A(\decode.id_ex_imm_reg[8] ),
    .B(\decode.id_ex_pc_reg[8] ),
    .Y(_05276_));
 sky130_fd_sc_hd__xor2_2 _20058_ (.A(_05275_),
    .B(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__o22a_2 _20059_ (.A1(_00556_),
    .A2(_05228_),
    .B1(_05277_),
    .B2(_05231_),
    .X(_00628_));
 sky130_fd_sc_hd__xor2_2 _20060_ (.A(\decode.id_ex_imm_reg[9] ),
    .B(_10706_),
    .X(_05278_));
 sky130_fd_sc_hd__o21bai_2 _20061_ (.A1(_05270_),
    .A2(_05272_),
    .B1_N(_05276_),
    .Y(_05279_));
 sky130_fd_sc_hd__a21bo_2 _20062_ (.A1(\decode.id_ex_imm_reg[8] ),
    .A2(\decode.id_ex_pc_reg[8] ),
    .B1_N(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__xor2_2 _20063_ (.A(_05278_),
    .B(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__o22a_2 _20064_ (.A1(_05281_),
    .A2(_05239_),
    .B1(_00557_),
    .B2(_05227_),
    .X(_00629_));
 sky130_fd_sc_hd__nor2_2 _20065_ (.A(\decode.id_ex_imm_reg[10] ),
    .B(\decode.id_ex_pc_reg[10] ),
    .Y(_05282_));
 sky130_fd_sc_hd__nand2_2 _20066_ (.A(\decode.id_ex_imm_reg[10] ),
    .B(\decode.id_ex_pc_reg[10] ),
    .Y(_05283_));
 sky130_fd_sc_hd__and2b_2 _20067_ (.A_N(_05282_),
    .B(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__a22oi_2 _20068_ (.A1(\decode.id_ex_imm_reg[8] ),
    .A2(\decode.id_ex_pc_reg[8] ),
    .B1(\decode.id_ex_pc_reg[9] ),
    .B2(\decode.id_ex_imm_reg[9] ),
    .Y(_05285_));
 sky130_fd_sc_hd__a2bb2o_2 _20069_ (.A1_N(\decode.id_ex_imm_reg[9] ),
    .A2_N(_10706_),
    .B1(_05285_),
    .B2(_05279_),
    .X(_05286_));
 sky130_fd_sc_hd__xnor2_2 _20070_ (.A(_05284_),
    .B(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__o22a_2 _20071_ (.A1(_00558_),
    .A2(_05228_),
    .B1(_05287_),
    .B2(_05231_),
    .X(_00630_));
 sky130_fd_sc_hd__and2_2 _20072_ (.A(\decode.id_ex_imm_reg[11] ),
    .B(_10689_),
    .X(_05288_));
 sky130_fd_sc_hd__nor2_2 _20073_ (.A(\decode.id_ex_imm_reg[11] ),
    .B(_10689_),
    .Y(_05289_));
 sky130_fd_sc_hd__o221ai_2 _20074_ (.A1(_05288_),
    .A2(_05289_),
    .B1(_05282_),
    .B2(_05286_),
    .C1(_05283_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand2_2 _20075_ (.A(_05279_),
    .B(_05285_),
    .Y(_05291_));
 sky130_fd_sc_hd__o211ai_2 _20076_ (.A1(\decode.id_ex_imm_reg[9] ),
    .A2(_10706_),
    .B1(_05284_),
    .C1(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__a211o_2 _20077_ (.A1(_05283_),
    .A2(_05292_),
    .B1(_05288_),
    .C1(_05289_),
    .X(_05293_));
 sky130_fd_sc_hd__and2_2 _20078_ (.A(_05290_),
    .B(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__o22a_2 _20079_ (.A1(_00559_),
    .A2(_05228_),
    .B1(_05294_),
    .B2(_05231_),
    .X(_00631_));
 sky130_fd_sc_hd__nor2_2 _20080_ (.A(\decode.id_ex_imm_reg[12] ),
    .B(\decode.id_ex_pc_reg[12] ),
    .Y(_05295_));
 sky130_fd_sc_hd__nand2_2 _20081_ (.A(\decode.id_ex_imm_reg[12] ),
    .B(\decode.id_ex_pc_reg[12] ),
    .Y(_05296_));
 sky130_fd_sc_hd__and2b_2 _20082_ (.A_N(_05295_),
    .B(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__nand2_2 _20083_ (.A(\decode.id_ex_imm_reg[11] ),
    .B(\decode.id_ex_pc_reg[11] ),
    .Y(_05298_));
 sky130_fd_sc_hd__a31o_2 _20084_ (.A1(_05283_),
    .A2(_05292_),
    .A3(_05298_),
    .B1(_05289_),
    .X(_05299_));
 sky130_fd_sc_hd__xor2_2 _20085_ (.A(_05297_),
    .B(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__a2bb2oi_2 _20086_ (.A1_N(_00560_),
    .A2_N(_05227_),
    .B1(_05300_),
    .B2(_05267_),
    .Y(_00632_));
 sky130_fd_sc_hd__and2_2 _20087_ (.A(\decode.id_ex_imm_reg[13] ),
    .B(_10710_),
    .X(_05301_));
 sky130_fd_sc_hd__nor2_2 _20088_ (.A(\decode.id_ex_imm_reg[13] ),
    .B(_10710_),
    .Y(_05302_));
 sky130_fd_sc_hd__o221ai_2 _20089_ (.A1(_05295_),
    .A2(_05299_),
    .B1(_05301_),
    .B2(_05302_),
    .C1(_05296_),
    .Y(_05303_));
 sky130_fd_sc_hd__nand3_2 _20090_ (.A(_05283_),
    .B(_05292_),
    .C(_05298_),
    .Y(_05304_));
 sky130_fd_sc_hd__o211ai_2 _20091_ (.A1(\decode.id_ex_imm_reg[11] ),
    .A2(_10689_),
    .B1(_05297_),
    .C1(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__a211o_2 _20092_ (.A1(_05296_),
    .A2(_05305_),
    .B1(_05301_),
    .C1(_05302_),
    .X(_05306_));
 sky130_fd_sc_hd__and2_2 _20093_ (.A(_05303_),
    .B(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__o22a_2 _20094_ (.A1(_00561_),
    .A2(_05228_),
    .B1(_05307_),
    .B2(_05231_),
    .X(_00633_));
 sky130_fd_sc_hd__nor2_2 _20095_ (.A(\decode.id_ex_imm_reg[14] ),
    .B(\decode.id_ex_pc_reg[14] ),
    .Y(_05308_));
 sky130_fd_sc_hd__nand2_2 _20096_ (.A(\decode.id_ex_imm_reg[14] ),
    .B(\decode.id_ex_pc_reg[14] ),
    .Y(_05309_));
 sky130_fd_sc_hd__and2b_2 _20097_ (.A_N(_05308_),
    .B(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__nand2_2 _20098_ (.A(\decode.id_ex_imm_reg[13] ),
    .B(\decode.id_ex_pc_reg[13] ),
    .Y(_05311_));
 sky130_fd_sc_hd__a31o_2 _20099_ (.A1(_05296_),
    .A2(_05305_),
    .A3(_05311_),
    .B1(_05302_),
    .X(_05312_));
 sky130_fd_sc_hd__xnor2_2 _20100_ (.A(_05310_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__o22a_2 _20101_ (.A1(_00562_),
    .A2(_05228_),
    .B1(_05313_),
    .B2(_05231_),
    .X(_00634_));
 sky130_fd_sc_hd__nand2_2 _20102_ (.A(\decode.id_ex_imm_reg[15] ),
    .B(_10681_),
    .Y(_05314_));
 sky130_fd_sc_hd__or2_2 _20103_ (.A(\decode.id_ex_imm_reg[15] ),
    .B(_10681_),
    .X(_05315_));
 sky130_fd_sc_hd__nand2_2 _20104_ (.A(_05314_),
    .B(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__o21ai_2 _20105_ (.A1(_05308_),
    .A2(_05312_),
    .B1(_05309_),
    .Y(_05317_));
 sky130_fd_sc_hd__xor2_2 _20106_ (.A(_05316_),
    .B(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__a2bb2oi_2 _20107_ (.A1_N(_00563_),
    .A2_N(_05227_),
    .B1(_05318_),
    .B2(_05267_),
    .Y(_00635_));
 sky130_fd_sc_hd__nor2_2 _20108_ (.A(\decode.id_ex_imm_reg[16] ),
    .B(\decode.id_ex_pc_reg[16] ),
    .Y(_05319_));
 sky130_fd_sc_hd__nand2_2 _20109_ (.A(\decode.id_ex_imm_reg[16] ),
    .B(\decode.id_ex_pc_reg[16] ),
    .Y(_05320_));
 sky130_fd_sc_hd__and2b_2 _20110_ (.A_N(_05319_),
    .B(_05320_),
    .X(_05321_));
 sky130_fd_sc_hd__nand3_2 _20111_ (.A(_05296_),
    .B(_05305_),
    .C(_05311_),
    .Y(_05322_));
 sky130_fd_sc_hd__o211ai_2 _20112_ (.A1(\decode.id_ex_imm_reg[13] ),
    .A2(_10710_),
    .B1(_05310_),
    .C1(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__nand3_2 _20113_ (.A(_05309_),
    .B(_05323_),
    .C(_05314_),
    .Y(_05324_));
 sky130_fd_sc_hd__o21ai_2 _20114_ (.A1(\decode.id_ex_imm_reg[15] ),
    .A2(_10681_),
    .B1(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__xnor2_2 _20115_ (.A(_05321_),
    .B(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__o22a_2 _20116_ (.A1(_00564_),
    .A2(_05226_),
    .B1(_05326_),
    .B2(_05231_),
    .X(_00636_));
 sky130_fd_sc_hd__nand2_2 _20117_ (.A(\decode.id_ex_imm_reg[17] ),
    .B(_10806_),
    .Y(_05327_));
 sky130_fd_sc_hd__or2_2 _20118_ (.A(\decode.id_ex_imm_reg[17] ),
    .B(_10806_),
    .X(_05328_));
 sky130_fd_sc_hd__and2_2 _20119_ (.A(_05327_),
    .B(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__o21ai_2 _20120_ (.A1(_05319_),
    .A2(_05325_),
    .B1(_05320_),
    .Y(_05330_));
 sky130_fd_sc_hd__xor2_2 _20121_ (.A(_05329_),
    .B(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__o22a_2 _20122_ (.A1(_00565_),
    .A2(_05226_),
    .B1(_05331_),
    .B2(_05239_),
    .X(_00637_));
 sky130_fd_sc_hd__nor2_2 _20123_ (.A(\decode.id_ex_imm_reg[18] ),
    .B(\decode.id_ex_pc_reg[18] ),
    .Y(_05332_));
 sky130_fd_sc_hd__nand2_2 _20124_ (.A(\decode.id_ex_imm_reg[18] ),
    .B(\decode.id_ex_pc_reg[18] ),
    .Y(_05333_));
 sky130_fd_sc_hd__and2b_2 _20125_ (.A_N(_05332_),
    .B(_05333_),
    .X(_05334_));
 sky130_fd_sc_hd__o211ai_2 _20126_ (.A1(\decode.id_ex_imm_reg[15] ),
    .A2(_10681_),
    .B1(_05321_),
    .C1(_05324_),
    .Y(_05335_));
 sky130_fd_sc_hd__nand3_2 _20127_ (.A(_05320_),
    .B(_05335_),
    .C(_05327_),
    .Y(_05336_));
 sky130_fd_sc_hd__o21ai_2 _20128_ (.A1(\decode.id_ex_imm_reg[17] ),
    .A2(_10806_),
    .B1(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__xnor2_2 _20129_ (.A(_05334_),
    .B(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__o22a_2 _20130_ (.A1(_00566_),
    .A2(_05226_),
    .B1(_05338_),
    .B2(_05239_),
    .X(_00638_));
 sky130_fd_sc_hd__nand2_2 _20131_ (.A(\decode.id_ex_imm_reg[19] ),
    .B(\decode.id_ex_pc_reg[19] ),
    .Y(_05339_));
 sky130_fd_sc_hd__buf_1 _20132_ (.A(\decode.id_ex_pc_reg[19] ),
    .X(_05340_));
 sky130_fd_sc_hd__or2_2 _20133_ (.A(\decode.id_ex_imm_reg[19] ),
    .B(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__nand2_2 _20134_ (.A(_05339_),
    .B(_05341_),
    .Y(_05342_));
 sky130_fd_sc_hd__o21ai_2 _20135_ (.A1(_05332_),
    .A2(_05337_),
    .B1(_05333_),
    .Y(_05343_));
 sky130_fd_sc_hd__xor2_2 _20136_ (.A(_05342_),
    .B(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__a2bb2oi_2 _20137_ (.A1_N(_00567_),
    .A2_N(_05227_),
    .B1(_05344_),
    .B2(_05267_),
    .Y(_00639_));
 sky130_fd_sc_hd__xor2_2 _20138_ (.A(\decode.id_ex_imm_reg[20] ),
    .B(_10867_),
    .X(_05345_));
 sky130_fd_sc_hd__o211ai_2 _20139_ (.A1(\decode.id_ex_imm_reg[17] ),
    .A2(_10806_),
    .B1(_05334_),
    .C1(_05336_),
    .Y(_05346_));
 sky130_fd_sc_hd__nand3_2 _20140_ (.A(_05333_),
    .B(_05346_),
    .C(_05339_),
    .Y(_05347_));
 sky130_fd_sc_hd__o21ai_2 _20141_ (.A1(\decode.id_ex_imm_reg[19] ),
    .A2(_05340_),
    .B1(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__xnor2_2 _20142_ (.A(_05345_),
    .B(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__o22a_2 _20143_ (.A1(_00568_),
    .A2(_05226_),
    .B1(_05349_),
    .B2(_05239_),
    .X(_00640_));
 sky130_fd_sc_hd__or2_2 _20144_ (.A(\decode.id_ex_imm_reg[21] ),
    .B(_10798_),
    .X(_05350_));
 sky130_fd_sc_hd__nand2_2 _20145_ (.A(\decode.id_ex_imm_reg[21] ),
    .B(_10798_),
    .Y(_05351_));
 sky130_fd_sc_hd__nand2_2 _20146_ (.A(_05350_),
    .B(_05351_),
    .Y(_05352_));
 sky130_fd_sc_hd__and3_2 _20147_ (.A(_05341_),
    .B(_05347_),
    .C(_05345_),
    .X(_05353_));
 sky130_fd_sc_hd__a21o_2 _20148_ (.A1(\decode.id_ex_imm_reg[20] ),
    .A2(_10867_),
    .B1(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__xnor2_2 _20149_ (.A(_05352_),
    .B(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__o22a_2 _20150_ (.A1(_05222_),
    .A2(_05355_),
    .B1(_05228_),
    .B2(_00569_),
    .X(_00641_));
 sky130_fd_sc_hd__a221o_2 _20151_ (.A1(\decode.id_ex_imm_reg[20] ),
    .A2(_10867_),
    .B1(_10798_),
    .B2(\decode.id_ex_imm_reg[21] ),
    .C1(_05353_),
    .X(_05356_));
 sky130_fd_sc_hd__xor2_2 _20152_ (.A(\decode.id_ex_imm_reg[22] ),
    .B(_10864_),
    .X(_05357_));
 sky130_fd_sc_hd__a21o_2 _20153_ (.A1(_05350_),
    .A2(_05356_),
    .B1(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__o211ai_2 _20154_ (.A1(\decode.id_ex_imm_reg[19] ),
    .A2(_05340_),
    .B1(_05345_),
    .C1(_05347_),
    .Y(_05359_));
 sky130_fd_sc_hd__a22oi_2 _20155_ (.A1(\decode.id_ex_imm_reg[20] ),
    .A2(_10867_),
    .B1(_10798_),
    .B2(\decode.id_ex_imm_reg[21] ),
    .Y(_05360_));
 sky130_fd_sc_hd__o21ai_2 _20156_ (.A1(\decode.id_ex_imm_reg[21] ),
    .A2(_10798_),
    .B1(_05357_),
    .Y(_05361_));
 sky130_fd_sc_hd__a21o_2 _20157_ (.A1(_05359_),
    .A2(_05360_),
    .B1(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__and2_2 _20158_ (.A(_05358_),
    .B(_05362_),
    .X(_05363_));
 sky130_fd_sc_hd__o22a_2 _20159_ (.A1(_00570_),
    .A2(_05226_),
    .B1(_05363_),
    .B2(_05239_),
    .X(_00642_));
 sky130_fd_sc_hd__xor2_2 _20160_ (.A(\decode.id_ex_imm_reg[23] ),
    .B(_10786_),
    .X(_05364_));
 sky130_fd_sc_hd__a21oi_2 _20161_ (.A1(_05359_),
    .A2(_05360_),
    .B1(_05361_),
    .Y(_05365_));
 sky130_fd_sc_hd__a21o_2 _20162_ (.A1(\decode.id_ex_imm_reg[22] ),
    .A2(_10864_),
    .B1(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__xor2_2 _20163_ (.A(_05364_),
    .B(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__o22a_2 _20164_ (.A1(_05222_),
    .A2(_05367_),
    .B1(_05228_),
    .B2(_00571_),
    .X(_00643_));
 sky130_fd_sc_hd__nor2_2 _20165_ (.A(\decode.id_ex_imm_reg[24] ),
    .B(\decode.id_ex_pc_reg[24] ),
    .Y(_05368_));
 sky130_fd_sc_hd__nand2_2 _20166_ (.A(\decode.id_ex_imm_reg[24] ),
    .B(\decode.id_ex_pc_reg[24] ),
    .Y(_05369_));
 sky130_fd_sc_hd__and2b_2 _20167_ (.A_N(_05368_),
    .B(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__a22o_2 _20168_ (.A1(\decode.id_ex_imm_reg[22] ),
    .A2(_10864_),
    .B1(_10786_),
    .B2(\decode.id_ex_imm_reg[23] ),
    .X(_05371_));
 sky130_fd_sc_hd__o22ai_2 _20169_ (.A1(\decode.id_ex_imm_reg[23] ),
    .A2(_10786_),
    .B1(_05371_),
    .B2(_05365_),
    .Y(_05372_));
 sky130_fd_sc_hd__xnor2_2 _20170_ (.A(_05370_),
    .B(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__o22a_2 _20171_ (.A1(_00572_),
    .A2(_05226_),
    .B1(_05373_),
    .B2(_05239_),
    .X(_00644_));
 sky130_fd_sc_hd__or2_2 _20172_ (.A(\decode.id_ex_imm_reg[25] ),
    .B(_10790_),
    .X(_05374_));
 sky130_fd_sc_hd__nand2_2 _20173_ (.A(\decode.id_ex_imm_reg[25] ),
    .B(_10790_),
    .Y(_05375_));
 sky130_fd_sc_hd__nand2_2 _20174_ (.A(_05374_),
    .B(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__o21a_2 _20175_ (.A1(_05368_),
    .A2(_05372_),
    .B1(_05369_),
    .X(_05377_));
 sky130_fd_sc_hd__xnor2_2 _20176_ (.A(_05376_),
    .B(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__a22oi_2 _20177_ (.A1(_05068_),
    .A2(_05247_),
    .B1(_05378_),
    .B2(_05267_),
    .Y(_00645_));
 sky130_fd_sc_hd__o221ai_2 _20178_ (.A1(\decode.id_ex_imm_reg[23] ),
    .A2(_10786_),
    .B1(_05371_),
    .B2(_05365_),
    .C1(_05370_),
    .Y(_05379_));
 sky130_fd_sc_hd__nand3_2 _20179_ (.A(_05369_),
    .B(_05379_),
    .C(_05375_),
    .Y(_05380_));
 sky130_fd_sc_hd__xor2_2 _20180_ (.A(\decode.id_ex_imm_reg[26] ),
    .B(\decode.id_ex_pc_reg[26] ),
    .X(_05381_));
 sky130_fd_sc_hd__a21oi_2 _20181_ (.A1(_05374_),
    .A2(_05380_),
    .B1(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__o211ai_2 _20182_ (.A1(\decode.id_ex_imm_reg[25] ),
    .A2(_10790_),
    .B1(_05381_),
    .C1(_05380_),
    .Y(_05383_));
 sky130_fd_sc_hd__and2b_2 _20183_ (.A_N(_05382_),
    .B(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__o22a_2 _20184_ (.A1(_00574_),
    .A2(_05226_),
    .B1(_05384_),
    .B2(_05239_),
    .X(_00646_));
 sky130_fd_sc_hd__or2_2 _20185_ (.A(\decode.id_ex_imm_reg[27] ),
    .B(_10854_),
    .X(_05385_));
 sky130_fd_sc_hd__nand2_2 _20186_ (.A(\decode.id_ex_imm_reg[27] ),
    .B(_10854_),
    .Y(_05386_));
 sky130_fd_sc_hd__nand2_2 _20187_ (.A(_05385_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__a32o_2 _20188_ (.A1(_05374_),
    .A2(_05380_),
    .A3(_05381_),
    .B1(\decode.id_ex_pc_reg[26] ),
    .B2(\decode.id_ex_imm_reg[26] ),
    .X(_05388_));
 sky130_fd_sc_hd__xor2_2 _20189_ (.A(_05387_),
    .B(_05388_),
    .X(_05389_));
 sky130_fd_sc_hd__inv_2 _20190_ (.A(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__o22a_2 _20191_ (.A1(_00575_),
    .A2(_05226_),
    .B1(_05390_),
    .B2(_05239_),
    .X(_00647_));
 sky130_fd_sc_hd__nand2_2 _20192_ (.A(\decode.id_ex_imm_reg[26] ),
    .B(\decode.id_ex_pc_reg[26] ),
    .Y(_05391_));
 sky130_fd_sc_hd__nand3_2 _20193_ (.A(_05391_),
    .B(_05383_),
    .C(_05386_),
    .Y(_05392_));
 sky130_fd_sc_hd__and2_2 _20194_ (.A(\decode.id_ex_imm_reg[28] ),
    .B(\decode.id_ex_pc_reg[28] ),
    .X(_05393_));
 sky130_fd_sc_hd__nor2_2 _20195_ (.A(\decode.id_ex_imm_reg[28] ),
    .B(\decode.id_ex_pc_reg[28] ),
    .Y(_05394_));
 sky130_fd_sc_hd__nor2_2 _20196_ (.A(_05393_),
    .B(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__a21oi_2 _20197_ (.A1(_05385_),
    .A2(_05392_),
    .B1(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__o211ai_2 _20198_ (.A1(\decode.id_ex_imm_reg[27] ),
    .A2(_10854_),
    .B1(_05395_),
    .C1(_05392_),
    .Y(_05397_));
 sky130_fd_sc_hd__or2b_2 _20199_ (.A(_05396_),
    .B_N(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__a2bb2oi_2 _20200_ (.A1_N(_00576_),
    .A2_N(_05227_),
    .B1(_05398_),
    .B2(_05267_),
    .Y(_00648_));
 sky130_fd_sc_hd__nor2_2 _20201_ (.A(\decode.id_ex_imm_reg[29] ),
    .B(_10697_),
    .Y(_05399_));
 sky130_fd_sc_hd__and2_2 _20202_ (.A(\decode.id_ex_imm_reg[29] ),
    .B(_10697_),
    .X(_05400_));
 sky130_fd_sc_hd__nor2_2 _20203_ (.A(_05399_),
    .B(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__a31oi_2 _20204_ (.A1(_05385_),
    .A2(_05392_),
    .A3(_05395_),
    .B1(_05393_),
    .Y(_05402_));
 sky130_fd_sc_hd__xor2_2 _20205_ (.A(_05401_),
    .B(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__a2bb2oi_2 _20206_ (.A1_N(_00577_),
    .A2_N(_05227_),
    .B1(_05403_),
    .B2(_05267_),
    .Y(_00649_));
 sky130_fd_sc_hd__o21bai_2 _20207_ (.A1(_05399_),
    .A2(_05402_),
    .B1_N(_05400_),
    .Y(_05404_));
 sky130_fd_sc_hd__xor2_2 _20208_ (.A(\decode.id_ex_imm_reg[30] ),
    .B(\decode.id_ex_pc_reg[30] ),
    .X(_05405_));
 sky130_fd_sc_hd__xnor2_2 _20209_ (.A(_05404_),
    .B(_05405_),
    .Y(_05406_));
 sky130_fd_sc_hd__a22oi_2 _20210_ (.A1(_05178_),
    .A2(_05247_),
    .B1(_05406_),
    .B2(_05267_),
    .Y(_00650_));
 sky130_fd_sc_hd__nand2_2 _20211_ (.A(\decode.id_ex_imm_reg[30] ),
    .B(\decode.id_ex_pc_reg[30] ),
    .Y(_05407_));
 sky130_fd_sc_hd__a21bo_2 _20212_ (.A1(_05404_),
    .A2(_05405_),
    .B1_N(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__xor2_2 _20213_ (.A(\decode.id_ex_imm_reg[31] ),
    .B(\decode.id_ex_pc_reg[31] ),
    .X(_05409_));
 sky130_fd_sc_hd__xnor2_2 _20214_ (.A(_05408_),
    .B(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__a22oi_2 _20215_ (.A1(_05410_),
    .A2(_05267_),
    .B1(_05200_),
    .B2(_05247_),
    .Y(_00651_));
 sky130_fd_sc_hd__buf_1 _20216_ (.A(\decode.id_ex_rdsel_reg ),
    .X(_05411_));
 sky130_fd_sc_hd__buf_1 _20217_ (.A(_05411_),
    .X(_05412_));
 sky130_fd_sc_hd__o21ai_2 _20218_ (.A1(_05223_),
    .A2(_05224_),
    .B1(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__buf_1 _20219_ (.A(_04459_),
    .X(_05414_));
 sky130_fd_sc_hd__o211a_2 _20220_ (.A1(\decode.id_ex_pc_reg[0] ),
    .A2(_05412_),
    .B1(_05413_),
    .C1(_05414_),
    .X(_00652_));
 sky130_fd_sc_hd__inv_2 _20221_ (.A(\decode.id_ex_rdsel_reg ),
    .Y(_05415_));
 sky130_fd_sc_hd__buf_1 _20222_ (.A(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__buf_1 _20223_ (.A(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__buf_1 _20224_ (.A(\decode.id_ex_rdsel_reg ),
    .X(_05418_));
 sky130_fd_sc_hd__or2_2 _20225_ (.A(\decode.id_ex_pc_reg[1] ),
    .B(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__o211a_2 _20226_ (.A1(_05417_),
    .A2(_05230_),
    .B1(_05419_),
    .C1(_05414_),
    .X(_00653_));
 sky130_fd_sc_hd__buf_1 _20227_ (.A(_05416_),
    .X(_05420_));
 sky130_fd_sc_hd__nand2_2 _20228_ (.A(_05420_),
    .B(_10834_),
    .Y(_05421_));
 sky130_fd_sc_hd__o211a_2 _20229_ (.A1(_05417_),
    .A2(_05238_),
    .B1(_05421_),
    .C1(_05414_),
    .X(_00654_));
 sky130_fd_sc_hd__nand2_2 _20230_ (.A(_10834_),
    .B(_10747_),
    .Y(_05422_));
 sky130_fd_sc_hd__o21a_2 _20231_ (.A1(_10834_),
    .A2(_10747_),
    .B1(_05415_),
    .X(_05423_));
 sky130_fd_sc_hd__a22o_2 _20232_ (.A1(_05422_),
    .A2(_05423_),
    .B1(_05245_),
    .B2(_05411_),
    .X(_05424_));
 sky130_fd_sc_hd__buf_1 _20233_ (.A(_03582_),
    .X(_05425_));
 sky130_fd_sc_hd__and3b_2 _20234_ (.A_N(_03581_),
    .B(_05424_),
    .C(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__buf_1 _20235_ (.A(_05426_),
    .X(_00655_));
 sky130_fd_sc_hd__and3_2 _20236_ (.A(_10834_),
    .B(_10747_),
    .C(\decode.id_ex_pc_reg[4] ),
    .X(_05427_));
 sky130_fd_sc_hd__a21oi_2 _20237_ (.A1(_10834_),
    .A2(_10747_),
    .B1(\decode.id_ex_pc_reg[4] ),
    .Y(_05428_));
 sky130_fd_sc_hd__o21a_2 _20238_ (.A1(_05427_),
    .A2(_05428_),
    .B1(_05415_),
    .X(_05429_));
 sky130_fd_sc_hd__a2111oi_2 _20239_ (.A1(_05412_),
    .A2(_05253_),
    .B1(_05429_),
    .C1(_03517_),
    .D1(_03551_),
    .Y(_00656_));
 sky130_fd_sc_hd__and4_2 _20240_ (.A(_10834_),
    .B(_10747_),
    .C(\decode.id_ex_pc_reg[4] ),
    .D(_10704_),
    .X(_05430_));
 sky130_fd_sc_hd__o21ai_2 _20241_ (.A1(_10704_),
    .A2(_05427_),
    .B1(_05416_),
    .Y(_05431_));
 sky130_fd_sc_hd__o2bb2a_2 _20242_ (.A1_N(_05418_),
    .A2_N(_05259_),
    .B1(_05430_),
    .B2(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__nor2_2 _20243_ (.A(_05432_),
    .B(_05219_),
    .Y(_00657_));
 sky130_fd_sc_hd__and3_2 _20244_ (.A(_10704_),
    .B(_10678_),
    .C(_05427_),
    .X(_05433_));
 sky130_fd_sc_hd__a21oi_2 _20245_ (.A1(_10704_),
    .A2(_05427_),
    .B1(_10678_),
    .Y(_05434_));
 sky130_fd_sc_hd__o21a_2 _20246_ (.A1(_05433_),
    .A2(_05434_),
    .B1(_05415_),
    .X(_05435_));
 sky130_fd_sc_hd__a2111oi_2 _20247_ (.A1(_05412_),
    .A2(_05266_),
    .B1(_05435_),
    .C1(_03517_),
    .D1(_03551_),
    .Y(_00658_));
 sky130_fd_sc_hd__a31o_2 _20248_ (.A1(_10704_),
    .A2(_10678_),
    .A3(_05427_),
    .B1(_10730_),
    .X(_05436_));
 sky130_fd_sc_hd__nand2_2 _20249_ (.A(_10730_),
    .B(_05433_),
    .Y(_05437_));
 sky130_fd_sc_hd__a21o_2 _20250_ (.A1(_05436_),
    .A2(_05437_),
    .B1(_05418_),
    .X(_05438_));
 sky130_fd_sc_hd__o211a_2 _20251_ (.A1(_05417_),
    .A2(_05274_),
    .B1(_05438_),
    .C1(_05414_),
    .X(_00659_));
 sky130_fd_sc_hd__buf_1 _20252_ (.A(_10910_),
    .X(_05439_));
 sky130_fd_sc_hd__and3_2 _20253_ (.A(_10730_),
    .B(\decode.id_ex_pc_reg[8] ),
    .C(_05433_),
    .X(_05440_));
 sky130_fd_sc_hd__nor2_2 _20254_ (.A(\decode.id_ex_rdsel_reg ),
    .B(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__a31o_2 _20255_ (.A1(_10678_),
    .A2(_10730_),
    .A3(_05430_),
    .B1(\decode.id_ex_pc_reg[8] ),
    .X(_05442_));
 sky130_fd_sc_hd__a22o_2 _20256_ (.A1(_05441_),
    .A2(_05442_),
    .B1(_05277_),
    .B2(_05411_),
    .X(_05443_));
 sky130_fd_sc_hd__and3b_2 _20257_ (.A_N(_05439_),
    .B(_05443_),
    .C(_05425_),
    .X(_05444_));
 sky130_fd_sc_hd__buf_1 _20258_ (.A(_05444_),
    .X(_00660_));
 sky130_fd_sc_hd__a31o_2 _20259_ (.A1(_10730_),
    .A2(\decode.id_ex_pc_reg[8] ),
    .A3(_05433_),
    .B1(_10706_),
    .X(_05445_));
 sky130_fd_sc_hd__or4b_2 _20260_ (.A(_10731_),
    .B(_10680_),
    .C(_10707_),
    .D_N(_05433_),
    .X(_05446_));
 sky130_fd_sc_hd__a21o_2 _20261_ (.A1(_05445_),
    .A2(_05446_),
    .B1(_05418_),
    .X(_05447_));
 sky130_fd_sc_hd__o211a_2 _20262_ (.A1(_05417_),
    .A2(_05281_),
    .B1(_05447_),
    .C1(_05414_),
    .X(_00661_));
 sky130_fd_sc_hd__a21oi_2 _20263_ (.A1(_10706_),
    .A2(_05440_),
    .B1(\decode.id_ex_pc_reg[10] ),
    .Y(_05448_));
 sky130_fd_sc_hd__and3_2 _20264_ (.A(_10706_),
    .B(\decode.id_ex_pc_reg[10] ),
    .C(_05440_),
    .X(_05449_));
 sky130_fd_sc_hd__o21ai_2 _20265_ (.A1(_05448_),
    .A2(_05449_),
    .B1(_05420_),
    .Y(_05450_));
 sky130_fd_sc_hd__o211a_2 _20266_ (.A1(_05417_),
    .A2(_05287_),
    .B1(_05450_),
    .C1(_05414_),
    .X(_00662_));
 sky130_fd_sc_hd__nor2_2 _20267_ (.A(_10689_),
    .B(_05449_),
    .Y(_05451_));
 sky130_fd_sc_hd__and4_2 _20268_ (.A(_10706_),
    .B(\decode.id_ex_pc_reg[10] ),
    .C(_10689_),
    .D(_05440_),
    .X(_05452_));
 sky130_fd_sc_hd__o21ai_2 _20269_ (.A1(_05451_),
    .A2(_05452_),
    .B1(_05420_),
    .Y(_05453_));
 sky130_fd_sc_hd__buf_1 _20270_ (.A(_05214_),
    .X(_05454_));
 sky130_fd_sc_hd__o211a_2 _20271_ (.A1(_05417_),
    .A2(_05294_),
    .B1(_05453_),
    .C1(_05454_),
    .X(_00663_));
 sky130_fd_sc_hd__a41o_2 _20272_ (.A1(_10706_),
    .A2(\decode.id_ex_pc_reg[10] ),
    .A3(_10689_),
    .A4(_05440_),
    .B1(_10694_),
    .X(_05455_));
 sky130_fd_sc_hd__nand2_2 _20273_ (.A(_10694_),
    .B(_05452_),
    .Y(_05456_));
 sky130_fd_sc_hd__a21oi_2 _20274_ (.A1(_05455_),
    .A2(_05456_),
    .B1(_05411_),
    .Y(_05457_));
 sky130_fd_sc_hd__a2111oi_2 _20275_ (.A1(_05412_),
    .A2(_05300_),
    .B1(_05457_),
    .C1(_03517_),
    .D1(_03551_),
    .Y(_00664_));
 sky130_fd_sc_hd__and3_2 _20276_ (.A(_10694_),
    .B(_10710_),
    .C(_05452_),
    .X(_05458_));
 sky130_fd_sc_hd__a21oi_2 _20277_ (.A1(_10694_),
    .A2(_05452_),
    .B1(_10710_),
    .Y(_05459_));
 sky130_fd_sc_hd__o21ai_2 _20278_ (.A1(_05458_),
    .A2(_05459_),
    .B1(_05420_),
    .Y(_05460_));
 sky130_fd_sc_hd__o211a_2 _20279_ (.A1(_05417_),
    .A2(_05307_),
    .B1(_05460_),
    .C1(_05454_),
    .X(_00665_));
 sky130_fd_sc_hd__nor2_2 _20280_ (.A(\decode.id_ex_pc_reg[14] ),
    .B(_05458_),
    .Y(_05461_));
 sky130_fd_sc_hd__and4_2 _20281_ (.A(_10694_),
    .B(_10710_),
    .C(\decode.id_ex_pc_reg[14] ),
    .D(_05452_),
    .X(_05462_));
 sky130_fd_sc_hd__o21ai_2 _20282_ (.A1(_05461_),
    .A2(_05462_),
    .B1(_05420_),
    .Y(_05463_));
 sky130_fd_sc_hd__o211a_2 _20283_ (.A1(_05417_),
    .A2(_05313_),
    .B1(_05463_),
    .C1(_05454_),
    .X(_00666_));
 sky130_fd_sc_hd__or3b_2 _20284_ (.A(_10702_),
    .B(_10682_),
    .C_N(_05458_),
    .X(_05464_));
 sky130_fd_sc_hd__a41o_2 _20285_ (.A1(_10694_),
    .A2(_10710_),
    .A3(\decode.id_ex_pc_reg[14] ),
    .A4(_05452_),
    .B1(_10681_),
    .X(_05465_));
 sky130_fd_sc_hd__a21oi_2 _20286_ (.A1(_05464_),
    .A2(_05465_),
    .B1(_05411_),
    .Y(_05466_));
 sky130_fd_sc_hd__a2111oi_2 _20287_ (.A1(_05412_),
    .A2(_05318_),
    .B1(_05466_),
    .C1(_03517_),
    .D1(_03551_),
    .Y(_00667_));
 sky130_fd_sc_hd__a21oi_2 _20288_ (.A1(_10681_),
    .A2(_05462_),
    .B1(\decode.id_ex_pc_reg[16] ),
    .Y(_05467_));
 sky130_fd_sc_hd__and3_2 _20289_ (.A(_10681_),
    .B(\decode.id_ex_pc_reg[16] ),
    .C(_05462_),
    .X(_05468_));
 sky130_fd_sc_hd__o21ai_2 _20290_ (.A1(_05467_),
    .A2(_05468_),
    .B1(_05420_),
    .Y(_05469_));
 sky130_fd_sc_hd__o211a_2 _20291_ (.A1(_05417_),
    .A2(_05326_),
    .B1(_05469_),
    .C1(_05454_),
    .X(_00668_));
 sky130_fd_sc_hd__and4_2 _20292_ (.A(_10681_),
    .B(\decode.id_ex_pc_reg[16] ),
    .C(_10806_),
    .D(_05462_),
    .X(_05470_));
 sky130_fd_sc_hd__o21ai_2 _20293_ (.A1(_10806_),
    .A2(_05468_),
    .B1(_05416_),
    .Y(_05471_));
 sky130_fd_sc_hd__o2bb2a_2 _20294_ (.A1_N(_05418_),
    .A2_N(_05331_),
    .B1(_05470_),
    .B2(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__nor2_2 _20295_ (.A(_05472_),
    .B(_05219_),
    .Y(_00669_));
 sky130_fd_sc_hd__and3_2 _20296_ (.A(_10806_),
    .B(\decode.id_ex_pc_reg[18] ),
    .C(_05468_),
    .X(_05473_));
 sky130_fd_sc_hd__o21ai_2 _20297_ (.A1(\decode.id_ex_pc_reg[18] ),
    .A2(_05470_),
    .B1(_05416_),
    .Y(_05474_));
 sky130_fd_sc_hd__o2bb2a_2 _20298_ (.A1_N(_05418_),
    .A2_N(_05338_),
    .B1(_05473_),
    .B2(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__nor2_2 _20299_ (.A(_05475_),
    .B(_05219_),
    .Y(_00670_));
 sky130_fd_sc_hd__a31o_2 _20300_ (.A1(_10806_),
    .A2(\decode.id_ex_pc_reg[18] ),
    .A3(_05468_),
    .B1(_05340_),
    .X(_05476_));
 sky130_fd_sc_hd__a21oi_2 _20301_ (.A1(_05340_),
    .A2(_05473_),
    .B1(_05411_),
    .Y(_05477_));
 sky130_fd_sc_hd__o2bb2a_2 _20302_ (.A1_N(_05476_),
    .A2_N(_05477_),
    .B1(_05416_),
    .B2(_05344_),
    .X(_05478_));
 sky130_fd_sc_hd__nor2_2 _20303_ (.A(_05478_),
    .B(_05219_),
    .Y(_00671_));
 sky130_fd_sc_hd__a21oi_2 _20304_ (.A1(_05340_),
    .A2(_05473_),
    .B1(_10867_),
    .Y(_05479_));
 sky130_fd_sc_hd__a31o_2 _20305_ (.A1(_05340_),
    .A2(_10867_),
    .A3(_05473_),
    .B1(\decode.id_ex_rdsel_reg ),
    .X(_05480_));
 sky130_fd_sc_hd__o2bb2a_2 _20306_ (.A1_N(_05411_),
    .A2_N(_05349_),
    .B1(_05479_),
    .B2(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__nor2_2 _20307_ (.A(_05481_),
    .B(_05219_),
    .Y(_00672_));
 sky130_fd_sc_hd__and4_2 _20308_ (.A(_05340_),
    .B(_10867_),
    .C(_10798_),
    .D(_05473_),
    .X(_05482_));
 sky130_fd_sc_hd__a31o_2 _20309_ (.A1(_05340_),
    .A2(_10867_),
    .A3(_05473_),
    .B1(_10798_),
    .X(_05483_));
 sky130_fd_sc_hd__or3b_2 _20310_ (.A(_05411_),
    .B(_05482_),
    .C_N(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__nand2_2 _20311_ (.A(_05355_),
    .B(_05412_),
    .Y(_05485_));
 sky130_fd_sc_hd__a21oi_2 _20312_ (.A1(_05484_),
    .A2(_05485_),
    .B1(_03588_),
    .Y(_00673_));
 sky130_fd_sc_hd__a41o_2 _20313_ (.A1(_05340_),
    .A2(_10867_),
    .A3(_10798_),
    .A4(_05473_),
    .B1(_10864_),
    .X(_05486_));
 sky130_fd_sc_hd__a21oi_2 _20314_ (.A1(_10864_),
    .A2(_05482_),
    .B1(\decode.id_ex_rdsel_reg ),
    .Y(_05487_));
 sky130_fd_sc_hd__a32o_2 _20315_ (.A1(_05358_),
    .A2(_05362_),
    .A3(\decode.id_ex_rdsel_reg ),
    .B1(_05486_),
    .B2(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__and3b_2 _20316_ (.A_N(_05439_),
    .B(_05488_),
    .C(_05425_),
    .X(_05489_));
 sky130_fd_sc_hd__buf_1 _20317_ (.A(_05489_),
    .X(_00674_));
 sky130_fd_sc_hd__and3_2 _20318_ (.A(_10864_),
    .B(_10786_),
    .C(_05482_),
    .X(_05490_));
 sky130_fd_sc_hd__a21oi_2 _20319_ (.A1(_10864_),
    .A2(_05482_),
    .B1(_10786_),
    .Y(_05491_));
 sky130_fd_sc_hd__o21ai_2 _20320_ (.A1(_05490_),
    .A2(_05491_),
    .B1(_05420_),
    .Y(_05492_));
 sky130_fd_sc_hd__o211a_2 _20321_ (.A1(_05417_),
    .A2(_05367_),
    .B1(_05492_),
    .C1(_05454_),
    .X(_00675_));
 sky130_fd_sc_hd__nor2_2 _20322_ (.A(\decode.id_ex_pc_reg[24] ),
    .B(_05490_),
    .Y(_05493_));
 sky130_fd_sc_hd__and4_2 _20323_ (.A(_10864_),
    .B(_10786_),
    .C(\decode.id_ex_pc_reg[24] ),
    .D(_05482_),
    .X(_05494_));
 sky130_fd_sc_hd__o21ai_2 _20324_ (.A1(_05493_),
    .A2(_05494_),
    .B1(_05416_),
    .Y(_05495_));
 sky130_fd_sc_hd__o211a_2 _20325_ (.A1(_05420_),
    .A2(_05373_),
    .B1(_05495_),
    .C1(_05454_),
    .X(_00676_));
 sky130_fd_sc_hd__or3b_2 _20326_ (.A(_10693_),
    .B(_10725_),
    .C_N(_05490_),
    .X(_05496_));
 sky130_fd_sc_hd__a41o_2 _20327_ (.A1(_10864_),
    .A2(_10786_),
    .A3(\decode.id_ex_pc_reg[24] ),
    .A4(_05482_),
    .B1(_10790_),
    .X(_05497_));
 sky130_fd_sc_hd__a21oi_2 _20328_ (.A1(_05496_),
    .A2(_05497_),
    .B1(_05411_),
    .Y(_05498_));
 sky130_fd_sc_hd__a2111oi_2 _20329_ (.A1(_05378_),
    .A2(_05412_),
    .B1(_03517_),
    .C1(_05498_),
    .D1(_03551_),
    .Y(_00677_));
 sky130_fd_sc_hd__a21oi_2 _20330_ (.A1(_10790_),
    .A2(_05494_),
    .B1(\decode.id_ex_pc_reg[26] ),
    .Y(_05499_));
 sky130_fd_sc_hd__and3_2 _20331_ (.A(_10790_),
    .B(\decode.id_ex_pc_reg[26] ),
    .C(_05494_),
    .X(_05500_));
 sky130_fd_sc_hd__o21ai_2 _20332_ (.A1(_05499_),
    .A2(_05500_),
    .B1(_05416_),
    .Y(_05501_));
 sky130_fd_sc_hd__o211a_2 _20333_ (.A1(_05420_),
    .A2(_05384_),
    .B1(_05501_),
    .C1(_05454_),
    .X(_00678_));
 sky130_fd_sc_hd__and4_2 _20334_ (.A(_10790_),
    .B(\decode.id_ex_pc_reg[26] ),
    .C(_10854_),
    .D(_05494_),
    .X(_05502_));
 sky130_fd_sc_hd__nor2_2 _20335_ (.A(_10854_),
    .B(_05500_),
    .Y(_05503_));
 sky130_fd_sc_hd__o21ai_2 _20336_ (.A1(_05502_),
    .A2(_05503_),
    .B1(_05416_),
    .Y(_05504_));
 sky130_fd_sc_hd__o211a_2 _20337_ (.A1(_05420_),
    .A2(_05390_),
    .B1(_05504_),
    .C1(_05454_),
    .X(_00679_));
 sky130_fd_sc_hd__a41o_2 _20338_ (.A1(_10790_),
    .A2(\decode.id_ex_pc_reg[26] ),
    .A3(_10854_),
    .A4(_05494_),
    .B1(\decode.id_ex_pc_reg[28] ),
    .X(_05505_));
 sky130_fd_sc_hd__nand2_2 _20339_ (.A(\decode.id_ex_pc_reg[28] ),
    .B(_05502_),
    .Y(_05506_));
 sky130_fd_sc_hd__a21oi_2 _20340_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_05418_),
    .Y(_05507_));
 sky130_fd_sc_hd__a2111oi_2 _20341_ (.A1(_05398_),
    .A2(_05412_),
    .B1(_03517_),
    .C1(_03551_),
    .D1(_05507_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand4_2 _20342_ (.A(_10854_),
    .B(\decode.id_ex_pc_reg[28] ),
    .C(_10697_),
    .D(_05500_),
    .Y(_05508_));
 sky130_fd_sc_hd__a31o_2 _20343_ (.A1(_10854_),
    .A2(\decode.id_ex_pc_reg[28] ),
    .A3(_05500_),
    .B1(_10697_),
    .X(_05509_));
 sky130_fd_sc_hd__a21oi_2 _20344_ (.A1(_05508_),
    .A2(_05509_),
    .B1(_05418_),
    .Y(_05510_));
 sky130_fd_sc_hd__a2111oi_2 _20345_ (.A1(_05403_),
    .A2(_05418_),
    .B1(_03517_),
    .C1(_03551_),
    .D1(_05510_),
    .Y(_00681_));
 sky130_fd_sc_hd__a21oi_2 _20346_ (.A1(_05508_),
    .A2(\decode.id_ex_pc_reg[30] ),
    .B1(_05411_),
    .Y(_05511_));
 sky130_fd_sc_hd__o21a_2 _20347_ (.A1(\decode.id_ex_pc_reg[30] ),
    .A2(_05508_),
    .B1(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__a2111oi_2 _20348_ (.A1(_05406_),
    .A2(_05418_),
    .B1(_03517_),
    .C1(_03551_),
    .D1(_05512_),
    .Y(_00682_));
 sky130_fd_sc_hd__or3_2 _20349_ (.A(_10684_),
    .B(\decode.id_ex_pc_reg[31] ),
    .C(_05508_),
    .X(_05513_));
 sky130_fd_sc_hd__and4_2 _20350_ (.A(\decode.id_ex_pc_reg[28] ),
    .B(_10697_),
    .C(\decode.id_ex_pc_reg[30] ),
    .D(_05502_),
    .X(_05514_));
 sky130_fd_sc_hd__o21a_2 _20351_ (.A1(_10733_),
    .A2(_05514_),
    .B1(_05416_),
    .X(_05515_));
 sky130_fd_sc_hd__a221oi_2 _20352_ (.A1(_05513_),
    .A2(_05515_),
    .B1(_05410_),
    .B2(_05412_),
    .C1(_03588_),
    .Y(_00683_));
 sky130_fd_sc_hd__buf_1 _20353_ (.A(\csr.io_csr_address[2] ),
    .X(_05516_));
 sky130_fd_sc_hd__and4_2 _20354_ (.A(_03721_),
    .B(_03737_),
    .C(_03755_),
    .D(_05516_),
    .X(_05517_));
 sky130_fd_sc_hd__a21oi_2 _20355_ (.A1(_03741_),
    .A2(_03755_),
    .B1(_05517_),
    .Y(_05518_));
 sky130_fd_sc_hd__or4b_2 _20356_ (.A(\csr.io_csr_address[4] ),
    .B(\csr.io_csr_address[5] ),
    .C(\csr.io_csr_address[7] ),
    .D_N(\csr.io_csr_address[6] ),
    .X(_05519_));
 sky130_fd_sc_hd__and3b_2 _20357_ (.A_N(\csr.io_csr_address[10] ),
    .B(\csr.io_csr_address[9] ),
    .C(\csr.io_csr_address[8] ),
    .X(_05520_));
 sky130_fd_sc_hd__or3b_2 _20358_ (.A(_05519_),
    .B(\csr.io_csr_address[11] ),
    .C_N(_05520_),
    .X(_05521_));
 sky130_fd_sc_hd__buf_1 _20359_ (.A(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__nor4_2 _20360_ (.A(\csr.io_csr_address[4] ),
    .B(\csr.io_csr_address[5] ),
    .C(\csr.io_csr_address[7] ),
    .D(\csr.io_csr_address[6] ),
    .Y(_05523_));
 sky130_fd_sc_hd__and3_2 _20361_ (.A(_03737_),
    .B(_03741_),
    .C(_03755_),
    .X(_05524_));
 sky130_fd_sc_hd__nor2_2 _20362_ (.A(\csr.io_csr_address[2] ),
    .B(\csr.io_csr_address[3] ),
    .Y(_05525_));
 sky130_fd_sc_hd__and3_2 _20363_ (.A(_05525_),
    .B(_03721_),
    .C(_03710_),
    .X(_05526_));
 sky130_fd_sc_hd__and3b_2 _20364_ (.A_N(\csr.io_csr_address[11] ),
    .B(_05523_),
    .C(_05520_),
    .X(_05527_));
 sky130_fd_sc_hd__and3_2 _20365_ (.A(_05527_),
    .B(_03755_),
    .C(_03737_),
    .X(_05528_));
 sky130_fd_sc_hd__a41o_2 _20366_ (.A1(\csr.io_csr_address[11] ),
    .A2(_05526_),
    .A3(_05523_),
    .A4(_05520_),
    .B1(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__a41o_2 _20367_ (.A1(\csr.io_csr_address[11] ),
    .A2(_05523_),
    .A3(_05520_),
    .A4(_05524_),
    .B1(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__o21ba_2 _20368_ (.A1(_05518_),
    .A2(_05522_),
    .B1_N(_05530_),
    .X(_05531_));
 sky130_fd_sc_hd__a21oi_2 _20369_ (.A1(\decode.csr_write_reg ),
    .A2(_05531_),
    .B1(\decode.exception_out_reg ),
    .Y(_05532_));
 sky130_fd_sc_hd__o21ai_2 _20370_ (.A1(\decode.csr_write_reg ),
    .A2(_05531_),
    .B1(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__buf_1 _20371_ (.A(\csr.io_csr_address[7] ),
    .X(_05534_));
 sky130_fd_sc_hd__or4_2 _20372_ (.A(\csr.io_csr_address[4] ),
    .B(\csr.io_csr_address[5] ),
    .C(\csr.io_csr_address[6] ),
    .D(\csr.io_csr_address[8] ),
    .X(_05535_));
 sky130_fd_sc_hd__and4bb_2 _20373_ (.A_N(\csr.io_csr_address[9] ),
    .B_N(_05535_),
    .C(\csr.io_csr_address[11] ),
    .D(\csr.io_csr_address[10] ),
    .X(_05536_));
 sky130_fd_sc_hd__or4bb_2 _20374_ (.A(_03710_),
    .B(_05534_),
    .C_N(_05525_),
    .D_N(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__nand2_2 _20375_ (.A(_05526_),
    .B(_05536_),
    .Y(_05538_));
 sky130_fd_sc_hd__or4_2 _20376_ (.A(_03718_),
    .B(_03710_),
    .C(\csr.io_csr_address[3] ),
    .D(_03741_),
    .X(_05539_));
 sky130_fd_sc_hd__buf_1 _20377_ (.A(_03721_),
    .X(_05540_));
 sky130_fd_sc_hd__buf_1 _20378_ (.A(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__a211o_2 _20379_ (.A1(_05541_),
    .A2(_03737_),
    .B1(_05516_),
    .C1(\csr.io_csr_address[3] ),
    .X(_05542_));
 sky130_fd_sc_hd__nand4_2 _20380_ (.A(\csr.io_csr_address[11] ),
    .B(\csr.io_csr_address[10] ),
    .C(\csr.io_csr_address[9] ),
    .D(\csr.io_csr_address[8] ),
    .Y(_05543_));
 sky130_fd_sc_hd__or4b_2 _20381_ (.A(\csr.io_csr_address[5] ),
    .B(_05534_),
    .C(\csr.io_csr_address[6] ),
    .D_N(\csr.io_csr_address[4] ),
    .X(_05544_));
 sky130_fd_sc_hd__a211o_2 _20382_ (.A1(_05539_),
    .A2(_05542_),
    .B1(_05543_),
    .C1(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__and3_2 _20383_ (.A(_05537_),
    .B(_05538_),
    .C(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__and3_2 _20384_ (.A(\decode.csr_read_reg ),
    .B(_05531_),
    .C(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__a21oi_2 _20385_ (.A1(_05531_),
    .A2(_05546_),
    .B1(\decode.csr_read_reg ),
    .Y(_05548_));
 sky130_fd_sc_hd__o31a_2 _20386_ (.A1(_05533_),
    .A2(_05547_),
    .A3(_05548_),
    .B1(_05414_),
    .X(_00684_));
 sky130_fd_sc_hd__and3b_2 _20387_ (.A_N(_05439_),
    .B(_05201_),
    .C(\decode.io_wfi_out ),
    .X(_05549_));
 sky130_fd_sc_hd__buf_1 _20388_ (.A(_05549_),
    .X(_00685_));
 sky130_fd_sc_hd__and3b_2 _20389_ (.A_N(_05439_),
    .B(_05201_),
    .C(\decode.io_mret_out ),
    .X(_05550_));
 sky130_fd_sc_hd__buf_1 _20390_ (.A(_05550_),
    .X(_00686_));
 sky130_fd_sc_hd__and4bb_2 _20391_ (.A_N(_03710_),
    .B_N(_05534_),
    .C(_05525_),
    .D(_05536_),
    .X(_05551_));
 sky130_fd_sc_hd__buf_1 _20392_ (.A(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__or3_2 _20393_ (.A(_05534_),
    .B(\csr.minstret[0] ),
    .C(_05538_),
    .X(_05553_));
 sky130_fd_sc_hd__or4_2 _20394_ (.A(_03710_),
    .B(_05516_),
    .C(\csr.io_csr_address[3] ),
    .D(_05522_),
    .X(_05554_));
 sky130_fd_sc_hd__and4_2 _20395_ (.A(_03710_),
    .B(_05525_),
    .C(_05536_),
    .D(_05540_),
    .X(_05555_));
 sky130_fd_sc_hd__nand2_2 _20396_ (.A(_05534_),
    .B(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__or3_2 _20397_ (.A(\csr.mscratch[0] ),
    .B(_03718_),
    .C(_05554_),
    .X(_05557_));
 sky130_fd_sc_hd__o311a_2 _20398_ (.A1(_05540_),
    .A2(_05554_),
    .A3(\csr.io_mret_vector[0] ),
    .B1(_05556_),
    .C1(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__nor2_2 _20399_ (.A(_05534_),
    .B(_05538_),
    .Y(_05559_));
 sky130_fd_sc_hd__a41o_2 _20400_ (.A1(\csr.io_csr_address[11] ),
    .A2(_05526_),
    .A3(_05523_),
    .A4(_05520_),
    .B1(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__and4_2 _20401_ (.A(\csr.io_csr_address[11] ),
    .B(_05523_),
    .C(_05520_),
    .D(_05524_),
    .X(_05561_));
 sky130_fd_sc_hd__or4_2 _20402_ (.A(_03718_),
    .B(_05516_),
    .C(\csr.io_csr_address[3] ),
    .D(_03737_),
    .X(_05562_));
 sky130_fd_sc_hd__nor2_2 _20403_ (.A(_05562_),
    .B(_05522_),
    .Y(_05563_));
 sky130_fd_sc_hd__and4b_2 _20404_ (.A_N(_05522_),
    .B(_03755_),
    .C(_03741_),
    .D(_03737_),
    .X(_05564_));
 sky130_fd_sc_hd__buf_1 _20405_ (.A(_05564_),
    .X(_05565_));
 sky130_fd_sc_hd__a221o_2 _20406_ (.A1(\csr.mcycle[0] ),
    .A2(_05561_),
    .B1(_05563_),
    .B2(\csr._csr_read_data_T_9[0] ),
    .C1(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__a21o_2 _20407_ (.A1(\csr.minstret[0] ),
    .A2(_05560_),
    .B1(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__a32o_2 _20408_ (.A1(\csr._minstret_T_3[32] ),
    .A2(_05526_),
    .A3(_05536_),
    .B1(_05558_),
    .B2(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__a22o_2 _20409_ (.A1(\csr.mcycle[0] ),
    .A2(_05552_),
    .B1(_05553_),
    .B2(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__and3b_2 _20410_ (.A_N(_05439_),
    .B(_05569_),
    .C(_05425_),
    .X(_05570_));
 sky130_fd_sc_hd__buf_1 _20411_ (.A(_05570_),
    .X(_00687_));
 sky130_fd_sc_hd__and4_2 _20412_ (.A(\csr.io_csr_address[11] ),
    .B(_05526_),
    .C(_05523_),
    .D(_05520_),
    .X(_05571_));
 sky130_fd_sc_hd__buf_1 _20413_ (.A(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__buf_1 _20414_ (.A(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__buf_1 _20415_ (.A(_05573_),
    .X(_05574_));
 sky130_fd_sc_hd__buf_1 _20416_ (.A(_05559_),
    .X(_05575_));
 sky130_fd_sc_hd__o21a_2 _20417_ (.A1(_05574_),
    .A2(_05575_),
    .B1(\csr.minstret[1] ),
    .X(_05576_));
 sky130_fd_sc_hd__buf_1 _20418_ (.A(_05534_),
    .X(_05577_));
 sky130_fd_sc_hd__buf_1 _20419_ (.A(_05555_),
    .X(_05578_));
 sky130_fd_sc_hd__a32o_2 _20420_ (.A1(\csr._minstret_T_3[33] ),
    .A2(_05577_),
    .A3(_05578_),
    .B1(_05563_),
    .B2(\csr._csr_read_data_T_9[1] ),
    .X(_05579_));
 sky130_fd_sc_hd__nor2_2 _20421_ (.A(_03721_),
    .B(_05554_),
    .Y(_05580_));
 sky130_fd_sc_hd__and4b_2 _20422_ (.A_N(_05522_),
    .B(_03737_),
    .C(_03721_),
    .D(_05525_),
    .X(_05581_));
 sky130_fd_sc_hd__buf_1 _20423_ (.A(_05561_),
    .X(_05582_));
 sky130_fd_sc_hd__o21a_2 _20424_ (.A1(_05582_),
    .A2(_05551_),
    .B1(\csr.mcycle[1] ),
    .X(_05583_));
 sky130_fd_sc_hd__a221o_2 _20425_ (.A1(\csr.io_mret_vector[1] ),
    .A2(_05580_),
    .B1(_05581_),
    .B2(\csr.mscratch[1] ),
    .C1(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__o31a_2 _20426_ (.A1(_05576_),
    .A2(_05579_),
    .A3(_05584_),
    .B1(_05414_),
    .X(_00688_));
 sky130_fd_sc_hd__buf_1 _20427_ (.A(_05582_),
    .X(_05585_));
 sky130_fd_sc_hd__buf_1 _20428_ (.A(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__buf_1 _20429_ (.A(_05551_),
    .X(_05587_));
 sky130_fd_sc_hd__buf_1 _20430_ (.A(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__o21a_2 _20431_ (.A1(_05586_),
    .A2(_05588_),
    .B1(\csr.mcycle[2] ),
    .X(_05589_));
 sky130_fd_sc_hd__a22o_2 _20432_ (.A1(\csr.io_mret_vector[2] ),
    .A2(_05580_),
    .B1(_05581_),
    .B2(\csr.mscratch[2] ),
    .X(_05590_));
 sky130_fd_sc_hd__buf_1 _20433_ (.A(_03718_),
    .X(_05591_));
 sky130_fd_sc_hd__buf_1 _20434_ (.A(_05591_),
    .X(_05592_));
 sky130_fd_sc_hd__buf_1 _20435_ (.A(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__buf_1 _20436_ (.A(_05559_),
    .X(_05594_));
 sky130_fd_sc_hd__and3_2 _20437_ (.A(_05534_),
    .B(_05526_),
    .C(_05536_),
    .X(_05595_));
 sky130_fd_sc_hd__a22o_2 _20438_ (.A1(\csr.minstret[2] ),
    .A2(_05573_),
    .B1(_05563_),
    .B2(\csr._csr_read_data_T_9[2] ),
    .X(_05596_));
 sky130_fd_sc_hd__a221o_2 _20439_ (.A1(\csr.minstret[2] ),
    .A2(_05594_),
    .B1(_05595_),
    .B2(\csr._minstret_T_3[34] ),
    .C1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__a41o_2 _20440_ (.A1(\csr._csr_read_data_T_8[2] ),
    .A2(_05593_),
    .A3(_05516_),
    .A4(_05528_),
    .B1(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__o31a_2 _20441_ (.A1(_05589_),
    .A2(_05590_),
    .A3(_05598_),
    .B1(_04459_),
    .X(_00689_));
 sky130_fd_sc_hd__and3_2 _20442_ (.A(_05527_),
    .B(_05540_),
    .C(_05524_),
    .X(_05599_));
 sky130_fd_sc_hd__a221o_2 _20443_ (.A1(\csr.minstret[3] ),
    .A2(_05594_),
    .B1(_05599_),
    .B2(\csr.ie ),
    .C1(_05552_),
    .X(_05600_));
 sky130_fd_sc_hd__a31o_2 _20444_ (.A1(\csr._minstret_T_3[35] ),
    .A2(_05577_),
    .A3(_05578_),
    .B1(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__buf_1 _20445_ (.A(_05565_),
    .X(_05602_));
 sky130_fd_sc_hd__buf_1 _20446_ (.A(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__nor2_2 _20447_ (.A(_05539_),
    .B(_05522_),
    .Y(_05604_));
 sky130_fd_sc_hd__a221o_2 _20448_ (.A1(\csr.mcycle[3] ),
    .A2(_05582_),
    .B1(_05581_),
    .B2(\csr.mscratch[3] ),
    .C1(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__a31o_2 _20449_ (.A1(_05592_),
    .A2(\csr.io_mret_vector[3] ),
    .A3(_05603_),
    .B1(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__a22o_2 _20450_ (.A1(\csr.minstret[3] ),
    .A2(_05572_),
    .B1(_05563_),
    .B2(\csr._csr_read_data_T_9[3] ),
    .X(_05607_));
 sky130_fd_sc_hd__a31o_2 _20451_ (.A1(\csr.msie ),
    .A2(_05517_),
    .A3(_05527_),
    .B1(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__a41o_2 _20452_ (.A1(\csr._csr_read_data_T_8[3] ),
    .A2(_05592_),
    .A3(_05516_),
    .A4(_05528_),
    .B1(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__o32a_2 _20453_ (.A1(\csr.msip ),
    .A2(_05539_),
    .A3(_05522_),
    .B1(_05606_),
    .B2(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__o221a_2 _20454_ (.A1(\csr.mcycle[3] ),
    .A2(_05537_),
    .B1(_05601_),
    .B2(_05610_),
    .C1(_03595_),
    .X(_00690_));
 sky130_fd_sc_hd__buf_1 _20455_ (.A(_05554_),
    .X(_05611_));
 sky130_fd_sc_hd__or3_2 _20456_ (.A(\csr.mscratch[4] ),
    .B(_05592_),
    .C(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__buf_1 _20457_ (.A(\csr.minstret[4] ),
    .X(_05613_));
 sky130_fd_sc_hd__o21a_2 _20458_ (.A1(_05541_),
    .A2(\csr.io_mret_vector[4] ),
    .B1(_05602_),
    .X(_05614_));
 sky130_fd_sc_hd__a221o_2 _20459_ (.A1(_05613_),
    .A2(_05574_),
    .B1(_05586_),
    .B2(\csr.mcycle[4] ),
    .C1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__buf_1 _20460_ (.A(_05595_),
    .X(_05616_));
 sky130_fd_sc_hd__and3_2 _20461_ (.A(_03718_),
    .B(_05516_),
    .C(_05528_),
    .X(_05617_));
 sky130_fd_sc_hd__buf_1 _20462_ (.A(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__a22o_2 _20463_ (.A1(\csr.mcycle[4] ),
    .A2(_05587_),
    .B1(_05594_),
    .B2(_05613_),
    .X(_05619_));
 sky130_fd_sc_hd__a221o_2 _20464_ (.A1(\csr._minstret_T_3[36] ),
    .A2(_05616_),
    .B1(_05618_),
    .B2(\csr._csr_read_data_T_8[4] ),
    .C1(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__a21oi_2 _20465_ (.A1(_05612_),
    .A2(_05615_),
    .B1(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__nor2_2 _20466_ (.A(_05621_),
    .B(_05219_),
    .Y(_00691_));
 sky130_fd_sc_hd__buf_1 _20467_ (.A(_05618_),
    .X(_05622_));
 sky130_fd_sc_hd__a22o_2 _20468_ (.A1(\csr.mcycle[5] ),
    .A2(_05552_),
    .B1(_05575_),
    .B2(\csr.minstret[5] ),
    .X(_05623_));
 sky130_fd_sc_hd__a221o_2 _20469_ (.A1(\csr._minstret_T_3[37] ),
    .A2(_05616_),
    .B1(_05622_),
    .B2(\csr._csr_read_data_T_8[5] ),
    .C1(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__buf_1 _20470_ (.A(_05611_),
    .X(_05625_));
 sky130_fd_sc_hd__a22o_2 _20471_ (.A1(\csr.minstret[5] ),
    .A2(_05574_),
    .B1(_05586_),
    .B2(\csr.mcycle[5] ),
    .X(_05626_));
 sky130_fd_sc_hd__buf_1 _20472_ (.A(_05541_),
    .X(_05627_));
 sky130_fd_sc_hd__o21a_2 _20473_ (.A1(_05627_),
    .A2(\csr.io_mret_vector[5] ),
    .B1(_05603_),
    .X(_05628_));
 sky130_fd_sc_hd__o32a_2 _20474_ (.A1(\csr.mscratch[5] ),
    .A2(_05593_),
    .A3(_05625_),
    .B1(_05626_),
    .B2(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__buf_1 _20475_ (.A(_03594_),
    .X(_05630_));
 sky130_fd_sc_hd__o21a_2 _20476_ (.A1(_05624_),
    .A2(_05629_),
    .B1(_05630_),
    .X(_00692_));
 sky130_fd_sc_hd__a22o_2 _20477_ (.A1(\csr.mcycle[6] ),
    .A2(_05552_),
    .B1(_05575_),
    .B2(\csr.minstret[6] ),
    .X(_05631_));
 sky130_fd_sc_hd__a221o_2 _20478_ (.A1(\csr._minstret_T_3[38] ),
    .A2(_05616_),
    .B1(_05622_),
    .B2(\csr._csr_read_data_T_8[6] ),
    .C1(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__a22o_2 _20479_ (.A1(\csr.minstret[6] ),
    .A2(_05574_),
    .B1(_05586_),
    .B2(\csr.mcycle[6] ),
    .X(_05633_));
 sky130_fd_sc_hd__o21a_2 _20480_ (.A1(_05627_),
    .A2(\csr.io_mret_vector[6] ),
    .B1(_05603_),
    .X(_05634_));
 sky130_fd_sc_hd__o32a_2 _20481_ (.A1(\csr.mscratch[6] ),
    .A2(_05593_),
    .A3(_05625_),
    .B1(_05633_),
    .B2(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__o21a_2 _20482_ (.A1(_05632_),
    .A2(_05635_),
    .B1(_05630_),
    .X(_00693_));
 sky130_fd_sc_hd__or3_2 _20483_ (.A(_05534_),
    .B(\csr.minstret[7] ),
    .C(_05538_),
    .X(_05636_));
 sky130_fd_sc_hd__and3_2 _20484_ (.A(\csr.mtie ),
    .B(_05517_),
    .C(_05527_),
    .X(_05637_));
 sky130_fd_sc_hd__a221o_2 _20485_ (.A1(\csr.minstret[7] ),
    .A2(_05571_),
    .B1(_05561_),
    .B2(\csr.mcycle[7] ),
    .C1(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__a221o_2 _20486_ (.A1(\csr.io_mret_vector[7] ),
    .A2(_05580_),
    .B1(_05581_),
    .B2(\csr.mscratch[7] ),
    .C1(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__a41o_2 _20487_ (.A1(\csr._csr_read_data_T_8[7] ),
    .A2(_05591_),
    .A3(_05516_),
    .A4(_05528_),
    .B1(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__a221o_2 _20488_ (.A1(\csr._minstret_T_3[39] ),
    .A2(_05555_),
    .B1(_05599_),
    .B2(\csr.pie ),
    .C1(_05559_),
    .X(_05641_));
 sky130_fd_sc_hd__a211o_2 _20489_ (.A1(\csr.mtip ),
    .A2(_05604_),
    .B1(_05640_),
    .C1(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__a22o_2 _20490_ (.A1(\csr.mcycle[7] ),
    .A2(_05552_),
    .B1(_05636_),
    .B2(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__and3b_2 _20491_ (.A_N(_10909_),
    .B(_05643_),
    .C(_09954_),
    .X(_05644_));
 sky130_fd_sc_hd__buf_1 _20492_ (.A(_05644_),
    .X(_00694_));
 sky130_fd_sc_hd__a22o_2 _20493_ (.A1(\csr.mcycle[8] ),
    .A2(_05588_),
    .B1(_05575_),
    .B2(\csr.minstret[8] ),
    .X(_05645_));
 sky130_fd_sc_hd__a31o_2 _20494_ (.A1(_05591_),
    .A2(_03741_),
    .A3(_05528_),
    .B1(_05595_),
    .X(_05646_));
 sky130_fd_sc_hd__a41o_2 _20495_ (.A1(\csr._csr_read_data_T_8[8] ),
    .A2(_05591_),
    .A3(_05516_),
    .A4(_05528_),
    .B1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__a22o_2 _20496_ (.A1(\csr.minstret[8] ),
    .A2(_05572_),
    .B1(_05582_),
    .B2(\csr.mcycle[8] ),
    .X(_05648_));
 sky130_fd_sc_hd__a221o_2 _20497_ (.A1(\csr.io_mret_vector[8] ),
    .A2(_05580_),
    .B1(_05581_),
    .B2(\csr.mscratch[8] ),
    .C1(_05648_),
    .X(_05649_));
 sky130_fd_sc_hd__o22a_2 _20498_ (.A1(_05556_),
    .A2(\csr._minstret_T_3[40] ),
    .B1(_05647_),
    .B2(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__o21a_2 _20499_ (.A1(_05645_),
    .A2(_05650_),
    .B1(_03595_),
    .X(_00695_));
 sky130_fd_sc_hd__or3_2 _20500_ (.A(\csr.mscratch[9] ),
    .B(_05592_),
    .C(_05611_),
    .X(_05651_));
 sky130_fd_sc_hd__o21a_2 _20501_ (.A1(_05541_),
    .A2(\csr.io_mret_vector[9] ),
    .B1(_05602_),
    .X(_05652_));
 sky130_fd_sc_hd__a221o_2 _20502_ (.A1(\csr.minstret[9] ),
    .A2(_05573_),
    .B1(_05585_),
    .B2(\csr.mcycle[9] ),
    .C1(_05652_),
    .X(_05653_));
 sky130_fd_sc_hd__a22o_2 _20503_ (.A1(\csr.mcycle[9] ),
    .A2(_05587_),
    .B1(_05594_),
    .B2(\csr.minstret[9] ),
    .X(_05654_));
 sky130_fd_sc_hd__a31o_2 _20504_ (.A1(\csr._minstret_T_3[41] ),
    .A2(_05577_),
    .A3(_05578_),
    .B1(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__a221o_2 _20505_ (.A1(\csr._csr_read_data_T_8[9] ),
    .A2(_05622_),
    .B1(_05651_),
    .B2(_05653_),
    .C1(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__and3b_2 _20506_ (.A_N(_05439_),
    .B(_05656_),
    .C(_03449_),
    .X(_05657_));
 sky130_fd_sc_hd__buf_1 _20507_ (.A(_05657_),
    .X(_00696_));
 sky130_fd_sc_hd__or3b_2 _20508_ (.A(_05534_),
    .B(_05562_),
    .C_N(_05536_),
    .X(_05658_));
 sky130_fd_sc_hd__a221o_2 _20509_ (.A1(\csr._minstret_T_3[42] ),
    .A2(_05578_),
    .B1(_05617_),
    .B2(\csr._csr_read_data_T_8[10] ),
    .C1(_05559_),
    .X(_05659_));
 sky130_fd_sc_hd__a22o_2 _20510_ (.A1(\csr.minstret[10] ),
    .A2(_05572_),
    .B1(_05582_),
    .B2(\csr.mcycle[10] ),
    .X(_05660_));
 sky130_fd_sc_hd__o21a_2 _20511_ (.A1(_05540_),
    .A2(\csr.io_mret_vector[10] ),
    .B1(_05602_),
    .X(_05661_));
 sky130_fd_sc_hd__o32a_2 _20512_ (.A1(\csr.mscratch[10] ),
    .A2(_05591_),
    .A3(_05611_),
    .B1(_05660_),
    .B2(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__o221a_2 _20513_ (.A1(\csr.minstret[10] ),
    .A2(_05658_),
    .B1(_05659_),
    .B2(_05662_),
    .C1(_05537_),
    .X(_05663_));
 sky130_fd_sc_hd__a21oi_2 _20514_ (.A1(\csr.mcycle[10] ),
    .A2(_05588_),
    .B1(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__nor2_2 _20515_ (.A(_05664_),
    .B(_03587_),
    .Y(_00697_));
 sky130_fd_sc_hd__and3_2 _20516_ (.A(\csr.meie ),
    .B(_05517_),
    .C(_05527_),
    .X(_05665_));
 sky130_fd_sc_hd__a221o_2 _20517_ (.A1(\csr.minstret[11] ),
    .A2(_05573_),
    .B1(_05585_),
    .B2(\csr.mcycle[11] ),
    .C1(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__a221o_2 _20518_ (.A1(\csr.io_mret_vector[11] ),
    .A2(_05580_),
    .B1(_05581_),
    .B2(\csr.mscratch[11] ),
    .C1(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__a22o_2 _20519_ (.A1(\csr.minstret[11] ),
    .A2(_05594_),
    .B1(_05595_),
    .B2(\csr._minstret_T_3[43] ),
    .X(_05668_));
 sky130_fd_sc_hd__a221o_2 _20520_ (.A1(\csr.mcycle[11] ),
    .A2(_05552_),
    .B1(_05604_),
    .B2(io_meip),
    .C1(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__a211oi_2 _20521_ (.A1(\csr._csr_read_data_T_8[11] ),
    .A2(_05622_),
    .B1(_05667_),
    .C1(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__buf_1 _20522_ (.A(_03588_),
    .X(_05671_));
 sky130_fd_sc_hd__nor2_2 _20523_ (.A(_05670_),
    .B(_05671_),
    .Y(_00698_));
 sky130_fd_sc_hd__or3b_2 _20524_ (.A(_05540_),
    .B(_03741_),
    .C_N(_05528_),
    .X(_05672_));
 sky130_fd_sc_hd__o21a_2 _20525_ (.A1(_03721_),
    .A2(\csr.io_mret_vector[12] ),
    .B1(_05565_),
    .X(_05673_));
 sky130_fd_sc_hd__a221o_2 _20526_ (.A1(\csr.minstret[12] ),
    .A2(_05571_),
    .B1(_05561_),
    .B2(\csr.mcycle[12] ),
    .C1(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__o311a_2 _20527_ (.A1(\csr.mscratch[12] ),
    .A2(_03718_),
    .A3(_05554_),
    .B1(_05672_),
    .C1(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__a221o_2 _20528_ (.A1(_05526_),
    .A2(_05536_),
    .B1(_05617_),
    .B2(\csr._csr_read_data_T_8[12] ),
    .C1(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__o221a_2 _20529_ (.A1(\csr._minstret_T_3[44] ),
    .A2(_05556_),
    .B1(\csr.minstret[12] ),
    .B2(_05658_),
    .C1(_05537_),
    .X(_05677_));
 sky130_fd_sc_hd__a22o_2 _20530_ (.A1(\csr.mcycle[12] ),
    .A2(_05552_),
    .B1(_05676_),
    .B2(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__and3b_2 _20531_ (.A_N(_10909_),
    .B(_05678_),
    .C(_09954_),
    .X(_05679_));
 sky130_fd_sc_hd__buf_1 _20532_ (.A(_05679_),
    .X(_00699_));
 sky130_fd_sc_hd__a32o_2 _20533_ (.A1(\csr._minstret_T_3[45] ),
    .A2(_05577_),
    .A3(_05578_),
    .B1(_05552_),
    .B2(\csr.mcycle[13] ),
    .X(_05680_));
 sky130_fd_sc_hd__a221o_2 _20534_ (.A1(\csr.minstret[13] ),
    .A2(_05575_),
    .B1(_05622_),
    .B2(\csr._csr_read_data_T_8[13] ),
    .C1(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__o21a_2 _20535_ (.A1(_05541_),
    .A2(\csr.io_mret_vector[13] ),
    .B1(_05602_),
    .X(_05682_));
 sky130_fd_sc_hd__a221o_2 _20536_ (.A1(\csr.minstret[13] ),
    .A2(_05574_),
    .B1(_05586_),
    .B2(\csr.mcycle[13] ),
    .C1(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__o311a_2 _20537_ (.A1(\csr.mscratch[13] ),
    .A2(_05593_),
    .A3(_05625_),
    .B1(_05672_),
    .C1(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__o21a_2 _20538_ (.A1(_05681_),
    .A2(_05684_),
    .B1(_05414_),
    .X(_00700_));
 sky130_fd_sc_hd__a22o_2 _20539_ (.A1(\csr.mcycle[14] ),
    .A2(_05588_),
    .B1(_05575_),
    .B2(\csr.minstret[14] ),
    .X(_05685_));
 sky130_fd_sc_hd__or3_2 _20540_ (.A(\csr.mscratch[14] ),
    .B(_05591_),
    .C(_05554_),
    .X(_05686_));
 sky130_fd_sc_hd__o21a_2 _20541_ (.A1(_05540_),
    .A2(\csr.io_mret_vector[14] ),
    .B1(_05565_),
    .X(_05687_));
 sky130_fd_sc_hd__a221o_2 _20542_ (.A1(\csr.minstret[14] ),
    .A2(_05572_),
    .B1(_05582_),
    .B2(\csr.mcycle[14] ),
    .C1(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__a221o_2 _20543_ (.A1(\csr._csr_read_data_T_8[14] ),
    .A2(_05617_),
    .B1(_05686_),
    .B2(_05688_),
    .C1(_05616_),
    .X(_05689_));
 sky130_fd_sc_hd__o211a_2 _20544_ (.A1(\csr._minstret_T_3[46] ),
    .A2(_05538_),
    .B1(_05658_),
    .C1(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__o21a_2 _20545_ (.A1(_05685_),
    .A2(_05690_),
    .B1(_05630_),
    .X(_00701_));
 sky130_fd_sc_hd__buf_1 _20546_ (.A(\csr.minstret[15] ),
    .X(_05691_));
 sky130_fd_sc_hd__a22o_2 _20547_ (.A1(_05691_),
    .A2(_05572_),
    .B1(_05561_),
    .B2(\csr.mcycle[15] ),
    .X(_05692_));
 sky130_fd_sc_hd__a31o_2 _20548_ (.A1(_05591_),
    .A2(\csr.io_mret_vector[15] ),
    .A3(_05565_),
    .B1(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__a221o_2 _20549_ (.A1(\csr._minstret_T_3[47] ),
    .A2(_05555_),
    .B1(_05581_),
    .B2(\csr.mscratch[15] ),
    .C1(_05559_),
    .X(_05694_));
 sky130_fd_sc_hd__a211o_2 _20550_ (.A1(\csr._csr_read_data_T_8[15] ),
    .A2(_05617_),
    .B1(_05693_),
    .C1(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__o311a_2 _20551_ (.A1(_05577_),
    .A2(_05538_),
    .A3(_05691_),
    .B1(_05537_),
    .C1(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__a21oi_2 _20552_ (.A1(\csr.mcycle[15] ),
    .A2(_05588_),
    .B1(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__nor2_2 _20553_ (.A(_05697_),
    .B(_03587_),
    .Y(_00702_));
 sky130_fd_sc_hd__or3_2 _20554_ (.A(\csr.mscratch[16] ),
    .B(_05592_),
    .C(_05611_),
    .X(_05698_));
 sky130_fd_sc_hd__o21a_2 _20555_ (.A1(_05541_),
    .A2(\csr.io_mret_vector[16] ),
    .B1(_05602_),
    .X(_05699_));
 sky130_fd_sc_hd__a221o_2 _20556_ (.A1(\csr.minstret[16] ),
    .A2(_05573_),
    .B1(_05585_),
    .B2(\csr.mcycle[16] ),
    .C1(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__a22o_2 _20557_ (.A1(\csr.mcycle[16] ),
    .A2(_05587_),
    .B1(_05559_),
    .B2(\csr.minstret[16] ),
    .X(_05701_));
 sky130_fd_sc_hd__a31o_2 _20558_ (.A1(\csr._minstret_T_3[48] ),
    .A2(_05577_),
    .A3(_05578_),
    .B1(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__a221o_2 _20559_ (.A1(\csr._csr_read_data_T_8[16] ),
    .A2(_05622_),
    .B1(_05698_),
    .B2(_05700_),
    .C1(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__and3b_2 _20560_ (.A_N(_05439_),
    .B(_05703_),
    .C(_03449_),
    .X(_05704_));
 sky130_fd_sc_hd__buf_1 _20561_ (.A(_05704_),
    .X(_00703_));
 sky130_fd_sc_hd__or3_2 _20562_ (.A(\csr.mscratch[17] ),
    .B(_05592_),
    .C(_05625_),
    .X(_05705_));
 sky130_fd_sc_hd__o21a_2 _20563_ (.A1(_05627_),
    .A2(\csr.io_mret_vector[17] ),
    .B1(_05603_),
    .X(_05706_));
 sky130_fd_sc_hd__a221o_2 _20564_ (.A1(\csr.minstret[17] ),
    .A2(_05574_),
    .B1(_05586_),
    .B2(\csr.mcycle[17] ),
    .C1(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__a22o_2 _20565_ (.A1(\csr.minstret[17] ),
    .A2(_05594_),
    .B1(_05595_),
    .B2(\csr._minstret_T_3[49] ),
    .X(_05708_));
 sky130_fd_sc_hd__a221o_2 _20566_ (.A1(\csr.mcycle[17] ),
    .A2(_05588_),
    .B1(_05618_),
    .B2(\csr._csr_read_data_T_8[17] ),
    .C1(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__a21oi_2 _20567_ (.A1(_05705_),
    .A2(_05707_),
    .B1(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__nor2_2 _20568_ (.A(_05710_),
    .B(_05671_),
    .Y(_00704_));
 sky130_fd_sc_hd__a22o_2 _20569_ (.A1(\csr.mcycle[18] ),
    .A2(_05551_),
    .B1(_05559_),
    .B2(\csr.minstret[18] ),
    .X(_05711_));
 sky130_fd_sc_hd__a31o_2 _20570_ (.A1(\csr._minstret_T_3[50] ),
    .A2(_05577_),
    .A3(_05578_),
    .B1(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__a22o_2 _20571_ (.A1(\csr.minstret[18] ),
    .A2(_05573_),
    .B1(_05585_),
    .B2(\csr.mcycle[18] ),
    .X(_05713_));
 sky130_fd_sc_hd__o21a_2 _20572_ (.A1(_05541_),
    .A2(\csr.io_mret_vector[18] ),
    .B1(_05602_),
    .X(_05714_));
 sky130_fd_sc_hd__o32a_2 _20573_ (.A1(\csr.mscratch[18] ),
    .A2(_05592_),
    .A3(_05611_),
    .B1(_05713_),
    .B2(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__a211o_2 _20574_ (.A1(\csr._csr_read_data_T_8[18] ),
    .A2(_05622_),
    .B1(_05712_),
    .C1(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__and3b_2 _20575_ (.A_N(_05439_),
    .B(_05716_),
    .C(_03449_),
    .X(_05717_));
 sky130_fd_sc_hd__buf_1 _20576_ (.A(_05717_),
    .X(_00705_));
 sky130_fd_sc_hd__or3_2 _20577_ (.A(\csr.mscratch[19] ),
    .B(_05592_),
    .C(_05611_),
    .X(_05718_));
 sky130_fd_sc_hd__o21a_2 _20578_ (.A1(_05541_),
    .A2(\csr.io_mret_vector[19] ),
    .B1(_05602_),
    .X(_05719_));
 sky130_fd_sc_hd__a221o_2 _20579_ (.A1(\csr.minstret[19] ),
    .A2(_05573_),
    .B1(_05585_),
    .B2(_03554_),
    .C1(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__a22o_2 _20580_ (.A1(_03554_),
    .A2(_05551_),
    .B1(_05559_),
    .B2(\csr.minstret[19] ),
    .X(_05721_));
 sky130_fd_sc_hd__a31o_2 _20581_ (.A1(\csr._minstret_T_3[51] ),
    .A2(_05577_),
    .A3(_05578_),
    .B1(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__a221o_2 _20582_ (.A1(\csr._csr_read_data_T_8[19] ),
    .A2(_05622_),
    .B1(_05718_),
    .B2(_05720_),
    .C1(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__and3b_2 _20583_ (.A_N(_05439_),
    .B(_05723_),
    .C(_03449_),
    .X(_05724_));
 sky130_fd_sc_hd__buf_1 _20584_ (.A(_05724_),
    .X(_00706_));
 sky130_fd_sc_hd__a22o_2 _20585_ (.A1(\csr.mcycle[20] ),
    .A2(_05587_),
    .B1(_05575_),
    .B2(\csr.minstret[20] ),
    .X(_05725_));
 sky130_fd_sc_hd__a221o_2 _20586_ (.A1(\csr._minstret_T_3[52] ),
    .A2(_05616_),
    .B1(_05622_),
    .B2(\csr._csr_read_data_T_8[20] ),
    .C1(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__a22o_2 _20587_ (.A1(\csr.minstret[20] ),
    .A2(_05574_),
    .B1(_05586_),
    .B2(\csr.mcycle[20] ),
    .X(_05727_));
 sky130_fd_sc_hd__o21a_2 _20588_ (.A1(_05627_),
    .A2(\csr.io_mret_vector[20] ),
    .B1(_05603_),
    .X(_05728_));
 sky130_fd_sc_hd__o32a_2 _20589_ (.A1(\csr.mscratch[20] ),
    .A2(_05593_),
    .A3(_05625_),
    .B1(_05727_),
    .B2(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__o21a_2 _20590_ (.A1(_05726_),
    .A2(_05729_),
    .B1(_05630_),
    .X(_00707_));
 sky130_fd_sc_hd__a22o_2 _20591_ (.A1(\csr.mcycle[21] ),
    .A2(_05587_),
    .B1(_05575_),
    .B2(\csr.minstret[21] ),
    .X(_05730_));
 sky130_fd_sc_hd__a221o_2 _20592_ (.A1(\csr._minstret_T_3[53] ),
    .A2(_05616_),
    .B1(_05618_),
    .B2(\csr._csr_read_data_T_8[21] ),
    .C1(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__a22o_2 _20593_ (.A1(\csr.minstret[21] ),
    .A2(_05574_),
    .B1(_05586_),
    .B2(\csr.mcycle[21] ),
    .X(_05732_));
 sky130_fd_sc_hd__o21a_2 _20594_ (.A1(_05627_),
    .A2(\csr.io_mret_vector[21] ),
    .B1(_05603_),
    .X(_05733_));
 sky130_fd_sc_hd__o32a_2 _20595_ (.A1(\csr.mscratch[21] ),
    .A2(_05593_),
    .A3(_05625_),
    .B1(_05732_),
    .B2(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__o21a_2 _20596_ (.A1(_05731_),
    .A2(_05734_),
    .B1(_05630_),
    .X(_00708_));
 sky130_fd_sc_hd__a221o_2 _20597_ (.A1(\csr._minstret_T_3[54] ),
    .A2(_05578_),
    .B1(_05617_),
    .B2(\csr._csr_read_data_T_8[22] ),
    .C1(_05559_),
    .X(_05735_));
 sky130_fd_sc_hd__a22o_2 _20598_ (.A1(\csr.minstret[22] ),
    .A2(_05572_),
    .B1(_05582_),
    .B2(_03555_),
    .X(_05736_));
 sky130_fd_sc_hd__o21a_2 _20599_ (.A1(_05541_),
    .A2(\csr.io_mret_vector[22] ),
    .B1(_05602_),
    .X(_05737_));
 sky130_fd_sc_hd__o32a_2 _20600_ (.A1(\csr.mscratch[22] ),
    .A2(_05591_),
    .A3(_05611_),
    .B1(_05736_),
    .B2(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__o221a_2 _20601_ (.A1(\csr.minstret[22] ),
    .A2(_05658_),
    .B1(_05735_),
    .B2(_05738_),
    .C1(_05537_),
    .X(_05739_));
 sky130_fd_sc_hd__a21oi_2 _20602_ (.A1(_03555_),
    .A2(_05588_),
    .B1(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__nor2_2 _20603_ (.A(_05740_),
    .B(_03588_),
    .Y(_00709_));
 sky130_fd_sc_hd__or3_2 _20604_ (.A(\csr.mscratch[23] ),
    .B(_03718_),
    .C(_05554_),
    .X(_05741_));
 sky130_fd_sc_hd__o21a_2 _20605_ (.A1(_05540_),
    .A2(\csr.io_mret_vector[23] ),
    .B1(_05565_),
    .X(_05742_));
 sky130_fd_sc_hd__a221o_2 _20606_ (.A1(\csr.minstret[23] ),
    .A2(_05572_),
    .B1(_05582_),
    .B2(\csr.mcycle[23] ),
    .C1(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__and3_2 _20607_ (.A(_03737_),
    .B(_03718_),
    .C(\csr._csr_read_data_T_8[23] ),
    .X(_05744_));
 sky130_fd_sc_hd__a41o_2 _20608_ (.A1(_05516_),
    .A2(_03755_),
    .A3(_05527_),
    .A4(_05744_),
    .B1(_05555_),
    .X(_05745_));
 sky130_fd_sc_hd__a31o_2 _20609_ (.A1(_05672_),
    .A2(_05741_),
    .A3(_05743_),
    .B1(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__o221a_2 _20610_ (.A1(\csr.minstret[23] ),
    .A2(_05658_),
    .B1(_05556_),
    .B2(\csr._minstret_T_3[55] ),
    .C1(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__or2_2 _20611_ (.A(_05588_),
    .B(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__o211a_2 _20612_ (.A1(\csr.mcycle[23] ),
    .A2(_05537_),
    .B1(_05748_),
    .C1(_05454_),
    .X(_00710_));
 sky130_fd_sc_hd__a22o_2 _20613_ (.A1(\csr.mcycle[24] ),
    .A2(_05587_),
    .B1(_05575_),
    .B2(\csr.minstret[24] ),
    .X(_05749_));
 sky130_fd_sc_hd__a221o_2 _20614_ (.A1(\csr._minstret_T_3[56] ),
    .A2(_05616_),
    .B1(_05618_),
    .B2(\csr._csr_read_data_T_8[24] ),
    .C1(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__a22o_2 _20615_ (.A1(\csr.minstret[24] ),
    .A2(_05574_),
    .B1(_05586_),
    .B2(\csr.mcycle[24] ),
    .X(_05751_));
 sky130_fd_sc_hd__o21a_2 _20616_ (.A1(_05627_),
    .A2(\csr.io_mret_vector[24] ),
    .B1(_05603_),
    .X(_05752_));
 sky130_fd_sc_hd__o32a_2 _20617_ (.A1(\csr.mscratch[24] ),
    .A2(_05593_),
    .A3(_05625_),
    .B1(_05751_),
    .B2(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__o21a_2 _20618_ (.A1(_05750_),
    .A2(_05753_),
    .B1(_05630_),
    .X(_00711_));
 sky130_fd_sc_hd__or3_2 _20619_ (.A(\csr.mscratch[25] ),
    .B(_05592_),
    .C(_05611_),
    .X(_05754_));
 sky130_fd_sc_hd__o21a_2 _20620_ (.A1(_05541_),
    .A2(\csr.io_mret_vector[25] ),
    .B1(_05602_),
    .X(_05755_));
 sky130_fd_sc_hd__a221o_2 _20621_ (.A1(\csr.minstret[25] ),
    .A2(_05574_),
    .B1(_05586_),
    .B2(\csr.mcycle[25] ),
    .C1(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__a22o_2 _20622_ (.A1(\csr.minstret[25] ),
    .A2(_05594_),
    .B1(_05595_),
    .B2(\csr._minstret_T_3[57] ),
    .X(_05757_));
 sky130_fd_sc_hd__a221o_2 _20623_ (.A1(\csr.mcycle[25] ),
    .A2(_05552_),
    .B1(_05618_),
    .B2(\csr._csr_read_data_T_8[25] ),
    .C1(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__a21oi_2 _20624_ (.A1(_05754_),
    .A2(_05756_),
    .B1(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__nor2_2 _20625_ (.A(_05759_),
    .B(_05671_),
    .Y(_00712_));
 sky130_fd_sc_hd__a22o_2 _20626_ (.A1(\csr.mcycle[26] ),
    .A2(_05587_),
    .B1(_05594_),
    .B2(\csr.minstret[26] ),
    .X(_05760_));
 sky130_fd_sc_hd__a221o_2 _20627_ (.A1(\csr._minstret_T_3[58] ),
    .A2(_05616_),
    .B1(_05618_),
    .B2(\csr._csr_read_data_T_8[26] ),
    .C1(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__a22o_2 _20628_ (.A1(\csr.minstret[26] ),
    .A2(_05573_),
    .B1(_05585_),
    .B2(\csr.mcycle[26] ),
    .X(_05762_));
 sky130_fd_sc_hd__o21a_2 _20629_ (.A1(_05627_),
    .A2(\csr.io_mret_vector[26] ),
    .B1(_05603_),
    .X(_05763_));
 sky130_fd_sc_hd__o32a_2 _20630_ (.A1(\csr.mscratch[26] ),
    .A2(_05593_),
    .A3(_05625_),
    .B1(_05762_),
    .B2(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__o21a_2 _20631_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_05630_),
    .X(_00713_));
 sky130_fd_sc_hd__a22o_2 _20632_ (.A1(\csr.mcycle[27] ),
    .A2(_05587_),
    .B1(_05594_),
    .B2(\csr.minstret[27] ),
    .X(_05765_));
 sky130_fd_sc_hd__a221o_2 _20633_ (.A1(\csr._minstret_T_3[59] ),
    .A2(_05616_),
    .B1(_05618_),
    .B2(\csr._csr_read_data_T_8[27] ),
    .C1(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__a22o_2 _20634_ (.A1(\csr.minstret[27] ),
    .A2(_05573_),
    .B1(_05585_),
    .B2(\csr.mcycle[27] ),
    .X(_05767_));
 sky130_fd_sc_hd__o21a_2 _20635_ (.A1(_05627_),
    .A2(\csr.io_mret_vector[27] ),
    .B1(_05603_),
    .X(_05768_));
 sky130_fd_sc_hd__o32a_2 _20636_ (.A1(\csr.mscratch[27] ),
    .A2(_05593_),
    .A3(_05625_),
    .B1(_05767_),
    .B2(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__o21a_2 _20637_ (.A1(_05766_),
    .A2(_05769_),
    .B1(_05630_),
    .X(_00714_));
 sky130_fd_sc_hd__a22o_2 _20638_ (.A1(\csr.mcycle[28] ),
    .A2(_05587_),
    .B1(_05594_),
    .B2(\csr.minstret[28] ),
    .X(_05770_));
 sky130_fd_sc_hd__a221o_2 _20639_ (.A1(\csr._minstret_T_3[60] ),
    .A2(_05616_),
    .B1(_05618_),
    .B2(\csr._csr_read_data_T_8[28] ),
    .C1(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__a22o_2 _20640_ (.A1(\csr.minstret[28] ),
    .A2(_05573_),
    .B1(_05585_),
    .B2(\csr.mcycle[28] ),
    .X(_05772_));
 sky130_fd_sc_hd__o21a_2 _20641_ (.A1(_05627_),
    .A2(\csr.io_mret_vector[28] ),
    .B1(_05603_),
    .X(_05773_));
 sky130_fd_sc_hd__o32a_2 _20642_ (.A1(\csr.mscratch[28] ),
    .A2(_05593_),
    .A3(_05625_),
    .B1(_05772_),
    .B2(_05773_),
    .X(_05774_));
 sky130_fd_sc_hd__o21a_2 _20643_ (.A1(_05771_),
    .A2(_05774_),
    .B1(_05630_),
    .X(_00715_));
 sky130_fd_sc_hd__o21a_2 _20644_ (.A1(_05540_),
    .A2(\csr.io_mret_vector[29] ),
    .B1(_05565_),
    .X(_05775_));
 sky130_fd_sc_hd__a221o_2 _20645_ (.A1(\csr.minstret[29] ),
    .A2(_05572_),
    .B1(_05582_),
    .B2(\csr.mcycle[29] ),
    .C1(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__o311a_2 _20646_ (.A1(\csr.mscratch[29] ),
    .A2(_05591_),
    .A3(_05611_),
    .B1(_05672_),
    .C1(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__a221o_2 _20647_ (.A1(_05526_),
    .A2(_05536_),
    .B1(_05618_),
    .B2(\csr._csr_read_data_T_8[29] ),
    .C1(_05777_),
    .X(_05778_));
 sky130_fd_sc_hd__o221a_2 _20648_ (.A1(\csr._minstret_T_3[61] ),
    .A2(_05556_),
    .B1(\csr.minstret[29] ),
    .B2(_05658_),
    .C1(_05537_),
    .X(_05779_));
 sky130_fd_sc_hd__a22oi_2 _20649_ (.A1(\csr.mcycle[29] ),
    .A2(_05588_),
    .B1(_05778_),
    .B2(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__nor2_2 _20650_ (.A(_05780_),
    .B(_05671_),
    .Y(_00716_));
 sky130_fd_sc_hd__or3_2 _20651_ (.A(\csr.mscratch[30] ),
    .B(_05591_),
    .C(_05554_),
    .X(_05781_));
 sky130_fd_sc_hd__o21a_2 _20652_ (.A1(_05540_),
    .A2(\csr.io_mret_vector[30] ),
    .B1(_05565_),
    .X(_05782_));
 sky130_fd_sc_hd__a221o_2 _20653_ (.A1(\csr.minstret[30] ),
    .A2(_05572_),
    .B1(_05582_),
    .B2(\csr.mcycle[30] ),
    .C1(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__a221o_2 _20654_ (.A1(\csr._csr_read_data_T_8[30] ),
    .A2(_05617_),
    .B1(_05781_),
    .B2(_05783_),
    .C1(_05646_),
    .X(_05784_));
 sky130_fd_sc_hd__o21a_2 _20655_ (.A1(\csr._minstret_T_3[62] ),
    .A2(_05556_),
    .B1(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__a22o_2 _20656_ (.A1(\csr.mcycle[30] ),
    .A2(_05588_),
    .B1(_05575_),
    .B2(\csr.minstret[30] ),
    .X(_05786_));
 sky130_fd_sc_hd__o21a_2 _20657_ (.A1(_05785_),
    .A2(_05786_),
    .B1(_03595_),
    .X(_00717_));
 sky130_fd_sc_hd__o21a_2 _20658_ (.A1(_05585_),
    .A2(_05552_),
    .B1(\csr.mcycle[31] ),
    .X(_05787_));
 sky130_fd_sc_hd__a221o_2 _20659_ (.A1(\csr.io_mret_vector[31] ),
    .A2(_05580_),
    .B1(_05581_),
    .B2(\csr.mscratch[31] ),
    .C1(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__a32o_2 _20660_ (.A1(\csr._minstret_T_3[63] ),
    .A2(_05577_),
    .A3(_05578_),
    .B1(_05563_),
    .B2(\csr._csr_read_data_T_9[31] ),
    .X(_05789_));
 sky130_fd_sc_hd__a221o_2 _20661_ (.A1(\csr.minstret[31] ),
    .A2(_05560_),
    .B1(_05622_),
    .B2(\csr._csr_read_data_T_8[31] ),
    .C1(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__o21a_2 _20662_ (.A1(_05788_),
    .A2(_05790_),
    .B1(_03595_),
    .X(_00718_));
 sky130_fd_sc_hd__and3_2 _20663_ (.A(\decode.id_ex_funct3_reg[1] ),
    .B(_03594_),
    .C(_05569_),
    .X(_05791_));
 sky130_fd_sc_hd__a21oi_2 _20664_ (.A1(\decode.id_ex_funct3_reg[0] ),
    .A2(\decode.id_ex_funct3_reg[1] ),
    .B1(_03587_),
    .Y(_05792_));
 sky130_fd_sc_hd__mux2_2 _20665_ (.A0(\decode.id_ex_rs1_data_reg[0] ),
    .A1(\decode.id_ex_ex_rs1_reg[0] ),
    .S(_05056_),
    .X(_05793_));
 sky130_fd_sc_hd__mux2_2 _20666_ (.A0(_05791_),
    .A1(_05792_),
    .S(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__buf_1 _20667_ (.A(_05794_),
    .X(_00719_));
 sky130_fd_sc_hd__o311a_2 _20668_ (.A1(_05576_),
    .A2(_05579_),
    .A3(_05584_),
    .B1(_03594_),
    .C1(\decode.id_ex_funct3_reg[1] ),
    .X(_05795_));
 sky130_fd_sc_hd__mux2_2 _20669_ (.A0(\decode.id_ex_rs1_data_reg[1] ),
    .A1(\decode.id_ex_ex_rs1_reg[1] ),
    .S(_05056_),
    .X(_05796_));
 sky130_fd_sc_hd__mux2_2 _20670_ (.A0(_05795_),
    .A1(_05792_),
    .S(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__buf_1 _20671_ (.A(_05797_),
    .X(_00720_));
 sky130_fd_sc_hd__buf_1 _20672_ (.A(_03585_),
    .X(_05798_));
 sky130_fd_sc_hd__mux2_2 _20673_ (.A0(\decode.id_ex_rs1_data_reg[2] ),
    .A1(\decode.id_ex_ex_rs1_reg[2] ),
    .S(_05056_),
    .X(_05799_));
 sky130_fd_sc_hd__nor2_2 _20674_ (.A(_05798_),
    .B(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__buf_1 _20675_ (.A(_05792_),
    .X(_05801_));
 sky130_fd_sc_hd__a22o_2 _20676_ (.A1(_00689_),
    .A2(_05800_),
    .B1(_05801_),
    .B2(_05799_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_2 _20677_ (.A0(\decode.id_ex_rs1_data_reg[3] ),
    .A1(\decode.id_ex_ex_rs1_reg[3] ),
    .S(_05056_),
    .X(_05802_));
 sky130_fd_sc_hd__nor2_2 _20678_ (.A(_05798_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__a22o_2 _20679_ (.A1(_00690_),
    .A2(_05803_),
    .B1(_05801_),
    .B2(_05802_),
    .X(_00722_));
 sky130_fd_sc_hd__buf_1 _20680_ (.A(\decode.id_ex_funct3_reg[1] ),
    .X(_05804_));
 sky130_fd_sc_hd__buf_1 _20681_ (.A(_05630_),
    .X(_05805_));
 sky130_fd_sc_hd__mux2_2 _20682_ (.A0(\decode.id_ex_rs1_data_reg[4] ),
    .A1(\decode.id_ex_ex_rs1_reg[4] ),
    .S(_05056_),
    .X(_05806_));
 sky130_fd_sc_hd__nor2_2 _20683_ (.A(_05621_),
    .B(_05806_),
    .Y(_05807_));
 sky130_fd_sc_hd__a32o_2 _20684_ (.A1(_05804_),
    .A2(_05805_),
    .A3(_05807_),
    .B1(_05806_),
    .B2(_05801_),
    .X(_00723_));
 sky130_fd_sc_hd__buf_1 _20685_ (.A(_03728_),
    .X(_05808_));
 sky130_fd_sc_hd__buf_1 _20686_ (.A(_03728_),
    .X(_05809_));
 sky130_fd_sc_hd__a21oi_2 _20687_ (.A1(_05809_),
    .A2(\decode.id_ex_rs1_data_reg[5] ),
    .B1(_05798_),
    .Y(_05810_));
 sky130_fd_sc_hd__a32o_2 _20688_ (.A1(_05801_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[5] ),
    .B1(_05810_),
    .B2(_00692_),
    .X(_00724_));
 sky130_fd_sc_hd__a21oi_2 _20689_ (.A1(_05809_),
    .A2(\decode.id_ex_rs1_data_reg[6] ),
    .B1(_05798_),
    .Y(_05811_));
 sky130_fd_sc_hd__a32o_2 _20690_ (.A1(_05801_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[6] ),
    .B1(_05811_),
    .B2(_00693_),
    .X(_00725_));
 sky130_fd_sc_hd__a21oi_2 _20691_ (.A1(_05809_),
    .A2(\decode.id_ex_rs1_data_reg[7] ),
    .B1(_05798_),
    .Y(_05812_));
 sky130_fd_sc_hd__a32o_2 _20692_ (.A1(_05801_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[7] ),
    .B1(_05812_),
    .B2(_00694_),
    .X(_00726_));
 sky130_fd_sc_hd__buf_1 _20693_ (.A(_03728_),
    .X(_05813_));
 sky130_fd_sc_hd__nand2_2 _20694_ (.A(_05813_),
    .B(\decode.id_ex_rs1_data_reg[8] ),
    .Y(_05814_));
 sky130_fd_sc_hd__a2111oi_2 _20695_ (.A1(\decode.id_ex_funct3_reg[0] ),
    .A2(\decode.id_ex_funct3_reg[1] ),
    .B1(_05056_),
    .C1(_10575_),
    .D1(_10909_),
    .Y(_05815_));
 sky130_fd_sc_hd__a32o_2 _20696_ (.A1(_05804_),
    .A2(_00695_),
    .A3(_05814_),
    .B1(_05815_),
    .B2(\decode.id_ex_rs1_data_reg[8] ),
    .X(_00727_));
 sky130_fd_sc_hd__nand2_2 _20697_ (.A(_05813_),
    .B(\decode.id_ex_rs1_data_reg[9] ),
    .Y(_05816_));
 sky130_fd_sc_hd__a32o_2 _20698_ (.A1(_00514_),
    .A2(_05656_),
    .A3(_05816_),
    .B1(_05815_),
    .B2(\decode.id_ex_rs1_data_reg[9] ),
    .X(_00728_));
 sky130_fd_sc_hd__a21oi_2 _20699_ (.A1(_05809_),
    .A2(\decode.id_ex_rs1_data_reg[10] ),
    .B1(_05798_),
    .Y(_05817_));
 sky130_fd_sc_hd__a32o_2 _20700_ (.A1(_05801_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[10] ),
    .B1(_05817_),
    .B2(_00697_),
    .X(_00729_));
 sky130_fd_sc_hd__buf_1 _20701_ (.A(_03728_),
    .X(_05818_));
 sky130_fd_sc_hd__a21oi_2 _20702_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[11] ),
    .B1(_05670_),
    .Y(_05819_));
 sky130_fd_sc_hd__a32o_2 _20703_ (.A1(_05804_),
    .A2(_03596_),
    .A3(_05819_),
    .B1(_05815_),
    .B2(\decode.id_ex_rs1_data_reg[11] ),
    .X(_00730_));
 sky130_fd_sc_hd__a21oi_2 _20704_ (.A1(_05809_),
    .A2(\decode.id_ex_rs1_data_reg[12] ),
    .B1(_05798_),
    .Y(_05820_));
 sky130_fd_sc_hd__a32o_2 _20705_ (.A1(_05801_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[12] ),
    .B1(_05820_),
    .B2(_00699_),
    .X(_00731_));
 sky130_fd_sc_hd__nand2_2 _20706_ (.A(_03728_),
    .B(\decode.id_ex_rs1_data_reg[13] ),
    .Y(_05821_));
 sky130_fd_sc_hd__a21oi_2 _20707_ (.A1(\decode.id_ex_funct3_reg[0] ),
    .A2(_05804_),
    .B1(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__o211a_2 _20708_ (.A1(_05681_),
    .A2(_05684_),
    .B1(_05821_),
    .C1(_05804_),
    .X(_05823_));
 sky130_fd_sc_hd__o21a_2 _20709_ (.A1(_05822_),
    .A2(_05823_),
    .B1(_05414_),
    .X(_00732_));
 sky130_fd_sc_hd__a21oi_2 _20710_ (.A1(_05809_),
    .A2(\decode.id_ex_rs1_data_reg[14] ),
    .B1(_05798_),
    .Y(_05824_));
 sky130_fd_sc_hd__a32o_2 _20711_ (.A1(_05801_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[14] ),
    .B1(_05824_),
    .B2(_00701_),
    .X(_00733_));
 sky130_fd_sc_hd__a21oi_2 _20712_ (.A1(_05809_),
    .A2(\decode.id_ex_rs1_data_reg[15] ),
    .B1(_05798_),
    .Y(_05825_));
 sky130_fd_sc_hd__a32o_2 _20713_ (.A1(_05801_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[15] ),
    .B1(_05825_),
    .B2(_00702_),
    .X(_00734_));
 sky130_fd_sc_hd__nand2_2 _20714_ (.A(_05813_),
    .B(\decode.id_ex_rs1_data_reg[16] ),
    .Y(_05826_));
 sky130_fd_sc_hd__a32o_2 _20715_ (.A1(_00514_),
    .A2(_05703_),
    .A3(_05826_),
    .B1(_05815_),
    .B2(\decode.id_ex_rs1_data_reg[16] ),
    .X(_00735_));
 sky130_fd_sc_hd__a21oi_2 _20716_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[17] ),
    .B1(_05710_),
    .Y(_05827_));
 sky130_fd_sc_hd__a32o_2 _20717_ (.A1(_05804_),
    .A2(_03596_),
    .A3(_05827_),
    .B1(_05815_),
    .B2(\decode.id_ex_rs1_data_reg[17] ),
    .X(_00736_));
 sky130_fd_sc_hd__inv_2 _20718_ (.A(\decode.id_ex_rs1_data_reg[18] ),
    .Y(_05828_));
 sky130_fd_sc_hd__o221a_2 _20719_ (.A1(_05056_),
    .A2(_05828_),
    .B1(\csr.mcycle[18] ),
    .B2(_05537_),
    .C1(_05716_),
    .X(_05829_));
 sky130_fd_sc_hd__a32o_2 _20720_ (.A1(_05804_),
    .A2(_03596_),
    .A3(_05829_),
    .B1(_05815_),
    .B2(\decode.id_ex_rs1_data_reg[18] ),
    .X(_00737_));
 sky130_fd_sc_hd__nand2_2 _20721_ (.A(_05809_),
    .B(\decode.id_ex_rs1_data_reg[19] ),
    .Y(_05830_));
 sky130_fd_sc_hd__a32o_2 _20722_ (.A1(_00514_),
    .A2(_05723_),
    .A3(_05830_),
    .B1(_05815_),
    .B2(\decode.id_ex_rs1_data_reg[19] ),
    .X(_00738_));
 sky130_fd_sc_hd__buf_1 _20723_ (.A(_05792_),
    .X(_05831_));
 sky130_fd_sc_hd__a21oi_2 _20724_ (.A1(_05809_),
    .A2(\decode.id_ex_rs1_data_reg[20] ),
    .B1(_05798_),
    .Y(_05832_));
 sky130_fd_sc_hd__a32o_2 _20725_ (.A1(_05831_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[20] ),
    .B1(_05832_),
    .B2(_00707_),
    .X(_00739_));
 sky130_fd_sc_hd__a21oi_2 _20726_ (.A1(_05809_),
    .A2(\decode.id_ex_rs1_data_reg[21] ),
    .B1(_03585_),
    .Y(_05833_));
 sky130_fd_sc_hd__a32o_2 _20727_ (.A1(_05831_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[21] ),
    .B1(_05833_),
    .B2(_00708_),
    .X(_00740_));
 sky130_fd_sc_hd__nand2_2 _20728_ (.A(_03728_),
    .B(\decode.id_ex_rs1_data_reg[22] ),
    .Y(_05834_));
 sky130_fd_sc_hd__a2111oi_2 _20729_ (.A1(\decode.id_ex_funct3_reg[0] ),
    .A2(_05804_),
    .B1(_05834_),
    .C1(_03517_),
    .D1(_03581_),
    .Y(_05835_));
 sky130_fd_sc_hd__a31o_2 _20730_ (.A1(_05804_),
    .A2(_00709_),
    .A3(_05834_),
    .B1(_05835_),
    .X(_00741_));
 sky130_fd_sc_hd__inv_2 _20731_ (.A(\decode.id_ex_rs1_data_reg[23] ),
    .Y(_05836_));
 sky130_fd_sc_hd__o221a_2 _20732_ (.A1(_05056_),
    .A2(_05836_),
    .B1(\csr.mcycle[23] ),
    .B2(_05537_),
    .C1(_05748_),
    .X(_05837_));
 sky130_fd_sc_hd__a32o_2 _20733_ (.A1(_05831_),
    .A2(_05808_),
    .A3(\decode.id_ex_rs1_data_reg[23] ),
    .B1(_05837_),
    .B2(_00514_),
    .X(_00742_));
 sky130_fd_sc_hd__a21oi_2 _20734_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[24] ),
    .B1(_03585_),
    .Y(_05838_));
 sky130_fd_sc_hd__a32o_2 _20735_ (.A1(_05831_),
    .A2(_05813_),
    .A3(\decode.id_ex_rs1_data_reg[24] ),
    .B1(_05838_),
    .B2(_00711_),
    .X(_00743_));
 sky130_fd_sc_hd__a21oi_2 _20736_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[25] ),
    .B1(_05759_),
    .Y(_05839_));
 sky130_fd_sc_hd__a32o_2 _20737_ (.A1(_05804_),
    .A2(_03596_),
    .A3(_05839_),
    .B1(_05815_),
    .B2(\decode.id_ex_rs1_data_reg[25] ),
    .X(_00744_));
 sky130_fd_sc_hd__a21oi_2 _20738_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[26] ),
    .B1(_03585_),
    .Y(_05840_));
 sky130_fd_sc_hd__a32o_2 _20739_ (.A1(_05831_),
    .A2(_05813_),
    .A3(\decode.id_ex_rs1_data_reg[26] ),
    .B1(_05840_),
    .B2(_00713_),
    .X(_00745_));
 sky130_fd_sc_hd__a21oi_2 _20740_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[27] ),
    .B1(_03585_),
    .Y(_05841_));
 sky130_fd_sc_hd__a32o_2 _20741_ (.A1(_05831_),
    .A2(_05813_),
    .A3(\decode.id_ex_rs1_data_reg[27] ),
    .B1(_05841_),
    .B2(_00714_),
    .X(_00746_));
 sky130_fd_sc_hd__a21oi_2 _20742_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[28] ),
    .B1(_03585_),
    .Y(_05842_));
 sky130_fd_sc_hd__a32o_2 _20743_ (.A1(_05831_),
    .A2(_05813_),
    .A3(\decode.id_ex_rs1_data_reg[28] ),
    .B1(_05842_),
    .B2(_00715_),
    .X(_00747_));
 sky130_fd_sc_hd__a21oi_2 _20744_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[29] ),
    .B1(_05780_),
    .Y(_05843_));
 sky130_fd_sc_hd__a32o_2 _20745_ (.A1(_05831_),
    .A2(_05813_),
    .A3(\decode.id_ex_rs1_data_reg[29] ),
    .B1(_05843_),
    .B2(_00514_),
    .X(_00748_));
 sky130_fd_sc_hd__a21oi_2 _20746_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[30] ),
    .B1(_03585_),
    .Y(_05844_));
 sky130_fd_sc_hd__a32o_2 _20747_ (.A1(_05831_),
    .A2(_05813_),
    .A3(\decode.id_ex_rs1_data_reg[30] ),
    .B1(_05844_),
    .B2(_00717_),
    .X(_00749_));
 sky130_fd_sc_hd__a21oi_2 _20748_ (.A1(_05818_),
    .A2(\decode.id_ex_rs1_data_reg[31] ),
    .B1(_03585_),
    .Y(_05845_));
 sky130_fd_sc_hd__a32o_2 _20749_ (.A1(_05831_),
    .A2(_05813_),
    .A3(\decode.id_ex_rs1_data_reg[31] ),
    .B1(_05845_),
    .B2(_00718_),
    .X(_00750_));
 sky130_fd_sc_hd__nor2_2 _20750_ (.A(_05627_),
    .B(_05671_),
    .Y(_00751_));
 sky130_fd_sc_hd__nor2_2 _20751_ (.A(_03737_),
    .B(_05671_),
    .Y(_00752_));
 sky130_fd_sc_hd__nor2_2 _20752_ (.A(_03741_),
    .B(_05671_),
    .Y(_00753_));
 sky130_fd_sc_hd__nor2_2 _20753_ (.A(_03755_),
    .B(_05671_),
    .Y(_00754_));
 sky130_fd_sc_hd__and2_2 _20754_ (.A(\csr.io_csr_address[4] ),
    .B(_05214_),
    .X(_05846_));
 sky130_fd_sc_hd__buf_1 _20755_ (.A(_05846_),
    .X(_00755_));
 sky130_fd_sc_hd__and3b_2 _20756_ (.A_N(_05439_),
    .B(_05201_),
    .C(\csr.io_csr_address[5] ),
    .X(_05847_));
 sky130_fd_sc_hd__buf_1 _20757_ (.A(_05847_),
    .X(_00756_));
 sky130_fd_sc_hd__and3b_2 _20758_ (.A_N(_03452_),
    .B(_05201_),
    .C(\csr.io_csr_address[6] ),
    .X(_05848_));
 sky130_fd_sc_hd__buf_1 _20759_ (.A(_05848_),
    .X(_00757_));
 sky130_fd_sc_hd__and3b_2 _20760_ (.A_N(_03452_),
    .B(_05425_),
    .C(_05577_),
    .X(_05849_));
 sky130_fd_sc_hd__buf_1 _20761_ (.A(_05849_),
    .X(_00758_));
 sky130_fd_sc_hd__and3b_2 _20762_ (.A_N(_03452_),
    .B(_05425_),
    .C(\csr.io_csr_address[8] ),
    .X(_05850_));
 sky130_fd_sc_hd__buf_1 _20763_ (.A(_05850_),
    .X(_00759_));
 sky130_fd_sc_hd__and3b_2 _20764_ (.A_N(_03452_),
    .B(_05425_),
    .C(\csr.io_csr_address[9] ),
    .X(_05851_));
 sky130_fd_sc_hd__buf_1 _20765_ (.A(_05851_),
    .X(_00760_));
 sky130_fd_sc_hd__and3b_2 _20766_ (.A_N(_03452_),
    .B(_05425_),
    .C(\csr.io_csr_address[10] ),
    .X(_05852_));
 sky130_fd_sc_hd__buf_1 _20767_ (.A(_05852_),
    .X(_00761_));
 sky130_fd_sc_hd__and3b_2 _20768_ (.A_N(_03452_),
    .B(_05425_),
    .C(\csr.io_csr_address[11] ),
    .X(_05853_));
 sky130_fd_sc_hd__buf_1 _20769_ (.A(_05853_),
    .X(_00762_));
 sky130_fd_sc_hd__and3b_2 _20770_ (.A_N(_03452_),
    .B(_05425_),
    .C(\decode.csr_write_reg ),
    .X(_05854_));
 sky130_fd_sc_hd__buf_1 _20771_ (.A(_05854_),
    .X(_00763_));
 sky130_fd_sc_hd__and4b_2 _20772_ (.A_N(_03452_),
    .B(_10668_),
    .C(_10916_),
    .D(_10018_),
    .X(_05855_));
 sky130_fd_sc_hd__buf_1 _20773_ (.A(_05855_),
    .X(_00764_));
 sky130_fd_sc_hd__buf_1 _20774_ (.A(_10018_),
    .X(_05856_));
 sky130_fd_sc_hd__buf_1 _20775_ (.A(_03590_),
    .X(_05857_));
 sky130_fd_sc_hd__buf_1 _20776_ (.A(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__or2_2 _20777_ (.A(io_memory_address[0]),
    .B(io_memory_size[0]),
    .X(_05859_));
 sky130_fd_sc_hd__nand2_2 _20778_ (.A(io_memory_address[0]),
    .B(io_memory_size[0]),
    .Y(_05860_));
 sky130_fd_sc_hd__o21bai_2 _20779_ (.A1(io_memory_size[0]),
    .A2(\execute.io_mem_zero ),
    .B1_N(io_memory_size[1]),
    .Y(_05861_));
 sky130_fd_sc_hd__a211oi_2 _20780_ (.A1(io_memory_size[0]),
    .A2(\execute.io_mem_zero ),
    .B1(io_load_store_unsigned),
    .C1(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__a31o_2 _20781_ (.A1(io_load_store_unsigned),
    .A2(_05859_),
    .A3(_05860_),
    .B1(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__buf_1 _20782_ (.A(_03590_),
    .X(_05864_));
 sky130_fd_sc_hd__and3_2 _20783_ (.A(_05864_),
    .B(_09954_),
    .C(\execute.io_mem_isbranch ),
    .X(_05865_));
 sky130_fd_sc_hd__buf_1 _20784_ (.A(_05865_),
    .X(_01176_));
 sky130_fd_sc_hd__a32o_2 _20785_ (.A1(_05856_),
    .A2(\execute.io_mem_isjump ),
    .A3(_05858_),
    .B1(_05863_),
    .B2(_01176_),
    .X(_00765_));
 sky130_fd_sc_hd__buf_1 _20786_ (.A(_03590_),
    .X(_05866_));
 sky130_fd_sc_hd__buf_1 _20787_ (.A(_05866_),
    .X(_05867_));
 sky130_fd_sc_hd__buf_1 _20788_ (.A(_09955_),
    .X(_05868_));
 sky130_fd_sc_hd__and3_2 _20789_ (.A(\execute.io_mem_rd[0] ),
    .B(_05867_),
    .C(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__buf_1 _20790_ (.A(_05869_),
    .X(_00766_));
 sky130_fd_sc_hd__and3_2 _20791_ (.A(\execute.io_mem_rd[1] ),
    .B(_05867_),
    .C(_05868_),
    .X(_05870_));
 sky130_fd_sc_hd__buf_1 _20792_ (.A(_05870_),
    .X(_00767_));
 sky130_fd_sc_hd__and3_2 _20793_ (.A(\execute.io_mem_rd[2] ),
    .B(_05867_),
    .C(_05868_),
    .X(_05871_));
 sky130_fd_sc_hd__buf_1 _20794_ (.A(_05871_),
    .X(_00768_));
 sky130_fd_sc_hd__and3_2 _20795_ (.A(\execute.io_mem_rd[3] ),
    .B(_05867_),
    .C(_05868_),
    .X(_05872_));
 sky130_fd_sc_hd__buf_1 _20796_ (.A(_05872_),
    .X(_00769_));
 sky130_fd_sc_hd__and3_2 _20797_ (.A(\execute.io_mem_rd[4] ),
    .B(_05867_),
    .C(_05868_),
    .X(_05873_));
 sky130_fd_sc_hd__buf_1 _20798_ (.A(_05873_),
    .X(_00770_));
 sky130_fd_sc_hd__and3_2 _20799_ (.A(\execute.io_mem_regwrite ),
    .B(_05867_),
    .C(_05868_),
    .X(_05874_));
 sky130_fd_sc_hd__buf_1 _20800_ (.A(_05874_),
    .X(_00771_));
 sky130_fd_sc_hd__buf_1 _20801_ (.A(_03582_),
    .X(_05875_));
 sky130_fd_sc_hd__and3_2 _20802_ (.A(\execute.io_mem_memtoreg[0] ),
    .B(_05867_),
    .C(_05875_),
    .X(_05876_));
 sky130_fd_sc_hd__buf_1 _20803_ (.A(_05876_),
    .X(_00772_));
 sky130_fd_sc_hd__and3_2 _20804_ (.A(\execute.io_mem_memtoreg[1] ),
    .B(_05867_),
    .C(_05875_),
    .X(_05877_));
 sky130_fd_sc_hd__buf_1 _20805_ (.A(_05877_),
    .X(_00773_));
 sky130_fd_sc_hd__and3_2 _20806_ (.A(io_memory_address[0]),
    .B(_05867_),
    .C(_05875_),
    .X(_05878_));
 sky130_fd_sc_hd__buf_1 _20807_ (.A(_05878_),
    .X(_00774_));
 sky130_fd_sc_hd__buf_1 _20808_ (.A(_05866_),
    .X(_05879_));
 sky130_fd_sc_hd__and3_2 _20809_ (.A(io_memory_address[1]),
    .B(_05879_),
    .C(_05875_),
    .X(_05880_));
 sky130_fd_sc_hd__buf_1 _20810_ (.A(_05880_),
    .X(_00775_));
 sky130_fd_sc_hd__and3_2 _20811_ (.A(io_memory_address[2]),
    .B(_05879_),
    .C(_05875_),
    .X(_05881_));
 sky130_fd_sc_hd__buf_1 _20812_ (.A(_05881_),
    .X(_00776_));
 sky130_fd_sc_hd__and3_2 _20813_ (.A(io_memory_address[3]),
    .B(_05879_),
    .C(_05875_),
    .X(_05882_));
 sky130_fd_sc_hd__buf_1 _20814_ (.A(_05882_),
    .X(_00777_));
 sky130_fd_sc_hd__and3_2 _20815_ (.A(io_memory_address[4]),
    .B(_05879_),
    .C(_05875_),
    .X(_05883_));
 sky130_fd_sc_hd__buf_1 _20816_ (.A(_05883_),
    .X(_00778_));
 sky130_fd_sc_hd__and3_2 _20817_ (.A(io_memory_address[5]),
    .B(_05879_),
    .C(_05875_),
    .X(_05884_));
 sky130_fd_sc_hd__buf_1 _20818_ (.A(_05884_),
    .X(_00779_));
 sky130_fd_sc_hd__and3_2 _20819_ (.A(io_memory_address[6]),
    .B(_05879_),
    .C(_05875_),
    .X(_05885_));
 sky130_fd_sc_hd__buf_1 _20820_ (.A(_05885_),
    .X(_00780_));
 sky130_fd_sc_hd__and3_2 _20821_ (.A(io_memory_address[7]),
    .B(_05879_),
    .C(_05875_),
    .X(_05886_));
 sky130_fd_sc_hd__buf_1 _20822_ (.A(_05886_),
    .X(_00781_));
 sky130_fd_sc_hd__buf_1 _20823_ (.A(_03582_),
    .X(_05887_));
 sky130_fd_sc_hd__and3_2 _20824_ (.A(io_memory_address[8]),
    .B(_05879_),
    .C(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__buf_1 _20825_ (.A(_05888_),
    .X(_00782_));
 sky130_fd_sc_hd__and3_2 _20826_ (.A(io_memory_address[9]),
    .B(_05879_),
    .C(_05887_),
    .X(_05889_));
 sky130_fd_sc_hd__buf_1 _20827_ (.A(_05889_),
    .X(_00783_));
 sky130_fd_sc_hd__and3_2 _20828_ (.A(io_memory_address[10]),
    .B(_05879_),
    .C(_05887_),
    .X(_05890_));
 sky130_fd_sc_hd__buf_1 _20829_ (.A(_05890_),
    .X(_00784_));
 sky130_fd_sc_hd__buf_1 _20830_ (.A(_05866_),
    .X(_05891_));
 sky130_fd_sc_hd__and3_2 _20831_ (.A(io_memory_address[11]),
    .B(_05891_),
    .C(_05887_),
    .X(_05892_));
 sky130_fd_sc_hd__buf_1 _20832_ (.A(_05892_),
    .X(_00785_));
 sky130_fd_sc_hd__and3_2 _20833_ (.A(io_memory_address[12]),
    .B(_05891_),
    .C(_05887_),
    .X(_05893_));
 sky130_fd_sc_hd__buf_1 _20834_ (.A(_05893_),
    .X(_00786_));
 sky130_fd_sc_hd__and3_2 _20835_ (.A(io_memory_address[13]),
    .B(_05891_),
    .C(_05887_),
    .X(_05894_));
 sky130_fd_sc_hd__buf_1 _20836_ (.A(_05894_),
    .X(_00787_));
 sky130_fd_sc_hd__and3_2 _20837_ (.A(io_memory_address[14]),
    .B(_05891_),
    .C(_05887_),
    .X(_05895_));
 sky130_fd_sc_hd__buf_1 _20838_ (.A(_05895_),
    .X(_00788_));
 sky130_fd_sc_hd__and3_2 _20839_ (.A(io_memory_address[15]),
    .B(_05891_),
    .C(_05887_),
    .X(_05896_));
 sky130_fd_sc_hd__buf_1 _20840_ (.A(_05896_),
    .X(_00789_));
 sky130_fd_sc_hd__and3_2 _20841_ (.A(io_memory_address[16]),
    .B(_05891_),
    .C(_05887_),
    .X(_05897_));
 sky130_fd_sc_hd__buf_1 _20842_ (.A(_05897_),
    .X(_00790_));
 sky130_fd_sc_hd__and3_2 _20843_ (.A(io_memory_address[17]),
    .B(_05891_),
    .C(_05887_),
    .X(_05898_));
 sky130_fd_sc_hd__buf_1 _20844_ (.A(_05898_),
    .X(_00791_));
 sky130_fd_sc_hd__buf_1 _20845_ (.A(_03582_),
    .X(_05899_));
 sky130_fd_sc_hd__and3_2 _20846_ (.A(io_memory_address[18]),
    .B(_05891_),
    .C(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__buf_1 _20847_ (.A(_05900_),
    .X(_00792_));
 sky130_fd_sc_hd__and3_2 _20848_ (.A(io_memory_address[19]),
    .B(_05891_),
    .C(_05899_),
    .X(_05901_));
 sky130_fd_sc_hd__buf_1 _20849_ (.A(_05901_),
    .X(_00793_));
 sky130_fd_sc_hd__and3_2 _20850_ (.A(io_memory_address[20]),
    .B(_05891_),
    .C(_05899_),
    .X(_05902_));
 sky130_fd_sc_hd__buf_1 _20851_ (.A(_05902_),
    .X(_00794_));
 sky130_fd_sc_hd__buf_1 _20852_ (.A(_05866_),
    .X(_05903_));
 sky130_fd_sc_hd__and3_2 _20853_ (.A(io_memory_address[21]),
    .B(_05903_),
    .C(_05899_),
    .X(_05904_));
 sky130_fd_sc_hd__buf_1 _20854_ (.A(_05904_),
    .X(_00795_));
 sky130_fd_sc_hd__and3_2 _20855_ (.A(io_memory_address[22]),
    .B(_05903_),
    .C(_05899_),
    .X(_05905_));
 sky130_fd_sc_hd__buf_1 _20856_ (.A(_05905_),
    .X(_00796_));
 sky130_fd_sc_hd__and3_2 _20857_ (.A(io_memory_address[23]),
    .B(_05903_),
    .C(_05899_),
    .X(_05906_));
 sky130_fd_sc_hd__buf_1 _20858_ (.A(_05906_),
    .X(_00797_));
 sky130_fd_sc_hd__and3_2 _20859_ (.A(io_memory_address[24]),
    .B(_05903_),
    .C(_05899_),
    .X(_05907_));
 sky130_fd_sc_hd__buf_1 _20860_ (.A(_05907_),
    .X(_00798_));
 sky130_fd_sc_hd__and3_2 _20861_ (.A(io_memory_address[25]),
    .B(_05903_),
    .C(_05899_),
    .X(_05908_));
 sky130_fd_sc_hd__buf_1 _20862_ (.A(_05908_),
    .X(_00799_));
 sky130_fd_sc_hd__and3_2 _20863_ (.A(io_memory_address[26]),
    .B(_05903_),
    .C(_05899_),
    .X(_05909_));
 sky130_fd_sc_hd__buf_1 _20864_ (.A(_05909_),
    .X(_00800_));
 sky130_fd_sc_hd__and3_2 _20865_ (.A(io_memory_address[27]),
    .B(_05903_),
    .C(_05899_),
    .X(_05910_));
 sky130_fd_sc_hd__buf_1 _20866_ (.A(_05910_),
    .X(_00801_));
 sky130_fd_sc_hd__buf_1 _20867_ (.A(_03582_),
    .X(_05911_));
 sky130_fd_sc_hd__and3_2 _20868_ (.A(io_memory_address[28]),
    .B(_05903_),
    .C(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__buf_1 _20869_ (.A(_05912_),
    .X(_00802_));
 sky130_fd_sc_hd__and3_2 _20870_ (.A(io_memory_address[29]),
    .B(_05903_),
    .C(_05911_),
    .X(_05913_));
 sky130_fd_sc_hd__buf_1 _20871_ (.A(_05913_),
    .X(_00803_));
 sky130_fd_sc_hd__and3_2 _20872_ (.A(io_memory_address[30]),
    .B(_05903_),
    .C(_05911_),
    .X(_05914_));
 sky130_fd_sc_hd__buf_1 _20873_ (.A(_05914_),
    .X(_00804_));
 sky130_fd_sc_hd__buf_1 _20874_ (.A(_05866_),
    .X(_05915_));
 sky130_fd_sc_hd__and3_2 _20875_ (.A(io_memory_address[31]),
    .B(_05915_),
    .C(_05911_),
    .X(_05916_));
 sky130_fd_sc_hd__buf_1 _20876_ (.A(_05916_),
    .X(_00805_));
 sky130_fd_sc_hd__and3_2 _20877_ (.A(_05858_),
    .B(_09956_),
    .C(io_memory_read_data[0]),
    .X(_05917_));
 sky130_fd_sc_hd__buf_1 _20878_ (.A(_05917_),
    .X(_00806_));
 sky130_fd_sc_hd__and3_2 _20879_ (.A(_05858_),
    .B(_09956_),
    .C(io_memory_read_data[1]),
    .X(_05918_));
 sky130_fd_sc_hd__buf_1 _20880_ (.A(_05918_),
    .X(_00807_));
 sky130_fd_sc_hd__and3_2 _20881_ (.A(_05858_),
    .B(_09956_),
    .C(io_memory_read_data[2]),
    .X(_05919_));
 sky130_fd_sc_hd__buf_1 _20882_ (.A(_05919_),
    .X(_00808_));
 sky130_fd_sc_hd__and3_2 _20883_ (.A(_05858_),
    .B(_09956_),
    .C(io_memory_read_data[3]),
    .X(_05920_));
 sky130_fd_sc_hd__buf_1 _20884_ (.A(_05920_),
    .X(_00809_));
 sky130_fd_sc_hd__buf_1 _20885_ (.A(_09955_),
    .X(_05921_));
 sky130_fd_sc_hd__and3_2 _20886_ (.A(_05858_),
    .B(_05921_),
    .C(io_memory_read_data[4]),
    .X(_05922_));
 sky130_fd_sc_hd__buf_1 _20887_ (.A(_05922_),
    .X(_00810_));
 sky130_fd_sc_hd__and3_2 _20888_ (.A(_05858_),
    .B(_05921_),
    .C(io_memory_read_data[5]),
    .X(_05923_));
 sky130_fd_sc_hd__buf_1 _20889_ (.A(_05923_),
    .X(_00811_));
 sky130_fd_sc_hd__and3_2 _20890_ (.A(_05858_),
    .B(_05921_),
    .C(io_memory_read_data[6]),
    .X(_05924_));
 sky130_fd_sc_hd__buf_1 _20891_ (.A(_05924_),
    .X(_00812_));
 sky130_fd_sc_hd__buf_1 _20892_ (.A(_05857_),
    .X(_05925_));
 sky130_fd_sc_hd__and3_2 _20893_ (.A(_05925_),
    .B(_05921_),
    .C(io_memory_read_data[7]),
    .X(_05926_));
 sky130_fd_sc_hd__buf_1 _20894_ (.A(_05926_),
    .X(_00813_));
 sky130_fd_sc_hd__and3_2 _20895_ (.A(_05925_),
    .B(_05921_),
    .C(io_memory_read_data[8]),
    .X(_05927_));
 sky130_fd_sc_hd__buf_1 _20896_ (.A(_05927_),
    .X(_00814_));
 sky130_fd_sc_hd__and3_2 _20897_ (.A(_05925_),
    .B(_05921_),
    .C(io_memory_read_data[9]),
    .X(_05928_));
 sky130_fd_sc_hd__buf_1 _20898_ (.A(_05928_),
    .X(_00815_));
 sky130_fd_sc_hd__and3_2 _20899_ (.A(_05925_),
    .B(_05921_),
    .C(io_memory_read_data[10]),
    .X(_05929_));
 sky130_fd_sc_hd__buf_1 _20900_ (.A(_05929_),
    .X(_00816_));
 sky130_fd_sc_hd__and3_2 _20901_ (.A(_05925_),
    .B(_05921_),
    .C(io_memory_read_data[11]),
    .X(_05930_));
 sky130_fd_sc_hd__buf_1 _20902_ (.A(_05930_),
    .X(_00817_));
 sky130_fd_sc_hd__and3_2 _20903_ (.A(_05925_),
    .B(_05921_),
    .C(io_memory_read_data[12]),
    .X(_05931_));
 sky130_fd_sc_hd__buf_1 _20904_ (.A(_05931_),
    .X(_00818_));
 sky130_fd_sc_hd__and3_2 _20905_ (.A(_05925_),
    .B(_05921_),
    .C(io_memory_read_data[13]),
    .X(_05932_));
 sky130_fd_sc_hd__buf_1 _20906_ (.A(_05932_),
    .X(_00819_));
 sky130_fd_sc_hd__buf_1 _20907_ (.A(_09955_),
    .X(_05933_));
 sky130_fd_sc_hd__and3_2 _20908_ (.A(_05925_),
    .B(_05933_),
    .C(io_memory_read_data[14]),
    .X(_05934_));
 sky130_fd_sc_hd__buf_1 _20909_ (.A(_05934_),
    .X(_00820_));
 sky130_fd_sc_hd__and3_2 _20910_ (.A(_05925_),
    .B(_05933_),
    .C(io_memory_read_data[15]),
    .X(_05935_));
 sky130_fd_sc_hd__buf_1 _20911_ (.A(_05935_),
    .X(_00821_));
 sky130_fd_sc_hd__and3_2 _20912_ (.A(_05925_),
    .B(_05933_),
    .C(io_memory_read_data[16]),
    .X(_05936_));
 sky130_fd_sc_hd__buf_1 _20913_ (.A(_05936_),
    .X(_00822_));
 sky130_fd_sc_hd__buf_1 _20914_ (.A(_05857_),
    .X(_05937_));
 sky130_fd_sc_hd__and3_2 _20915_ (.A(_05937_),
    .B(_05933_),
    .C(io_memory_read_data[17]),
    .X(_05938_));
 sky130_fd_sc_hd__buf_1 _20916_ (.A(_05938_),
    .X(_00823_));
 sky130_fd_sc_hd__and3_2 _20917_ (.A(_05937_),
    .B(_05933_),
    .C(io_memory_read_data[18]),
    .X(_05939_));
 sky130_fd_sc_hd__buf_1 _20918_ (.A(_05939_),
    .X(_00824_));
 sky130_fd_sc_hd__and3_2 _20919_ (.A(_05937_),
    .B(_05933_),
    .C(io_memory_read_data[19]),
    .X(_05940_));
 sky130_fd_sc_hd__buf_1 _20920_ (.A(_05940_),
    .X(_00825_));
 sky130_fd_sc_hd__and3_2 _20921_ (.A(_05937_),
    .B(_05933_),
    .C(io_memory_read_data[20]),
    .X(_05941_));
 sky130_fd_sc_hd__buf_1 _20922_ (.A(_05941_),
    .X(_00826_));
 sky130_fd_sc_hd__and3_2 _20923_ (.A(_05937_),
    .B(_05933_),
    .C(io_memory_read_data[21]),
    .X(_05942_));
 sky130_fd_sc_hd__buf_1 _20924_ (.A(_05942_),
    .X(_00827_));
 sky130_fd_sc_hd__and3_2 _20925_ (.A(_05937_),
    .B(_05933_),
    .C(io_memory_read_data[22]),
    .X(_05943_));
 sky130_fd_sc_hd__buf_1 _20926_ (.A(_05943_),
    .X(_00828_));
 sky130_fd_sc_hd__and3_2 _20927_ (.A(_05937_),
    .B(_05933_),
    .C(io_memory_read_data[23]),
    .X(_05944_));
 sky130_fd_sc_hd__buf_1 _20928_ (.A(_05944_),
    .X(_00829_));
 sky130_fd_sc_hd__buf_1 _20929_ (.A(_09955_),
    .X(_05945_));
 sky130_fd_sc_hd__and3_2 _20930_ (.A(_05937_),
    .B(_05945_),
    .C(io_memory_read_data[24]),
    .X(_05946_));
 sky130_fd_sc_hd__buf_1 _20931_ (.A(_05946_),
    .X(_00830_));
 sky130_fd_sc_hd__and3_2 _20932_ (.A(_05937_),
    .B(_05945_),
    .C(io_memory_read_data[25]),
    .X(_05947_));
 sky130_fd_sc_hd__buf_1 _20933_ (.A(_05947_),
    .X(_00831_));
 sky130_fd_sc_hd__and3_2 _20934_ (.A(_05937_),
    .B(_05945_),
    .C(io_memory_read_data[26]),
    .X(_05948_));
 sky130_fd_sc_hd__buf_1 _20935_ (.A(_05948_),
    .X(_00832_));
 sky130_fd_sc_hd__buf_1 _20936_ (.A(_05857_),
    .X(_05949_));
 sky130_fd_sc_hd__and3_2 _20937_ (.A(_05949_),
    .B(_05945_),
    .C(io_memory_read_data[27]),
    .X(_05950_));
 sky130_fd_sc_hd__buf_1 _20938_ (.A(_05950_),
    .X(_00833_));
 sky130_fd_sc_hd__and3_2 _20939_ (.A(_05949_),
    .B(_05945_),
    .C(io_memory_read_data[28]),
    .X(_05951_));
 sky130_fd_sc_hd__buf_1 _20940_ (.A(_05951_),
    .X(_00834_));
 sky130_fd_sc_hd__and3_2 _20941_ (.A(_05949_),
    .B(_05945_),
    .C(io_memory_read_data[29]),
    .X(_05952_));
 sky130_fd_sc_hd__buf_1 _20942_ (.A(_05952_),
    .X(_00835_));
 sky130_fd_sc_hd__and3_2 _20943_ (.A(_05949_),
    .B(_05945_),
    .C(io_memory_read_data[30]),
    .X(_05953_));
 sky130_fd_sc_hd__buf_1 _20944_ (.A(_05953_),
    .X(_00836_));
 sky130_fd_sc_hd__and3_2 _20945_ (.A(_05949_),
    .B(_05945_),
    .C(io_memory_read_data[31]),
    .X(_05954_));
 sky130_fd_sc_hd__buf_1 _20946_ (.A(_05954_),
    .X(_00837_));
 sky130_fd_sc_hd__and3_2 _20947_ (.A(\execute.io_reg_pc[0] ),
    .B(_05915_),
    .C(_05911_),
    .X(_05955_));
 sky130_fd_sc_hd__buf_1 _20948_ (.A(_05955_),
    .X(_00838_));
 sky130_fd_sc_hd__and3_2 _20949_ (.A(\execute.io_reg_pc[1] ),
    .B(_05915_),
    .C(_05911_),
    .X(_05956_));
 sky130_fd_sc_hd__buf_1 _20950_ (.A(_05956_),
    .X(_00839_));
 sky130_fd_sc_hd__and3_2 _20951_ (.A(\execute.io_reg_pc[2] ),
    .B(_05915_),
    .C(_05911_),
    .X(_05957_));
 sky130_fd_sc_hd__buf_1 _20952_ (.A(_05957_),
    .X(_00840_));
 sky130_fd_sc_hd__and3_2 _20953_ (.A(\execute.io_reg_pc[3] ),
    .B(_05915_),
    .C(_05911_),
    .X(_05958_));
 sky130_fd_sc_hd__buf_1 _20954_ (.A(_05958_),
    .X(_00841_));
 sky130_fd_sc_hd__and3_2 _20955_ (.A(\execute.io_reg_pc[4] ),
    .B(_05915_),
    .C(_05911_),
    .X(_05959_));
 sky130_fd_sc_hd__buf_1 _20956_ (.A(_05959_),
    .X(_00842_));
 sky130_fd_sc_hd__and3_2 _20957_ (.A(\execute.io_reg_pc[5] ),
    .B(_05915_),
    .C(_05911_),
    .X(_05960_));
 sky130_fd_sc_hd__buf_1 _20958_ (.A(_05960_),
    .X(_00843_));
 sky130_fd_sc_hd__buf_1 _20959_ (.A(_03582_),
    .X(_05961_));
 sky130_fd_sc_hd__and3_2 _20960_ (.A(\execute.io_reg_pc[6] ),
    .B(_05915_),
    .C(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__buf_1 _20961_ (.A(_05962_),
    .X(_00844_));
 sky130_fd_sc_hd__and3_2 _20962_ (.A(\execute.io_reg_pc[7] ),
    .B(_05915_),
    .C(_05961_),
    .X(_05963_));
 sky130_fd_sc_hd__buf_1 _20963_ (.A(_05963_),
    .X(_00845_));
 sky130_fd_sc_hd__and3_2 _20964_ (.A(\execute.io_reg_pc[8] ),
    .B(_05915_),
    .C(_05961_),
    .X(_05964_));
 sky130_fd_sc_hd__buf_1 _20965_ (.A(_05964_),
    .X(_00846_));
 sky130_fd_sc_hd__buf_1 _20966_ (.A(_05866_),
    .X(_05965_));
 sky130_fd_sc_hd__and3_2 _20967_ (.A(\execute.io_reg_pc[9] ),
    .B(_05965_),
    .C(_05961_),
    .X(_05966_));
 sky130_fd_sc_hd__buf_1 _20968_ (.A(_05966_),
    .X(_00847_));
 sky130_fd_sc_hd__and3_2 _20969_ (.A(\execute.io_reg_pc[10] ),
    .B(_05965_),
    .C(_05961_),
    .X(_05967_));
 sky130_fd_sc_hd__buf_1 _20970_ (.A(_05967_),
    .X(_00848_));
 sky130_fd_sc_hd__and3_2 _20971_ (.A(\execute.io_reg_pc[11] ),
    .B(_05965_),
    .C(_05961_),
    .X(_05968_));
 sky130_fd_sc_hd__buf_1 _20972_ (.A(_05968_),
    .X(_00849_));
 sky130_fd_sc_hd__and3_2 _20973_ (.A(\execute.io_reg_pc[12] ),
    .B(_05965_),
    .C(_05961_),
    .X(_05969_));
 sky130_fd_sc_hd__buf_1 _20974_ (.A(_05969_),
    .X(_00850_));
 sky130_fd_sc_hd__and3_2 _20975_ (.A(\execute.io_reg_pc[13] ),
    .B(_05965_),
    .C(_05961_),
    .X(_05970_));
 sky130_fd_sc_hd__buf_1 _20976_ (.A(_05970_),
    .X(_00851_));
 sky130_fd_sc_hd__and3_2 _20977_ (.A(\execute.io_reg_pc[14] ),
    .B(_05965_),
    .C(_05961_),
    .X(_05971_));
 sky130_fd_sc_hd__buf_1 _20978_ (.A(_05971_),
    .X(_00852_));
 sky130_fd_sc_hd__and3_2 _20979_ (.A(\execute.io_reg_pc[15] ),
    .B(_05965_),
    .C(_05961_),
    .X(_05972_));
 sky130_fd_sc_hd__buf_1 _20980_ (.A(_05972_),
    .X(_00853_));
 sky130_fd_sc_hd__buf_1 _20981_ (.A(_03582_),
    .X(_05973_));
 sky130_fd_sc_hd__and3_2 _20982_ (.A(\execute.io_reg_pc[16] ),
    .B(_05965_),
    .C(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__buf_1 _20983_ (.A(_05974_),
    .X(_00854_));
 sky130_fd_sc_hd__and3_2 _20984_ (.A(\execute.io_reg_pc[17] ),
    .B(_05965_),
    .C(_05973_),
    .X(_05975_));
 sky130_fd_sc_hd__buf_1 _20985_ (.A(_05975_),
    .X(_00855_));
 sky130_fd_sc_hd__and3_2 _20986_ (.A(\execute.io_reg_pc[18] ),
    .B(_05965_),
    .C(_05973_),
    .X(_05976_));
 sky130_fd_sc_hd__buf_1 _20987_ (.A(_05976_),
    .X(_00856_));
 sky130_fd_sc_hd__buf_1 _20988_ (.A(_05866_),
    .X(_05977_));
 sky130_fd_sc_hd__and3_2 _20989_ (.A(\execute.io_reg_pc[19] ),
    .B(_05977_),
    .C(_05973_),
    .X(_05978_));
 sky130_fd_sc_hd__buf_1 _20990_ (.A(_05978_),
    .X(_00857_));
 sky130_fd_sc_hd__and3_2 _20991_ (.A(\execute.io_reg_pc[20] ),
    .B(_05977_),
    .C(_05973_),
    .X(_05979_));
 sky130_fd_sc_hd__buf_1 _20992_ (.A(_05979_),
    .X(_00858_));
 sky130_fd_sc_hd__and3_2 _20993_ (.A(\execute.io_reg_pc[21] ),
    .B(_05977_),
    .C(_05973_),
    .X(_05980_));
 sky130_fd_sc_hd__buf_1 _20994_ (.A(_05980_),
    .X(_00859_));
 sky130_fd_sc_hd__and3_2 _20995_ (.A(\execute.io_reg_pc[22] ),
    .B(_05977_),
    .C(_05973_),
    .X(_05981_));
 sky130_fd_sc_hd__buf_1 _20996_ (.A(_05981_),
    .X(_00860_));
 sky130_fd_sc_hd__and3_2 _20997_ (.A(\execute.io_reg_pc[23] ),
    .B(_05977_),
    .C(_05973_),
    .X(_05982_));
 sky130_fd_sc_hd__buf_1 _20998_ (.A(_05982_),
    .X(_00861_));
 sky130_fd_sc_hd__and3_2 _20999_ (.A(\execute.io_reg_pc[24] ),
    .B(_05977_),
    .C(_05973_),
    .X(_05983_));
 sky130_fd_sc_hd__buf_1 _21000_ (.A(_05983_),
    .X(_00862_));
 sky130_fd_sc_hd__and3_2 _21001_ (.A(\execute.io_reg_pc[25] ),
    .B(_05977_),
    .C(_05973_),
    .X(_05984_));
 sky130_fd_sc_hd__buf_1 _21002_ (.A(_05984_),
    .X(_00863_));
 sky130_fd_sc_hd__buf_1 _21003_ (.A(_03582_),
    .X(_05985_));
 sky130_fd_sc_hd__and3_2 _21004_ (.A(\execute.io_reg_pc[26] ),
    .B(_05977_),
    .C(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__buf_1 _21005_ (.A(_05986_),
    .X(_00864_));
 sky130_fd_sc_hd__and3_2 _21006_ (.A(\execute.io_reg_pc[27] ),
    .B(_05977_),
    .C(_05985_),
    .X(_05987_));
 sky130_fd_sc_hd__buf_1 _21007_ (.A(_05987_),
    .X(_00865_));
 sky130_fd_sc_hd__and3_2 _21008_ (.A(\execute.io_reg_pc[28] ),
    .B(_05977_),
    .C(_05985_),
    .X(_05988_));
 sky130_fd_sc_hd__buf_1 _21009_ (.A(_05988_),
    .X(_00866_));
 sky130_fd_sc_hd__buf_1 _21010_ (.A(_05864_),
    .X(_05989_));
 sky130_fd_sc_hd__and3_2 _21011_ (.A(\execute.io_reg_pc[29] ),
    .B(_05989_),
    .C(_05985_),
    .X(_05990_));
 sky130_fd_sc_hd__buf_1 _21012_ (.A(_05990_),
    .X(_00867_));
 sky130_fd_sc_hd__and3_2 _21013_ (.A(\execute.io_reg_pc[30] ),
    .B(_05989_),
    .C(_05985_),
    .X(_05991_));
 sky130_fd_sc_hd__buf_1 _21014_ (.A(_05991_),
    .X(_00868_));
 sky130_fd_sc_hd__and3_2 _21015_ (.A(\execute.io_reg_pc[31] ),
    .B(_05989_),
    .C(_05985_),
    .X(_05992_));
 sky130_fd_sc_hd__buf_1 _21016_ (.A(_05992_),
    .X(_00869_));
 sky130_fd_sc_hd__and3_2 _21017_ (.A(_05949_),
    .B(_05945_),
    .C(\execute.io_mret_out ),
    .X(_05993_));
 sky130_fd_sc_hd__buf_1 _21018_ (.A(_05993_),
    .X(_00870_));
 sky130_fd_sc_hd__and3_2 _21019_ (.A(\execute.csr_read_data_out_reg[0] ),
    .B(_05989_),
    .C(_05985_),
    .X(_05994_));
 sky130_fd_sc_hd__buf_1 _21020_ (.A(_05994_),
    .X(_00871_));
 sky130_fd_sc_hd__and3_2 _21021_ (.A(\execute.csr_read_data_out_reg[1] ),
    .B(_05989_),
    .C(_05985_),
    .X(_05995_));
 sky130_fd_sc_hd__buf_1 _21022_ (.A(_05995_),
    .X(_00872_));
 sky130_fd_sc_hd__and3_2 _21023_ (.A(\execute.csr_read_data_out_reg[2] ),
    .B(_05989_),
    .C(_05985_),
    .X(_05996_));
 sky130_fd_sc_hd__buf_1 _21024_ (.A(_05996_),
    .X(_00873_));
 sky130_fd_sc_hd__and3_2 _21025_ (.A(\execute.csr_read_data_out_reg[3] ),
    .B(_05989_),
    .C(_05985_),
    .X(_05997_));
 sky130_fd_sc_hd__buf_1 _21026_ (.A(_05997_),
    .X(_00874_));
 sky130_fd_sc_hd__buf_1 _21027_ (.A(_03582_),
    .X(_05998_));
 sky130_fd_sc_hd__and3_2 _21028_ (.A(\execute.csr_read_data_out_reg[4] ),
    .B(_05989_),
    .C(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__buf_1 _21029_ (.A(_05999_),
    .X(_00875_));
 sky130_fd_sc_hd__and3_2 _21030_ (.A(\execute.csr_read_data_out_reg[5] ),
    .B(_05989_),
    .C(_05998_),
    .X(_06000_));
 sky130_fd_sc_hd__buf_1 _21031_ (.A(_06000_),
    .X(_00876_));
 sky130_fd_sc_hd__and3_2 _21032_ (.A(\execute.csr_read_data_out_reg[6] ),
    .B(_05989_),
    .C(_05998_),
    .X(_06001_));
 sky130_fd_sc_hd__buf_1 _21033_ (.A(_06001_),
    .X(_00877_));
 sky130_fd_sc_hd__buf_1 _21034_ (.A(_05864_),
    .X(_06002_));
 sky130_fd_sc_hd__and3_2 _21035_ (.A(\execute.csr_read_data_out_reg[7] ),
    .B(_06002_),
    .C(_05998_),
    .X(_06003_));
 sky130_fd_sc_hd__buf_1 _21036_ (.A(_06003_),
    .X(_00878_));
 sky130_fd_sc_hd__and3_2 _21037_ (.A(\execute.csr_read_data_out_reg[8] ),
    .B(_06002_),
    .C(_05998_),
    .X(_06004_));
 sky130_fd_sc_hd__buf_1 _21038_ (.A(_06004_),
    .X(_00879_));
 sky130_fd_sc_hd__and3_2 _21039_ (.A(\execute.csr_read_data_out_reg[9] ),
    .B(_06002_),
    .C(_05998_),
    .X(_06005_));
 sky130_fd_sc_hd__buf_1 _21040_ (.A(_06005_),
    .X(_00880_));
 sky130_fd_sc_hd__and3_2 _21041_ (.A(\execute.csr_read_data_out_reg[10] ),
    .B(_06002_),
    .C(_05998_),
    .X(_06006_));
 sky130_fd_sc_hd__buf_1 _21042_ (.A(_06006_),
    .X(_00881_));
 sky130_fd_sc_hd__and3_2 _21043_ (.A(\execute.csr_read_data_out_reg[11] ),
    .B(_06002_),
    .C(_05998_),
    .X(_06007_));
 sky130_fd_sc_hd__buf_1 _21044_ (.A(_06007_),
    .X(_00882_));
 sky130_fd_sc_hd__and3_2 _21045_ (.A(\execute.csr_read_data_out_reg[12] ),
    .B(_06002_),
    .C(_05998_),
    .X(_06008_));
 sky130_fd_sc_hd__buf_1 _21046_ (.A(_06008_),
    .X(_00883_));
 sky130_fd_sc_hd__and3_2 _21047_ (.A(\execute.csr_read_data_out_reg[13] ),
    .B(_06002_),
    .C(_05998_),
    .X(_06009_));
 sky130_fd_sc_hd__buf_1 _21048_ (.A(_06009_),
    .X(_00884_));
 sky130_fd_sc_hd__buf_1 _21049_ (.A(_09954_),
    .X(_06010_));
 sky130_fd_sc_hd__and3_2 _21050_ (.A(\execute.csr_read_data_out_reg[14] ),
    .B(_06002_),
    .C(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__buf_1 _21051_ (.A(_06011_),
    .X(_00885_));
 sky130_fd_sc_hd__and3_2 _21052_ (.A(\execute.csr_read_data_out_reg[15] ),
    .B(_06002_),
    .C(_06010_),
    .X(_06012_));
 sky130_fd_sc_hd__buf_1 _21053_ (.A(_06012_),
    .X(_00886_));
 sky130_fd_sc_hd__and3_2 _21054_ (.A(\execute.csr_read_data_out_reg[16] ),
    .B(_06002_),
    .C(_06010_),
    .X(_06013_));
 sky130_fd_sc_hd__buf_1 _21055_ (.A(_06013_),
    .X(_00887_));
 sky130_fd_sc_hd__buf_1 _21056_ (.A(_05864_),
    .X(_06014_));
 sky130_fd_sc_hd__and3_2 _21057_ (.A(\execute.csr_read_data_out_reg[17] ),
    .B(_06014_),
    .C(_06010_),
    .X(_06015_));
 sky130_fd_sc_hd__buf_1 _21058_ (.A(_06015_),
    .X(_00888_));
 sky130_fd_sc_hd__and3_2 _21059_ (.A(\execute.csr_read_data_out_reg[18] ),
    .B(_06014_),
    .C(_06010_),
    .X(_06016_));
 sky130_fd_sc_hd__buf_1 _21060_ (.A(_06016_),
    .X(_00889_));
 sky130_fd_sc_hd__and3_2 _21061_ (.A(\execute.csr_read_data_out_reg[19] ),
    .B(_06014_),
    .C(_06010_),
    .X(_06017_));
 sky130_fd_sc_hd__buf_1 _21062_ (.A(_06017_),
    .X(_00890_));
 sky130_fd_sc_hd__and3_2 _21063_ (.A(\execute.csr_read_data_out_reg[20] ),
    .B(_06014_),
    .C(_06010_),
    .X(_06018_));
 sky130_fd_sc_hd__buf_1 _21064_ (.A(_06018_),
    .X(_00891_));
 sky130_fd_sc_hd__and3_2 _21065_ (.A(\execute.csr_read_data_out_reg[21] ),
    .B(_06014_),
    .C(_06010_),
    .X(_06019_));
 sky130_fd_sc_hd__buf_1 _21066_ (.A(_06019_),
    .X(_00892_));
 sky130_fd_sc_hd__and3_2 _21067_ (.A(\execute.csr_read_data_out_reg[22] ),
    .B(_06014_),
    .C(_06010_),
    .X(_06020_));
 sky130_fd_sc_hd__buf_1 _21068_ (.A(_06020_),
    .X(_00893_));
 sky130_fd_sc_hd__and3_2 _21069_ (.A(\execute.csr_read_data_out_reg[23] ),
    .B(_06014_),
    .C(_06010_),
    .X(_06021_));
 sky130_fd_sc_hd__buf_1 _21070_ (.A(_06021_),
    .X(_00894_));
 sky130_fd_sc_hd__and3_2 _21071_ (.A(\execute.csr_read_data_out_reg[24] ),
    .B(_06014_),
    .C(_03583_),
    .X(_06022_));
 sky130_fd_sc_hd__buf_1 _21072_ (.A(_06022_),
    .X(_00895_));
 sky130_fd_sc_hd__and3_2 _21073_ (.A(\execute.csr_read_data_out_reg[25] ),
    .B(_06014_),
    .C(_03583_),
    .X(_06023_));
 sky130_fd_sc_hd__buf_1 _21074_ (.A(_06023_),
    .X(_00896_));
 sky130_fd_sc_hd__and3_2 _21075_ (.A(\execute.csr_read_data_out_reg[26] ),
    .B(_06014_),
    .C(_03583_),
    .X(_06024_));
 sky130_fd_sc_hd__buf_1 _21076_ (.A(_06024_),
    .X(_00897_));
 sky130_fd_sc_hd__buf_1 _21077_ (.A(_05864_),
    .X(_06025_));
 sky130_fd_sc_hd__and3_2 _21078_ (.A(\execute.csr_read_data_out_reg[27] ),
    .B(_06025_),
    .C(_03583_),
    .X(_06026_));
 sky130_fd_sc_hd__buf_1 _21079_ (.A(_06026_),
    .X(_00898_));
 sky130_fd_sc_hd__and3_2 _21080_ (.A(\execute.csr_read_data_out_reg[28] ),
    .B(_06025_),
    .C(_03583_),
    .X(_06027_));
 sky130_fd_sc_hd__buf_1 _21081_ (.A(_06027_),
    .X(_00899_));
 sky130_fd_sc_hd__and3_2 _21082_ (.A(\execute.csr_read_data_out_reg[29] ),
    .B(_06025_),
    .C(_03583_),
    .X(_06028_));
 sky130_fd_sc_hd__buf_1 _21083_ (.A(_06028_),
    .X(_00900_));
 sky130_fd_sc_hd__and3_2 _21084_ (.A(\execute.csr_read_data_out_reg[30] ),
    .B(_06025_),
    .C(_03583_),
    .X(_06029_));
 sky130_fd_sc_hd__buf_1 _21085_ (.A(_06029_),
    .X(_00901_));
 sky130_fd_sc_hd__and3_2 _21086_ (.A(\execute.csr_read_data_out_reg[31] ),
    .B(_06025_),
    .C(_03583_),
    .X(_06030_));
 sky130_fd_sc_hd__buf_1 _21087_ (.A(_06030_),
    .X(_00902_));
 sky130_fd_sc_hd__a21oi_2 _21088_ (.A1(_09921_),
    .A2(io_memory_read),
    .B1(_09922_),
    .Y(_06031_));
 sky130_fd_sc_hd__buf_1 _21089_ (.A(_10971_),
    .X(_06032_));
 sky130_fd_sc_hd__nor2_2 _21090_ (.A(_10576_),
    .B(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__and4bb_2 _21091_ (.A_N(\execute.io_wfi_out ),
    .B_N(_09925_),
    .C(_06031_),
    .D(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__buf_1 _21092_ (.A(_06034_),
    .X(_00903_));
 sky130_fd_sc_hd__a31o_2 _21093_ (.A1(\csr.mtie ),
    .A2(\csr.ie ),
    .A3(\csr.mtip ),
    .B1(_09924_),
    .X(_06035_));
 sky130_fd_sc_hd__and3_2 _21094_ (.A(_10019_),
    .B(_06035_),
    .C(_06025_),
    .X(_06036_));
 sky130_fd_sc_hd__buf_1 _21095_ (.A(_06036_),
    .X(_00904_));
 sky130_fd_sc_hd__buf_1 _21096_ (.A(\csr.io_trapped ),
    .X(_06037_));
 sky130_fd_sc_hd__buf_1 _21097_ (.A(_06037_),
    .X(_06038_));
 sky130_fd_sc_hd__buf_1 _21098_ (.A(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__buf_1 _21099_ (.A(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__buf_1 _21100_ (.A(_10970_),
    .X(_06041_));
 sky130_fd_sc_hd__nor4_2 _21101_ (.A(_06040_),
    .B(_06041_),
    .C(_10577_),
    .D(_09926_),
    .Y(_00905_));
 sky130_fd_sc_hd__and4b_2 _21102_ (.A_N(\execute.exception_out_reg ),
    .B(_06033_),
    .C(_09921_),
    .D(io_memory_read),
    .X(_06042_));
 sky130_fd_sc_hd__a31o_2 _21103_ (.A1(_05856_),
    .A2(_06035_),
    .A3(_05858_),
    .B1(_06042_),
    .X(_00906_));
 sky130_fd_sc_hd__o21ai_2 _21104_ (.A1(io_memory_address[0]),
    .A2(io_memory_address[1]),
    .B1(\execute.io_mem_memwrite ),
    .Y(_06043_));
 sky130_fd_sc_hd__nor2_2 _21105_ (.A(io_memory_read),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__o311a_2 _21106_ (.A1(\execute.exception_out_reg ),
    .A2(_06044_),
    .A3(_06035_),
    .B1(_05856_),
    .C1(_05858_),
    .X(_00907_));
 sky130_fd_sc_hd__and3_2 _21107_ (.A(_05949_),
    .B(_05945_),
    .C(\execute.csr_write_data_out_reg[0] ),
    .X(_06045_));
 sky130_fd_sc_hd__buf_1 _21108_ (.A(_06045_),
    .X(_00908_));
 sky130_fd_sc_hd__buf_1 _21109_ (.A(_09955_),
    .X(_06046_));
 sky130_fd_sc_hd__and3_2 _21110_ (.A(_05949_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[1] ),
    .X(_06047_));
 sky130_fd_sc_hd__buf_1 _21111_ (.A(_06047_),
    .X(_00909_));
 sky130_fd_sc_hd__and3_2 _21112_ (.A(_05949_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[2] ),
    .X(_06048_));
 sky130_fd_sc_hd__buf_1 _21113_ (.A(_06048_),
    .X(_00910_));
 sky130_fd_sc_hd__and3_2 _21114_ (.A(_05949_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[3] ),
    .X(_06049_));
 sky130_fd_sc_hd__buf_1 _21115_ (.A(_06049_),
    .X(_00911_));
 sky130_fd_sc_hd__buf_1 _21116_ (.A(_05857_),
    .X(_06050_));
 sky130_fd_sc_hd__and3_2 _21117_ (.A(_06050_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[4] ),
    .X(_06051_));
 sky130_fd_sc_hd__buf_1 _21118_ (.A(_06051_),
    .X(_00912_));
 sky130_fd_sc_hd__and3_2 _21119_ (.A(_06050_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[5] ),
    .X(_06052_));
 sky130_fd_sc_hd__buf_1 _21120_ (.A(_06052_),
    .X(_00913_));
 sky130_fd_sc_hd__and3_2 _21121_ (.A(_06050_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[6] ),
    .X(_06053_));
 sky130_fd_sc_hd__buf_1 _21122_ (.A(_06053_),
    .X(_00914_));
 sky130_fd_sc_hd__and3_2 _21123_ (.A(_06050_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[7] ),
    .X(_06054_));
 sky130_fd_sc_hd__buf_1 _21124_ (.A(_06054_),
    .X(_00915_));
 sky130_fd_sc_hd__and3_2 _21125_ (.A(_06050_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[8] ),
    .X(_06055_));
 sky130_fd_sc_hd__buf_1 _21126_ (.A(_06055_),
    .X(_00916_));
 sky130_fd_sc_hd__and3_2 _21127_ (.A(_06050_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[9] ),
    .X(_06056_));
 sky130_fd_sc_hd__buf_1 _21128_ (.A(_06056_),
    .X(_00917_));
 sky130_fd_sc_hd__and3_2 _21129_ (.A(_06050_),
    .B(_06046_),
    .C(\execute.csr_write_data_out_reg[10] ),
    .X(_06057_));
 sky130_fd_sc_hd__buf_1 _21130_ (.A(_06057_),
    .X(_00918_));
 sky130_fd_sc_hd__buf_1 _21131_ (.A(_09955_),
    .X(_06058_));
 sky130_fd_sc_hd__and3_2 _21132_ (.A(_06050_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[11] ),
    .X(_06059_));
 sky130_fd_sc_hd__buf_1 _21133_ (.A(_06059_),
    .X(_00919_));
 sky130_fd_sc_hd__and3_2 _21134_ (.A(_06050_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[12] ),
    .X(_06060_));
 sky130_fd_sc_hd__buf_1 _21135_ (.A(_06060_),
    .X(_00920_));
 sky130_fd_sc_hd__and3_2 _21136_ (.A(_06050_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[13] ),
    .X(_06061_));
 sky130_fd_sc_hd__buf_1 _21137_ (.A(_06061_),
    .X(_00921_));
 sky130_fd_sc_hd__buf_1 _21138_ (.A(_05866_),
    .X(_06062_));
 sky130_fd_sc_hd__and3_2 _21139_ (.A(_06062_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[14] ),
    .X(_06063_));
 sky130_fd_sc_hd__buf_1 _21140_ (.A(_06063_),
    .X(_00922_));
 sky130_fd_sc_hd__and3_2 _21141_ (.A(_06062_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[15] ),
    .X(_06064_));
 sky130_fd_sc_hd__buf_1 _21142_ (.A(_06064_),
    .X(_00923_));
 sky130_fd_sc_hd__and3_2 _21143_ (.A(_06062_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[16] ),
    .X(_06065_));
 sky130_fd_sc_hd__buf_1 _21144_ (.A(_06065_),
    .X(_00924_));
 sky130_fd_sc_hd__and3_2 _21145_ (.A(_06062_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[17] ),
    .X(_06066_));
 sky130_fd_sc_hd__buf_1 _21146_ (.A(_06066_),
    .X(_00925_));
 sky130_fd_sc_hd__and3_2 _21147_ (.A(_06062_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[18] ),
    .X(_06067_));
 sky130_fd_sc_hd__buf_1 _21148_ (.A(_06067_),
    .X(_00926_));
 sky130_fd_sc_hd__and3_2 _21149_ (.A(_06062_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[19] ),
    .X(_06068_));
 sky130_fd_sc_hd__buf_1 _21150_ (.A(_06068_),
    .X(_00927_));
 sky130_fd_sc_hd__and3_2 _21151_ (.A(_06062_),
    .B(_06058_),
    .C(\execute.csr_write_data_out_reg[20] ),
    .X(_06069_));
 sky130_fd_sc_hd__buf_1 _21152_ (.A(_06069_),
    .X(_00928_));
 sky130_fd_sc_hd__buf_1 _21153_ (.A(_09955_),
    .X(_06070_));
 sky130_fd_sc_hd__and3_2 _21154_ (.A(_06062_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[21] ),
    .X(_06071_));
 sky130_fd_sc_hd__buf_1 _21155_ (.A(_06071_),
    .X(_00929_));
 sky130_fd_sc_hd__and3_2 _21156_ (.A(_06062_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[22] ),
    .X(_06072_));
 sky130_fd_sc_hd__buf_1 _21157_ (.A(_06072_),
    .X(_00930_));
 sky130_fd_sc_hd__and3_2 _21158_ (.A(_06062_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[23] ),
    .X(_06073_));
 sky130_fd_sc_hd__buf_1 _21159_ (.A(_06073_),
    .X(_00931_));
 sky130_fd_sc_hd__buf_1 _21160_ (.A(_05866_),
    .X(_06074_));
 sky130_fd_sc_hd__and3_2 _21161_ (.A(_06074_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[24] ),
    .X(_06075_));
 sky130_fd_sc_hd__buf_1 _21162_ (.A(_06075_),
    .X(_00932_));
 sky130_fd_sc_hd__and3_2 _21163_ (.A(_06074_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[25] ),
    .X(_06076_));
 sky130_fd_sc_hd__buf_1 _21164_ (.A(_06076_),
    .X(_00933_));
 sky130_fd_sc_hd__and3_2 _21165_ (.A(_06074_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[26] ),
    .X(_06077_));
 sky130_fd_sc_hd__buf_1 _21166_ (.A(_06077_),
    .X(_00934_));
 sky130_fd_sc_hd__and3_2 _21167_ (.A(_06074_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[27] ),
    .X(_06078_));
 sky130_fd_sc_hd__buf_1 _21168_ (.A(_06078_),
    .X(_00935_));
 sky130_fd_sc_hd__and3_2 _21169_ (.A(_06074_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[28] ),
    .X(_06079_));
 sky130_fd_sc_hd__buf_1 _21170_ (.A(_06079_),
    .X(_00936_));
 sky130_fd_sc_hd__and3_2 _21171_ (.A(_06074_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[29] ),
    .X(_06080_));
 sky130_fd_sc_hd__buf_1 _21172_ (.A(_06080_),
    .X(_00937_));
 sky130_fd_sc_hd__and3_2 _21173_ (.A(_06074_),
    .B(_06070_),
    .C(\execute.csr_write_data_out_reg[30] ),
    .X(_06081_));
 sky130_fd_sc_hd__buf_1 _21174_ (.A(_06081_),
    .X(_00938_));
 sky130_fd_sc_hd__buf_1 _21175_ (.A(_09955_),
    .X(_06082_));
 sky130_fd_sc_hd__and3_2 _21176_ (.A(_06074_),
    .B(_06082_),
    .C(\execute.csr_write_data_out_reg[31] ),
    .X(_06083_));
 sky130_fd_sc_hd__buf_1 _21177_ (.A(_06083_),
    .X(_00939_));
 sky130_fd_sc_hd__and3_2 _21178_ (.A(_06074_),
    .B(_06082_),
    .C(\execute.csr_write_address_out_reg[0] ),
    .X(_06084_));
 sky130_fd_sc_hd__buf_1 _21179_ (.A(_06084_),
    .X(_00940_));
 sky130_fd_sc_hd__and3_2 _21180_ (.A(_06074_),
    .B(_06082_),
    .C(\execute.csr_write_address_out_reg[1] ),
    .X(_06085_));
 sky130_fd_sc_hd__buf_1 _21181_ (.A(_06085_),
    .X(_00941_));
 sky130_fd_sc_hd__buf_1 _21182_ (.A(_05866_),
    .X(_06086_));
 sky130_fd_sc_hd__and3_2 _21183_ (.A(_06086_),
    .B(_06082_),
    .C(\execute.csr_write_address_out_reg[2] ),
    .X(_06087_));
 sky130_fd_sc_hd__buf_1 _21184_ (.A(_06087_),
    .X(_00942_));
 sky130_fd_sc_hd__and3_2 _21185_ (.A(_06086_),
    .B(_06082_),
    .C(\execute.csr_write_address_out_reg[3] ),
    .X(_06088_));
 sky130_fd_sc_hd__buf_1 _21186_ (.A(_06088_),
    .X(_00943_));
 sky130_fd_sc_hd__and3_2 _21187_ (.A(_06086_),
    .B(_06082_),
    .C(\execute.csr_write_address_out_reg[4] ),
    .X(_06089_));
 sky130_fd_sc_hd__buf_1 _21188_ (.A(_06089_),
    .X(_00944_));
 sky130_fd_sc_hd__and3_2 _21189_ (.A(_06086_),
    .B(_06082_),
    .C(\execute.csr_write_address_out_reg[5] ),
    .X(_06090_));
 sky130_fd_sc_hd__buf_1 _21190_ (.A(_06090_),
    .X(_00945_));
 sky130_fd_sc_hd__and3_2 _21191_ (.A(_06086_),
    .B(_06082_),
    .C(\execute.csr_write_address_out_reg[6] ),
    .X(_06091_));
 sky130_fd_sc_hd__buf_1 _21192_ (.A(_06091_),
    .X(_00946_));
 sky130_fd_sc_hd__and3_2 _21193_ (.A(_06086_),
    .B(_06082_),
    .C(\execute.csr_write_address_out_reg[7] ),
    .X(_06092_));
 sky130_fd_sc_hd__buf_1 _21194_ (.A(_06092_),
    .X(_00947_));
 sky130_fd_sc_hd__and3_2 _21195_ (.A(_06086_),
    .B(_06082_),
    .C(\execute.csr_write_address_out_reg[8] ),
    .X(_06093_));
 sky130_fd_sc_hd__buf_1 _21196_ (.A(_06093_),
    .X(_00948_));
 sky130_fd_sc_hd__and3_2 _21197_ (.A(_06086_),
    .B(_05868_),
    .C(\execute.csr_write_address_out_reg[9] ),
    .X(_06094_));
 sky130_fd_sc_hd__buf_1 _21198_ (.A(_06094_),
    .X(_00949_));
 sky130_fd_sc_hd__and3_2 _21199_ (.A(_06086_),
    .B(_05868_),
    .C(\execute.csr_write_address_out_reg[10] ),
    .X(_06095_));
 sky130_fd_sc_hd__buf_1 _21200_ (.A(_06095_),
    .X(_00950_));
 sky130_fd_sc_hd__and3_2 _21201_ (.A(_06086_),
    .B(_05868_),
    .C(\execute.csr_write_address_out_reg[11] ),
    .X(_06096_));
 sky130_fd_sc_hd__buf_1 _21202_ (.A(_06096_),
    .X(_00951_));
 sky130_fd_sc_hd__and3_2 _21203_ (.A(_05867_),
    .B(_05868_),
    .C(\execute.csr_write_enable_out_reg ),
    .X(_06097_));
 sky130_fd_sc_hd__buf_1 _21204_ (.A(_06097_),
    .X(_00952_));
 sky130_fd_sc_hd__and2_2 _21205_ (.A(\decode.id_ex_ex_rd_reg[0] ),
    .B(_05214_),
    .X(_06098_));
 sky130_fd_sc_hd__buf_1 _21206_ (.A(_06098_),
    .X(_00953_));
 sky130_fd_sc_hd__nor2_2 _21207_ (.A(_10613_),
    .B(_05671_),
    .Y(_00954_));
 sky130_fd_sc_hd__and2_2 _21208_ (.A(\decode.id_ex_ex_rd_reg[2] ),
    .B(_05214_),
    .X(_06099_));
 sky130_fd_sc_hd__buf_1 _21209_ (.A(_06099_),
    .X(_00955_));
 sky130_fd_sc_hd__nor2_2 _21210_ (.A(_10596_),
    .B(_05671_),
    .Y(_00956_));
 sky130_fd_sc_hd__and2_2 _21211_ (.A(\decode.id_ex_ex_rd_reg[4] ),
    .B(_05214_),
    .X(_06100_));
 sky130_fd_sc_hd__buf_1 _21212_ (.A(_06100_),
    .X(_00957_));
 sky130_fd_sc_hd__buf_1 _21213_ (.A(_10820_),
    .X(_06101_));
 sky130_fd_sc_hd__mux2_2 _21214_ (.A0(\fetch.bht.bhtTable_tag[8][0] ),
    .A1(_06101_),
    .S(_09912_),
    .X(_06102_));
 sky130_fd_sc_hd__buf_1 _21215_ (.A(_06102_),
    .X(_00958_));
 sky130_fd_sc_hd__buf_1 _21216_ (.A(_10821_),
    .X(_06103_));
 sky130_fd_sc_hd__mux2_2 _21217_ (.A0(\fetch.bht.bhtTable_tag[8][1] ),
    .A1(_06103_),
    .S(_09912_),
    .X(_06104_));
 sky130_fd_sc_hd__buf_1 _21218_ (.A(_06104_),
    .X(_00959_));
 sky130_fd_sc_hd__buf_1 _21219_ (.A(_10881_),
    .X(_06105_));
 sky130_fd_sc_hd__mux2_2 _21220_ (.A0(\fetch.bht.bhtTable_tag[8][2] ),
    .A1(_06105_),
    .S(_09912_),
    .X(_06106_));
 sky130_fd_sc_hd__buf_1 _21221_ (.A(_06106_),
    .X(_00960_));
 sky130_fd_sc_hd__buf_1 _21222_ (.A(_10817_),
    .X(_06107_));
 sky130_fd_sc_hd__mux2_2 _21223_ (.A0(\fetch.bht.bhtTable_tag[8][3] ),
    .A1(_06107_),
    .S(_09912_),
    .X(_06108_));
 sky130_fd_sc_hd__buf_1 _21224_ (.A(_06108_),
    .X(_00961_));
 sky130_fd_sc_hd__buf_1 _21225_ (.A(_10878_),
    .X(_06109_));
 sky130_fd_sc_hd__mux2_2 _21226_ (.A0(\fetch.bht.bhtTable_tag[8][4] ),
    .A1(_06109_),
    .S(_09912_),
    .X(_06110_));
 sky130_fd_sc_hd__buf_1 _21227_ (.A(_06110_),
    .X(_00962_));
 sky130_fd_sc_hd__buf_1 _21228_ (.A(_10812_),
    .X(_06111_));
 sky130_fd_sc_hd__mux2_2 _21229_ (.A0(\fetch.bht.bhtTable_tag[8][5] ),
    .A1(_06111_),
    .S(_09912_),
    .X(_06112_));
 sky130_fd_sc_hd__buf_1 _21230_ (.A(_06112_),
    .X(_00963_));
 sky130_fd_sc_hd__buf_1 _21231_ (.A(\csr.io_mem_pc[12] ),
    .X(_06113_));
 sky130_fd_sc_hd__mux2_2 _21232_ (.A0(\fetch.bht.bhtTable_tag[8][6] ),
    .A1(_06113_),
    .S(_09912_),
    .X(_06114_));
 sky130_fd_sc_hd__buf_1 _21233_ (.A(_06114_),
    .X(_00964_));
 sky130_fd_sc_hd__buf_1 _21234_ (.A(_10871_),
    .X(_06115_));
 sky130_fd_sc_hd__mux2_2 _21235_ (.A0(\fetch.bht.bhtTable_tag[8][7] ),
    .A1(_06115_),
    .S(_09912_),
    .X(_06116_));
 sky130_fd_sc_hd__buf_1 _21236_ (.A(_06116_),
    .X(_00965_));
 sky130_fd_sc_hd__buf_1 _21237_ (.A(_10872_),
    .X(_06117_));
 sky130_fd_sc_hd__mux2_2 _21238_ (.A0(\fetch.bht.bhtTable_tag[8][8] ),
    .A1(_06117_),
    .S(_09912_),
    .X(_06118_));
 sky130_fd_sc_hd__buf_1 _21239_ (.A(_06118_),
    .X(_00966_));
 sky130_fd_sc_hd__buf_1 _21240_ (.A(_10807_),
    .X(_06119_));
 sky130_fd_sc_hd__buf_1 _21241_ (.A(_09910_),
    .X(_06120_));
 sky130_fd_sc_hd__mux2_2 _21242_ (.A0(\fetch.bht.bhtTable_tag[8][9] ),
    .A1(_06119_),
    .S(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__buf_1 _21243_ (.A(_06121_),
    .X(_00967_));
 sky130_fd_sc_hd__buf_1 _21244_ (.A(_10868_),
    .X(_06122_));
 sky130_fd_sc_hd__mux2_2 _21245_ (.A0(\fetch.bht.bhtTable_tag[8][10] ),
    .A1(_06122_),
    .S(_06120_),
    .X(_06123_));
 sky130_fd_sc_hd__buf_1 _21246_ (.A(_06123_),
    .X(_00968_));
 sky130_fd_sc_hd__buf_1 _21247_ (.A(_10803_),
    .X(_06124_));
 sky130_fd_sc_hd__mux2_2 _21248_ (.A0(\fetch.bht.bhtTable_tag[8][11] ),
    .A1(_06124_),
    .S(_06120_),
    .X(_06125_));
 sky130_fd_sc_hd__buf_1 _21249_ (.A(_06125_),
    .X(_00969_));
 sky130_fd_sc_hd__buf_1 _21250_ (.A(\csr.io_mem_pc[18] ),
    .X(_06126_));
 sky130_fd_sc_hd__mux2_2 _21251_ (.A0(\fetch.bht.bhtTable_tag[8][12] ),
    .A1(_06126_),
    .S(_06120_),
    .X(_06127_));
 sky130_fd_sc_hd__buf_1 _21252_ (.A(_06127_),
    .X(_00970_));
 sky130_fd_sc_hd__buf_1 _21253_ (.A(_10800_),
    .X(_06128_));
 sky130_fd_sc_hd__mux2_2 _21254_ (.A0(\fetch.bht.bhtTable_tag[8][13] ),
    .A1(_06128_),
    .S(_06120_),
    .X(_06129_));
 sky130_fd_sc_hd__buf_1 _21255_ (.A(_06129_),
    .X(_00971_));
 sky130_fd_sc_hd__buf_1 _21256_ (.A(_10795_),
    .X(_06130_));
 sky130_fd_sc_hd__mux2_2 _21257_ (.A0(\fetch.bht.bhtTable_tag[8][14] ),
    .A1(_06130_),
    .S(_06120_),
    .X(_06131_));
 sky130_fd_sc_hd__buf_1 _21258_ (.A(_06131_),
    .X(_00972_));
 sky130_fd_sc_hd__buf_1 _21259_ (.A(\csr.io_mem_pc[21] ),
    .X(_06132_));
 sky130_fd_sc_hd__mux2_2 _21260_ (.A0(\fetch.bht.bhtTable_tag[8][15] ),
    .A1(_06132_),
    .S(_06120_),
    .X(_06133_));
 sky130_fd_sc_hd__buf_1 _21261_ (.A(_06133_),
    .X(_00973_));
 sky130_fd_sc_hd__buf_1 _21262_ (.A(_10787_),
    .X(_06134_));
 sky130_fd_sc_hd__mux2_2 _21263_ (.A0(\fetch.bht.bhtTable_tag[8][16] ),
    .A1(_06134_),
    .S(_06120_),
    .X(_06135_));
 sky130_fd_sc_hd__buf_1 _21264_ (.A(_06135_),
    .X(_00974_));
 sky130_fd_sc_hd__buf_1 _21265_ (.A(\csr.io_mem_pc[23] ),
    .X(_06136_));
 sky130_fd_sc_hd__mux2_2 _21266_ (.A0(\fetch.bht.bhtTable_tag[8][17] ),
    .A1(_06136_),
    .S(_06120_),
    .X(_06137_));
 sky130_fd_sc_hd__buf_1 _21267_ (.A(_06137_),
    .X(_00975_));
 sky130_fd_sc_hd__buf_1 _21268_ (.A(_10772_),
    .X(_06138_));
 sky130_fd_sc_hd__mux2_2 _21269_ (.A0(\fetch.bht.bhtTable_tag[8][18] ),
    .A1(_06138_),
    .S(_06120_),
    .X(_06139_));
 sky130_fd_sc_hd__buf_1 _21270_ (.A(_06139_),
    .X(_00976_));
 sky130_fd_sc_hd__buf_1 _21271_ (.A(_10773_),
    .X(_06140_));
 sky130_fd_sc_hd__buf_1 _21272_ (.A(_09910_),
    .X(_06141_));
 sky130_fd_sc_hd__mux2_2 _21273_ (.A0(\fetch.bht.bhtTable_tag[8][19] ),
    .A1(_06140_),
    .S(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__buf_1 _21274_ (.A(_06142_),
    .X(_00977_));
 sky130_fd_sc_hd__buf_1 _21275_ (.A(_10760_),
    .X(_06143_));
 sky130_fd_sc_hd__mux2_2 _21276_ (.A0(\fetch.bht.bhtTable_tag[8][20] ),
    .A1(_06143_),
    .S(_06141_),
    .X(_06144_));
 sky130_fd_sc_hd__buf_1 _21277_ (.A(_06144_),
    .X(_00978_));
 sky130_fd_sc_hd__buf_1 _21278_ (.A(_10759_),
    .X(_06145_));
 sky130_fd_sc_hd__mux2_2 _21279_ (.A0(\fetch.bht.bhtTable_tag[8][21] ),
    .A1(_06145_),
    .S(_06141_),
    .X(_06146_));
 sky130_fd_sc_hd__buf_1 _21280_ (.A(_06146_),
    .X(_00979_));
 sky130_fd_sc_hd__buf_1 _21281_ (.A(_10771_),
    .X(_06147_));
 sky130_fd_sc_hd__mux2_2 _21282_ (.A0(\fetch.bht.bhtTable_tag[8][22] ),
    .A1(_06147_),
    .S(_06141_),
    .X(_06148_));
 sky130_fd_sc_hd__buf_1 _21283_ (.A(_06148_),
    .X(_00980_));
 sky130_fd_sc_hd__buf_1 _21284_ (.A(\csr.io_mem_pc[29] ),
    .X(_06149_));
 sky130_fd_sc_hd__mux2_2 _21285_ (.A0(\fetch.bht.bhtTable_tag[8][23] ),
    .A1(_06149_),
    .S(_06141_),
    .X(_06150_));
 sky130_fd_sc_hd__buf_1 _21286_ (.A(_06150_),
    .X(_00981_));
 sky130_fd_sc_hd__buf_1 _21287_ (.A(_10777_),
    .X(_06151_));
 sky130_fd_sc_hd__mux2_2 _21288_ (.A0(\fetch.bht.bhtTable_tag[8][24] ),
    .A1(_06151_),
    .S(_06141_),
    .X(_06152_));
 sky130_fd_sc_hd__buf_1 _21289_ (.A(_06152_),
    .X(_00982_));
 sky130_fd_sc_hd__buf_1 _21290_ (.A(\csr.io_mem_pc[31] ),
    .X(_06153_));
 sky130_fd_sc_hd__mux2_2 _21291_ (.A0(\fetch.bht.bhtTable_tag[8][25] ),
    .A1(_06153_),
    .S(_06141_),
    .X(_06154_));
 sky130_fd_sc_hd__buf_1 _21292_ (.A(_06154_),
    .X(_00983_));
 sky130_fd_sc_hd__and3_2 _21293_ (.A(_09885_),
    .B(_09890_),
    .C(_09917_),
    .X(_06155_));
 sky130_fd_sc_hd__buf_1 _21294_ (.A(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__buf_1 _21295_ (.A(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__mux2_2 _21296_ (.A0(\fetch.bht.bhtTable_tag[1][0] ),
    .A1(_06101_),
    .S(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__buf_1 _21297_ (.A(_06158_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_2 _21298_ (.A0(\fetch.bht.bhtTable_tag[1][1] ),
    .A1(_10821_),
    .S(_06157_),
    .X(_06159_));
 sky130_fd_sc_hd__buf_1 _21299_ (.A(_06159_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_2 _21300_ (.A0(\fetch.bht.bhtTable_tag[1][2] ),
    .A1(_10881_),
    .S(_06157_),
    .X(_06160_));
 sky130_fd_sc_hd__buf_1 _21301_ (.A(_06160_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_2 _21302_ (.A0(\fetch.bht.bhtTable_tag[1][3] ),
    .A1(_10817_),
    .S(_06157_),
    .X(_06161_));
 sky130_fd_sc_hd__buf_1 _21303_ (.A(_06161_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_2 _21304_ (.A0(\fetch.bht.bhtTable_tag[1][4] ),
    .A1(_10878_),
    .S(_06157_),
    .X(_06162_));
 sky130_fd_sc_hd__buf_1 _21305_ (.A(_06162_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_2 _21306_ (.A0(\fetch.bht.bhtTable_tag[1][5] ),
    .A1(_10812_),
    .S(_06157_),
    .X(_06163_));
 sky130_fd_sc_hd__buf_1 _21307_ (.A(_06163_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_2 _21308_ (.A0(\fetch.bht.bhtTable_tag[1][6] ),
    .A1(\csr.io_mem_pc[12] ),
    .S(_06157_),
    .X(_06164_));
 sky130_fd_sc_hd__buf_1 _21309_ (.A(_06164_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_2 _21310_ (.A0(\fetch.bht.bhtTable_tag[1][7] ),
    .A1(_10871_),
    .S(_06157_),
    .X(_06165_));
 sky130_fd_sc_hd__buf_1 _21311_ (.A(_06165_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_2 _21312_ (.A0(\fetch.bht.bhtTable_tag[1][8] ),
    .A1(_10872_),
    .S(_06157_),
    .X(_06166_));
 sky130_fd_sc_hd__buf_1 _21313_ (.A(_06166_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_2 _21314_ (.A0(\fetch.bht.bhtTable_tag[1][9] ),
    .A1(_10807_),
    .S(_06157_),
    .X(_06167_));
 sky130_fd_sc_hd__buf_1 _21315_ (.A(_06167_),
    .X(_00993_));
 sky130_fd_sc_hd__buf_1 _21316_ (.A(_06156_),
    .X(_06168_));
 sky130_fd_sc_hd__mux2_2 _21317_ (.A0(\fetch.bht.bhtTable_tag[1][10] ),
    .A1(_10868_),
    .S(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__buf_1 _21318_ (.A(_06169_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_2 _21319_ (.A0(\fetch.bht.bhtTable_tag[1][11] ),
    .A1(_10803_),
    .S(_06168_),
    .X(_06170_));
 sky130_fd_sc_hd__buf_1 _21320_ (.A(_06170_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_2 _21321_ (.A0(\fetch.bht.bhtTable_tag[1][12] ),
    .A1(\csr.io_mem_pc[18] ),
    .S(_06168_),
    .X(_06171_));
 sky130_fd_sc_hd__buf_1 _21322_ (.A(_06171_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_2 _21323_ (.A0(\fetch.bht.bhtTable_tag[1][13] ),
    .A1(_10800_),
    .S(_06168_),
    .X(_06172_));
 sky130_fd_sc_hd__buf_1 _21324_ (.A(_06172_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_2 _21325_ (.A0(\fetch.bht.bhtTable_tag[1][14] ),
    .A1(_10795_),
    .S(_06168_),
    .X(_06173_));
 sky130_fd_sc_hd__buf_1 _21326_ (.A(_06173_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_2 _21327_ (.A0(\fetch.bht.bhtTable_tag[1][15] ),
    .A1(\csr.io_mem_pc[21] ),
    .S(_06168_),
    .X(_06174_));
 sky130_fd_sc_hd__buf_1 _21328_ (.A(_06174_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_2 _21329_ (.A0(\fetch.bht.bhtTable_tag[1][16] ),
    .A1(_10787_),
    .S(_06168_),
    .X(_06175_));
 sky130_fd_sc_hd__buf_1 _21330_ (.A(_06175_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_2 _21331_ (.A0(\fetch.bht.bhtTable_tag[1][17] ),
    .A1(\csr.io_mem_pc[23] ),
    .S(_06168_),
    .X(_06176_));
 sky130_fd_sc_hd__buf_1 _21332_ (.A(_06176_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_2 _21333_ (.A0(\fetch.bht.bhtTable_tag[1][18] ),
    .A1(_10772_),
    .S(_06168_),
    .X(_06177_));
 sky130_fd_sc_hd__buf_1 _21334_ (.A(_06177_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_2 _21335_ (.A0(\fetch.bht.bhtTable_tag[1][19] ),
    .A1(_10773_),
    .S(_06168_),
    .X(_06178_));
 sky130_fd_sc_hd__buf_1 _21336_ (.A(_06178_),
    .X(_01003_));
 sky130_fd_sc_hd__buf_1 _21337_ (.A(_06155_),
    .X(_06179_));
 sky130_fd_sc_hd__mux2_2 _21338_ (.A0(\fetch.bht.bhtTable_tag[1][20] ),
    .A1(_10760_),
    .S(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__buf_1 _21339_ (.A(_06180_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_2 _21340_ (.A0(\fetch.bht.bhtTable_tag[1][21] ),
    .A1(_10759_),
    .S(_06179_),
    .X(_06181_));
 sky130_fd_sc_hd__buf_1 _21341_ (.A(_06181_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_2 _21342_ (.A0(\fetch.bht.bhtTable_tag[1][22] ),
    .A1(_10771_),
    .S(_06179_),
    .X(_06182_));
 sky130_fd_sc_hd__buf_1 _21343_ (.A(_06182_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_2 _21344_ (.A0(\fetch.bht.bhtTable_tag[1][23] ),
    .A1(\csr.io_mem_pc[29] ),
    .S(_06179_),
    .X(_06183_));
 sky130_fd_sc_hd__buf_1 _21345_ (.A(_06183_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_2 _21346_ (.A0(\fetch.bht.bhtTable_tag[1][24] ),
    .A1(_10777_),
    .S(_06179_),
    .X(_06184_));
 sky130_fd_sc_hd__buf_1 _21347_ (.A(_06184_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_2 _21348_ (.A0(\fetch.bht.bhtTable_tag[1][25] ),
    .A1(\csr.io_mem_pc[31] ),
    .S(_06179_),
    .X(_06185_));
 sky130_fd_sc_hd__buf_1 _21349_ (.A(_06185_),
    .X(_01009_));
 sky130_fd_sc_hd__nand4_2 _21350_ (.A(_10556_),
    .B(_10557_),
    .C(_09885_),
    .D(_09916_),
    .Y(_06186_));
 sky130_fd_sc_hd__buf_1 _21351_ (.A(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__buf_1 _21352_ (.A(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__mux2_2 _21353_ (.A0(_06101_),
    .A1(\fetch.bht.bhtTable_tag[7][0] ),
    .S(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__buf_1 _21354_ (.A(_06189_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_2 _21355_ (.A0(_06103_),
    .A1(\fetch.bht.bhtTable_tag[7][1] ),
    .S(_06188_),
    .X(_06190_));
 sky130_fd_sc_hd__buf_1 _21356_ (.A(_06190_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_2 _21357_ (.A0(_06105_),
    .A1(\fetch.bht.bhtTable_tag[7][2] ),
    .S(_06188_),
    .X(_06191_));
 sky130_fd_sc_hd__buf_1 _21358_ (.A(_06191_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_2 _21359_ (.A0(_06107_),
    .A1(\fetch.bht.bhtTable_tag[7][3] ),
    .S(_06188_),
    .X(_06192_));
 sky130_fd_sc_hd__buf_1 _21360_ (.A(_06192_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_2 _21361_ (.A0(_06109_),
    .A1(\fetch.bht.bhtTable_tag[7][4] ),
    .S(_06188_),
    .X(_06193_));
 sky130_fd_sc_hd__buf_1 _21362_ (.A(_06193_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_2 _21363_ (.A0(_06111_),
    .A1(\fetch.bht.bhtTable_tag[7][5] ),
    .S(_06188_),
    .X(_06194_));
 sky130_fd_sc_hd__buf_1 _21364_ (.A(_06194_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_2 _21365_ (.A0(_06113_),
    .A1(\fetch.bht.bhtTable_tag[7][6] ),
    .S(_06188_),
    .X(_06195_));
 sky130_fd_sc_hd__buf_1 _21366_ (.A(_06195_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_2 _21367_ (.A0(_06115_),
    .A1(\fetch.bht.bhtTable_tag[7][7] ),
    .S(_06188_),
    .X(_06196_));
 sky130_fd_sc_hd__buf_1 _21368_ (.A(_06196_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_2 _21369_ (.A0(_06117_),
    .A1(\fetch.bht.bhtTable_tag[7][8] ),
    .S(_06188_),
    .X(_06197_));
 sky130_fd_sc_hd__buf_1 _21370_ (.A(_06197_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_2 _21371_ (.A0(_06119_),
    .A1(\fetch.bht.bhtTable_tag[7][9] ),
    .S(_06188_),
    .X(_06198_));
 sky130_fd_sc_hd__buf_1 _21372_ (.A(_06198_),
    .X(_01019_));
 sky130_fd_sc_hd__buf_1 _21373_ (.A(_06187_),
    .X(_06199_));
 sky130_fd_sc_hd__mux2_2 _21374_ (.A0(_06122_),
    .A1(\fetch.bht.bhtTable_tag[7][10] ),
    .S(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__buf_1 _21375_ (.A(_06200_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_2 _21376_ (.A0(_06124_),
    .A1(\fetch.bht.bhtTable_tag[7][11] ),
    .S(_06199_),
    .X(_06201_));
 sky130_fd_sc_hd__buf_1 _21377_ (.A(_06201_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_2 _21378_ (.A0(_06126_),
    .A1(\fetch.bht.bhtTable_tag[7][12] ),
    .S(_06199_),
    .X(_06202_));
 sky130_fd_sc_hd__buf_1 _21379_ (.A(_06202_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_2 _21380_ (.A0(_06128_),
    .A1(\fetch.bht.bhtTable_tag[7][13] ),
    .S(_06199_),
    .X(_06203_));
 sky130_fd_sc_hd__buf_1 _21381_ (.A(_06203_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_2 _21382_ (.A0(_06130_),
    .A1(\fetch.bht.bhtTable_tag[7][14] ),
    .S(_06199_),
    .X(_06204_));
 sky130_fd_sc_hd__buf_1 _21383_ (.A(_06204_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_2 _21384_ (.A0(_06132_),
    .A1(\fetch.bht.bhtTable_tag[7][15] ),
    .S(_06199_),
    .X(_06205_));
 sky130_fd_sc_hd__buf_1 _21385_ (.A(_06205_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_2 _21386_ (.A0(_06134_),
    .A1(\fetch.bht.bhtTable_tag[7][16] ),
    .S(_06199_),
    .X(_06206_));
 sky130_fd_sc_hd__buf_1 _21387_ (.A(_06206_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_2 _21388_ (.A0(_06136_),
    .A1(\fetch.bht.bhtTable_tag[7][17] ),
    .S(_06199_),
    .X(_06207_));
 sky130_fd_sc_hd__buf_1 _21389_ (.A(_06207_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_2 _21390_ (.A0(_06138_),
    .A1(\fetch.bht.bhtTable_tag[7][18] ),
    .S(_06199_),
    .X(_06208_));
 sky130_fd_sc_hd__buf_1 _21391_ (.A(_06208_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_2 _21392_ (.A0(_06140_),
    .A1(\fetch.bht.bhtTable_tag[7][19] ),
    .S(_06199_),
    .X(_06209_));
 sky130_fd_sc_hd__buf_1 _21393_ (.A(_06209_),
    .X(_01029_));
 sky130_fd_sc_hd__buf_1 _21394_ (.A(_06186_),
    .X(_06210_));
 sky130_fd_sc_hd__mux2_2 _21395_ (.A0(_06143_),
    .A1(\fetch.bht.bhtTable_tag[7][20] ),
    .S(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__buf_1 _21396_ (.A(_06211_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_2 _21397_ (.A0(_06145_),
    .A1(\fetch.bht.bhtTable_tag[7][21] ),
    .S(_06210_),
    .X(_06212_));
 sky130_fd_sc_hd__buf_1 _21398_ (.A(_06212_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_2 _21399_ (.A0(_06147_),
    .A1(\fetch.bht.bhtTable_tag[7][22] ),
    .S(_06210_),
    .X(_06213_));
 sky130_fd_sc_hd__buf_1 _21400_ (.A(_06213_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_2 _21401_ (.A0(_06149_),
    .A1(\fetch.bht.bhtTable_tag[7][23] ),
    .S(_06210_),
    .X(_06214_));
 sky130_fd_sc_hd__buf_1 _21402_ (.A(_06214_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_2 _21403_ (.A0(_06151_),
    .A1(\fetch.bht.bhtTable_tag[7][24] ),
    .S(_06210_),
    .X(_06215_));
 sky130_fd_sc_hd__buf_1 _21404_ (.A(_06215_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_2 _21405_ (.A0(_06153_),
    .A1(\fetch.bht.bhtTable_tag[7][25] ),
    .S(_06210_),
    .X(_06216_));
 sky130_fd_sc_hd__buf_1 _21406_ (.A(_06216_),
    .X(_01035_));
 sky130_fd_sc_hd__or4bb_2 _21407_ (.A(_09900_),
    .B(_10556_),
    .C_N(_10557_),
    .D_N(_09916_),
    .X(_06217_));
 sky130_fd_sc_hd__buf_1 _21408_ (.A(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__buf_1 _21409_ (.A(_06218_),
    .X(_06219_));
 sky130_fd_sc_hd__mux2_2 _21410_ (.A0(_06101_),
    .A1(\fetch.bht.bhtTable_tag[6][0] ),
    .S(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__buf_1 _21411_ (.A(_06220_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_2 _21412_ (.A0(_06103_),
    .A1(\fetch.bht.bhtTable_tag[6][1] ),
    .S(_06219_),
    .X(_06221_));
 sky130_fd_sc_hd__buf_1 _21413_ (.A(_06221_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_2 _21414_ (.A0(_06105_),
    .A1(\fetch.bht.bhtTable_tag[6][2] ),
    .S(_06219_),
    .X(_06222_));
 sky130_fd_sc_hd__buf_1 _21415_ (.A(_06222_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_2 _21416_ (.A0(_06107_),
    .A1(\fetch.bht.bhtTable_tag[6][3] ),
    .S(_06219_),
    .X(_06223_));
 sky130_fd_sc_hd__buf_1 _21417_ (.A(_06223_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_2 _21418_ (.A0(_06109_),
    .A1(\fetch.bht.bhtTable_tag[6][4] ),
    .S(_06219_),
    .X(_06224_));
 sky130_fd_sc_hd__buf_1 _21419_ (.A(_06224_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_2 _21420_ (.A0(_06111_),
    .A1(\fetch.bht.bhtTable_tag[6][5] ),
    .S(_06219_),
    .X(_06225_));
 sky130_fd_sc_hd__buf_1 _21421_ (.A(_06225_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_2 _21422_ (.A0(_06113_),
    .A1(\fetch.bht.bhtTable_tag[6][6] ),
    .S(_06219_),
    .X(_06226_));
 sky130_fd_sc_hd__buf_1 _21423_ (.A(_06226_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_2 _21424_ (.A0(_06115_),
    .A1(\fetch.bht.bhtTable_tag[6][7] ),
    .S(_06219_),
    .X(_06227_));
 sky130_fd_sc_hd__buf_1 _21425_ (.A(_06227_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_2 _21426_ (.A0(_06117_),
    .A1(\fetch.bht.bhtTable_tag[6][8] ),
    .S(_06219_),
    .X(_06228_));
 sky130_fd_sc_hd__buf_1 _21427_ (.A(_06228_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_2 _21428_ (.A0(_06119_),
    .A1(\fetch.bht.bhtTable_tag[6][9] ),
    .S(_06219_),
    .X(_06229_));
 sky130_fd_sc_hd__buf_1 _21429_ (.A(_06229_),
    .X(_01045_));
 sky130_fd_sc_hd__buf_1 _21430_ (.A(_06218_),
    .X(_06230_));
 sky130_fd_sc_hd__mux2_2 _21431_ (.A0(_06122_),
    .A1(\fetch.bht.bhtTable_tag[6][10] ),
    .S(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__buf_1 _21432_ (.A(_06231_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_2 _21433_ (.A0(_06124_),
    .A1(\fetch.bht.bhtTable_tag[6][11] ),
    .S(_06230_),
    .X(_06232_));
 sky130_fd_sc_hd__buf_1 _21434_ (.A(_06232_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_2 _21435_ (.A0(_06126_),
    .A1(\fetch.bht.bhtTable_tag[6][12] ),
    .S(_06230_),
    .X(_06233_));
 sky130_fd_sc_hd__buf_1 _21436_ (.A(_06233_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_2 _21437_ (.A0(_06128_),
    .A1(\fetch.bht.bhtTable_tag[6][13] ),
    .S(_06230_),
    .X(_06234_));
 sky130_fd_sc_hd__buf_1 _21438_ (.A(_06234_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_2 _21439_ (.A0(_06130_),
    .A1(\fetch.bht.bhtTable_tag[6][14] ),
    .S(_06230_),
    .X(_06235_));
 sky130_fd_sc_hd__buf_1 _21440_ (.A(_06235_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_2 _21441_ (.A0(_06132_),
    .A1(\fetch.bht.bhtTable_tag[6][15] ),
    .S(_06230_),
    .X(_06236_));
 sky130_fd_sc_hd__buf_1 _21442_ (.A(_06236_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_2 _21443_ (.A0(_06134_),
    .A1(\fetch.bht.bhtTable_tag[6][16] ),
    .S(_06230_),
    .X(_06237_));
 sky130_fd_sc_hd__buf_1 _21444_ (.A(_06237_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_2 _21445_ (.A0(_06136_),
    .A1(\fetch.bht.bhtTable_tag[6][17] ),
    .S(_06230_),
    .X(_06238_));
 sky130_fd_sc_hd__buf_1 _21446_ (.A(_06238_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_2 _21447_ (.A0(_06138_),
    .A1(\fetch.bht.bhtTable_tag[6][18] ),
    .S(_06230_),
    .X(_06239_));
 sky130_fd_sc_hd__buf_1 _21448_ (.A(_06239_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_2 _21449_ (.A0(_06140_),
    .A1(\fetch.bht.bhtTable_tag[6][19] ),
    .S(_06230_),
    .X(_06240_));
 sky130_fd_sc_hd__buf_1 _21450_ (.A(_06240_),
    .X(_01055_));
 sky130_fd_sc_hd__buf_1 _21451_ (.A(_06217_),
    .X(_06241_));
 sky130_fd_sc_hd__mux2_2 _21452_ (.A0(_06143_),
    .A1(\fetch.bht.bhtTable_tag[6][20] ),
    .S(_06241_),
    .X(_06242_));
 sky130_fd_sc_hd__buf_1 _21453_ (.A(_06242_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_2 _21454_ (.A0(_06145_),
    .A1(\fetch.bht.bhtTable_tag[6][21] ),
    .S(_06241_),
    .X(_06243_));
 sky130_fd_sc_hd__buf_1 _21455_ (.A(_06243_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_2 _21456_ (.A0(_06147_),
    .A1(\fetch.bht.bhtTable_tag[6][22] ),
    .S(_06241_),
    .X(_06244_));
 sky130_fd_sc_hd__buf_1 _21457_ (.A(_06244_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_2 _21458_ (.A0(_06149_),
    .A1(\fetch.bht.bhtTable_tag[6][23] ),
    .S(_06241_),
    .X(_06245_));
 sky130_fd_sc_hd__buf_1 _21459_ (.A(_06245_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_2 _21460_ (.A0(_06151_),
    .A1(\fetch.bht.bhtTable_tag[6][24] ),
    .S(_06241_),
    .X(_06246_));
 sky130_fd_sc_hd__buf_1 _21461_ (.A(_06246_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_2 _21462_ (.A0(_06153_),
    .A1(\fetch.bht.bhtTable_tag[6][25] ),
    .S(_06241_),
    .X(_06247_));
 sky130_fd_sc_hd__buf_1 _21463_ (.A(_06247_),
    .X(_01061_));
 sky130_fd_sc_hd__o31a_2 _21464_ (.A1(io_fetch_data[0]),
    .A2(_10673_),
    .A3(_10911_),
    .B1(_09957_),
    .X(_01062_));
 sky130_fd_sc_hd__o31a_2 _21465_ (.A1(io_fetch_data[1]),
    .A2(_10673_),
    .A3(_10911_),
    .B1(_09957_),
    .X(_01063_));
 sky130_fd_sc_hd__buf_1 _21466_ (.A(_05246_),
    .X(_06248_));
 sky130_fd_sc_hd__or4_2 _21467_ (.A(_10964_),
    .B(_06248_),
    .C(_10915_),
    .D(_10908_),
    .X(_06249_));
 sky130_fd_sc_hd__o211a_2 _21468_ (.A1(io_fetch_data[4]),
    .A2(_10972_),
    .B1(_06249_),
    .C1(_10546_),
    .X(_01064_));
 sky130_fd_sc_hd__or4bb_2 _21469_ (.A(_10557_),
    .B(_09900_),
    .C_N(_09916_),
    .D_N(_10556_),
    .X(_06250_));
 sky130_fd_sc_hd__buf_1 _21470_ (.A(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__buf_1 _21471_ (.A(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__mux2_2 _21472_ (.A0(_06101_),
    .A1(\fetch.bht.bhtTable_tag[5][0] ),
    .S(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__buf_1 _21473_ (.A(_06253_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_2 _21474_ (.A0(_06103_),
    .A1(\fetch.bht.bhtTable_tag[5][1] ),
    .S(_06252_),
    .X(_06254_));
 sky130_fd_sc_hd__buf_1 _21475_ (.A(_06254_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_2 _21476_ (.A0(_06105_),
    .A1(\fetch.bht.bhtTable_tag[5][2] ),
    .S(_06252_),
    .X(_06255_));
 sky130_fd_sc_hd__buf_1 _21477_ (.A(_06255_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_2 _21478_ (.A0(_06107_),
    .A1(\fetch.bht.bhtTable_tag[5][3] ),
    .S(_06252_),
    .X(_06256_));
 sky130_fd_sc_hd__buf_1 _21479_ (.A(_06256_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_2 _21480_ (.A0(_06109_),
    .A1(\fetch.bht.bhtTable_tag[5][4] ),
    .S(_06252_),
    .X(_06257_));
 sky130_fd_sc_hd__buf_1 _21481_ (.A(_06257_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_2 _21482_ (.A0(_06111_),
    .A1(\fetch.bht.bhtTable_tag[5][5] ),
    .S(_06252_),
    .X(_06258_));
 sky130_fd_sc_hd__buf_1 _21483_ (.A(_06258_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_2 _21484_ (.A0(_06113_),
    .A1(\fetch.bht.bhtTable_tag[5][6] ),
    .S(_06252_),
    .X(_06259_));
 sky130_fd_sc_hd__buf_1 _21485_ (.A(_06259_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_2 _21486_ (.A0(_06115_),
    .A1(\fetch.bht.bhtTable_tag[5][7] ),
    .S(_06252_),
    .X(_06260_));
 sky130_fd_sc_hd__buf_1 _21487_ (.A(_06260_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_2 _21488_ (.A0(_06117_),
    .A1(\fetch.bht.bhtTable_tag[5][8] ),
    .S(_06252_),
    .X(_06261_));
 sky130_fd_sc_hd__buf_1 _21489_ (.A(_06261_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_2 _21490_ (.A0(_06119_),
    .A1(\fetch.bht.bhtTable_tag[5][9] ),
    .S(_06252_),
    .X(_06262_));
 sky130_fd_sc_hd__buf_1 _21491_ (.A(_06262_),
    .X(_01074_));
 sky130_fd_sc_hd__buf_1 _21492_ (.A(_06251_),
    .X(_06263_));
 sky130_fd_sc_hd__mux2_2 _21493_ (.A0(_06122_),
    .A1(\fetch.bht.bhtTable_tag[5][10] ),
    .S(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__buf_1 _21494_ (.A(_06264_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_2 _21495_ (.A0(_06124_),
    .A1(\fetch.bht.bhtTable_tag[5][11] ),
    .S(_06263_),
    .X(_06265_));
 sky130_fd_sc_hd__buf_1 _21496_ (.A(_06265_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_2 _21497_ (.A0(_06126_),
    .A1(\fetch.bht.bhtTable_tag[5][12] ),
    .S(_06263_),
    .X(_06266_));
 sky130_fd_sc_hd__buf_1 _21498_ (.A(_06266_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_2 _21499_ (.A0(_06128_),
    .A1(\fetch.bht.bhtTable_tag[5][13] ),
    .S(_06263_),
    .X(_06267_));
 sky130_fd_sc_hd__buf_1 _21500_ (.A(_06267_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_2 _21501_ (.A0(_06130_),
    .A1(\fetch.bht.bhtTable_tag[5][14] ),
    .S(_06263_),
    .X(_06268_));
 sky130_fd_sc_hd__buf_1 _21502_ (.A(_06268_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_2 _21503_ (.A0(_06132_),
    .A1(\fetch.bht.bhtTable_tag[5][15] ),
    .S(_06263_),
    .X(_06269_));
 sky130_fd_sc_hd__buf_1 _21504_ (.A(_06269_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_2 _21505_ (.A0(_06134_),
    .A1(\fetch.bht.bhtTable_tag[5][16] ),
    .S(_06263_),
    .X(_06270_));
 sky130_fd_sc_hd__buf_1 _21506_ (.A(_06270_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_2 _21507_ (.A0(_06136_),
    .A1(\fetch.bht.bhtTable_tag[5][17] ),
    .S(_06263_),
    .X(_06271_));
 sky130_fd_sc_hd__buf_1 _21508_ (.A(_06271_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_2 _21509_ (.A0(_06138_),
    .A1(\fetch.bht.bhtTable_tag[5][18] ),
    .S(_06263_),
    .X(_06272_));
 sky130_fd_sc_hd__buf_1 _21510_ (.A(_06272_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_2 _21511_ (.A0(_06140_),
    .A1(\fetch.bht.bhtTable_tag[5][19] ),
    .S(_06263_),
    .X(_06273_));
 sky130_fd_sc_hd__buf_1 _21512_ (.A(_06273_),
    .X(_01084_));
 sky130_fd_sc_hd__buf_1 _21513_ (.A(_06250_),
    .X(_06274_));
 sky130_fd_sc_hd__mux2_2 _21514_ (.A0(_06143_),
    .A1(\fetch.bht.bhtTable_tag[5][20] ),
    .S(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__buf_1 _21515_ (.A(_06275_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_2 _21516_ (.A0(_06145_),
    .A1(\fetch.bht.bhtTable_tag[5][21] ),
    .S(_06274_),
    .X(_06276_));
 sky130_fd_sc_hd__buf_1 _21517_ (.A(_06276_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_2 _21518_ (.A0(_06147_),
    .A1(\fetch.bht.bhtTable_tag[5][22] ),
    .S(_06274_),
    .X(_06277_));
 sky130_fd_sc_hd__buf_1 _21519_ (.A(_06277_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_2 _21520_ (.A0(_06149_),
    .A1(\fetch.bht.bhtTable_tag[5][23] ),
    .S(_06274_),
    .X(_06278_));
 sky130_fd_sc_hd__buf_1 _21521_ (.A(_06278_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_2 _21522_ (.A0(_06151_),
    .A1(\fetch.bht.bhtTable_tag[5][24] ),
    .S(_06274_),
    .X(_06279_));
 sky130_fd_sc_hd__buf_1 _21523_ (.A(_06279_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_2 _21524_ (.A0(_06153_),
    .A1(\fetch.bht.bhtTable_tag[5][25] ),
    .S(_06274_),
    .X(_06280_));
 sky130_fd_sc_hd__buf_1 _21525_ (.A(_06280_),
    .X(_01090_));
 sky130_fd_sc_hd__nand2_2 _21526_ (.A(_09879_),
    .B(_09882_),
    .Y(_06281_));
 sky130_fd_sc_hd__or4b_2 _21527_ (.A(_10557_),
    .B(_09900_),
    .C(_06281_),
    .D_N(_10556_),
    .X(_06282_));
 sky130_fd_sc_hd__buf_1 _21528_ (.A(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__buf_1 _21529_ (.A(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__mux2_2 _21530_ (.A0(_06101_),
    .A1(\fetch.bht.bhtTable_tag[13][0] ),
    .S(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__buf_1 _21531_ (.A(_06285_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_2 _21532_ (.A0(_06103_),
    .A1(\fetch.bht.bhtTable_tag[13][1] ),
    .S(_06284_),
    .X(_06286_));
 sky130_fd_sc_hd__buf_1 _21533_ (.A(_06286_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_2 _21534_ (.A0(_06105_),
    .A1(\fetch.bht.bhtTable_tag[13][2] ),
    .S(_06284_),
    .X(_06287_));
 sky130_fd_sc_hd__buf_1 _21535_ (.A(_06287_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_2 _21536_ (.A0(_06107_),
    .A1(\fetch.bht.bhtTable_tag[13][3] ),
    .S(_06284_),
    .X(_06288_));
 sky130_fd_sc_hd__buf_1 _21537_ (.A(_06288_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_2 _21538_ (.A0(_06109_),
    .A1(\fetch.bht.bhtTable_tag[13][4] ),
    .S(_06284_),
    .X(_06289_));
 sky130_fd_sc_hd__buf_1 _21539_ (.A(_06289_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_2 _21540_ (.A0(_06111_),
    .A1(\fetch.bht.bhtTable_tag[13][5] ),
    .S(_06284_),
    .X(_06290_));
 sky130_fd_sc_hd__buf_1 _21541_ (.A(_06290_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_2 _21542_ (.A0(_06113_),
    .A1(\fetch.bht.bhtTable_tag[13][6] ),
    .S(_06284_),
    .X(_06291_));
 sky130_fd_sc_hd__buf_1 _21543_ (.A(_06291_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_2 _21544_ (.A0(_06115_),
    .A1(\fetch.bht.bhtTable_tag[13][7] ),
    .S(_06284_),
    .X(_06292_));
 sky130_fd_sc_hd__buf_1 _21545_ (.A(_06292_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_2 _21546_ (.A0(_06117_),
    .A1(\fetch.bht.bhtTable_tag[13][8] ),
    .S(_06284_),
    .X(_06293_));
 sky130_fd_sc_hd__buf_1 _21547_ (.A(_06293_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_2 _21548_ (.A0(_06119_),
    .A1(\fetch.bht.bhtTable_tag[13][9] ),
    .S(_06284_),
    .X(_06294_));
 sky130_fd_sc_hd__buf_1 _21549_ (.A(_06294_),
    .X(_01100_));
 sky130_fd_sc_hd__buf_1 _21550_ (.A(_06283_),
    .X(_06295_));
 sky130_fd_sc_hd__mux2_2 _21551_ (.A0(_06122_),
    .A1(\fetch.bht.bhtTable_tag[13][10] ),
    .S(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__buf_1 _21552_ (.A(_06296_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_2 _21553_ (.A0(_06124_),
    .A1(\fetch.bht.bhtTable_tag[13][11] ),
    .S(_06295_),
    .X(_06297_));
 sky130_fd_sc_hd__buf_1 _21554_ (.A(_06297_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_2 _21555_ (.A0(_06126_),
    .A1(\fetch.bht.bhtTable_tag[13][12] ),
    .S(_06295_),
    .X(_06298_));
 sky130_fd_sc_hd__buf_1 _21556_ (.A(_06298_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_2 _21557_ (.A0(_06128_),
    .A1(\fetch.bht.bhtTable_tag[13][13] ),
    .S(_06295_),
    .X(_06299_));
 sky130_fd_sc_hd__buf_1 _21558_ (.A(_06299_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_2 _21559_ (.A0(_06130_),
    .A1(\fetch.bht.bhtTable_tag[13][14] ),
    .S(_06295_),
    .X(_06300_));
 sky130_fd_sc_hd__buf_1 _21560_ (.A(_06300_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_2 _21561_ (.A0(_06132_),
    .A1(\fetch.bht.bhtTable_tag[13][15] ),
    .S(_06295_),
    .X(_06301_));
 sky130_fd_sc_hd__buf_1 _21562_ (.A(_06301_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_2 _21563_ (.A0(_06134_),
    .A1(\fetch.bht.bhtTable_tag[13][16] ),
    .S(_06295_),
    .X(_06302_));
 sky130_fd_sc_hd__buf_1 _21564_ (.A(_06302_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_2 _21565_ (.A0(_06136_),
    .A1(\fetch.bht.bhtTable_tag[13][17] ),
    .S(_06295_),
    .X(_06303_));
 sky130_fd_sc_hd__buf_1 _21566_ (.A(_06303_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_2 _21567_ (.A0(_06138_),
    .A1(\fetch.bht.bhtTable_tag[13][18] ),
    .S(_06295_),
    .X(_06304_));
 sky130_fd_sc_hd__buf_1 _21568_ (.A(_06304_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_2 _21569_ (.A0(_06140_),
    .A1(\fetch.bht.bhtTable_tag[13][19] ),
    .S(_06295_),
    .X(_06305_));
 sky130_fd_sc_hd__buf_1 _21570_ (.A(_06305_),
    .X(_01110_));
 sky130_fd_sc_hd__buf_1 _21571_ (.A(_06282_),
    .X(_06306_));
 sky130_fd_sc_hd__mux2_2 _21572_ (.A0(_06143_),
    .A1(\fetch.bht.bhtTable_tag[13][20] ),
    .S(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__buf_1 _21573_ (.A(_06307_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_2 _21574_ (.A0(_06145_),
    .A1(\fetch.bht.bhtTable_tag[13][21] ),
    .S(_06306_),
    .X(_06308_));
 sky130_fd_sc_hd__buf_1 _21575_ (.A(_06308_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_2 _21576_ (.A0(_06147_),
    .A1(\fetch.bht.bhtTable_tag[13][22] ),
    .S(_06306_),
    .X(_06309_));
 sky130_fd_sc_hd__buf_1 _21577_ (.A(_06309_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_2 _21578_ (.A0(_06149_),
    .A1(\fetch.bht.bhtTable_tag[13][23] ),
    .S(_06306_),
    .X(_06310_));
 sky130_fd_sc_hd__buf_1 _21579_ (.A(_06310_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_2 _21580_ (.A0(_06151_),
    .A1(\fetch.bht.bhtTable_tag[13][24] ),
    .S(_06306_),
    .X(_06311_));
 sky130_fd_sc_hd__buf_1 _21581_ (.A(_06311_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_2 _21582_ (.A0(_06153_),
    .A1(\fetch.bht.bhtTable_tag[13][25] ),
    .S(_06306_),
    .X(_06312_));
 sky130_fd_sc_hd__buf_1 _21583_ (.A(_06312_),
    .X(_01116_));
 sky130_fd_sc_hd__nor4_2 _21584_ (.A(\csr.io_csr_write_address[5] ),
    .B(\csr.io_csr_write_address[4] ),
    .C(\csr.io_csr_write_address[7] ),
    .D(\csr.io_csr_write_address[6] ),
    .Y(_06313_));
 sky130_fd_sc_hd__and3b_2 _21585_ (.A_N(\csr.io_csr_write_address[10] ),
    .B(\csr.io_csr_write_address[8] ),
    .C(\csr.io_csr_write_address[9] ),
    .X(_06314_));
 sky130_fd_sc_hd__or3b_2 _21586_ (.A(\csr.io_csr_write_address[3] ),
    .B(\csr.io_csr_write_address[2] ),
    .C_N(\csr.io_csr_write_enable ),
    .X(_06315_));
 sky130_fd_sc_hd__nor3b_2 _21587_ (.A(\csr.io_csr_write_address[0] ),
    .B(_06315_),
    .C_N(\csr.io_csr_write_address[1] ),
    .Y(_06316_));
 sky130_fd_sc_hd__nand4_2 _21588_ (.A(\csr.io_csr_write_address[11] ),
    .B(_06313_),
    .C(_06314_),
    .D(_06316_),
    .Y(_06317_));
 sky130_fd_sc_hd__buf_1 _21589_ (.A(_10576_),
    .X(_06318_));
 sky130_fd_sc_hd__and4_2 _21590_ (.A(\csr.io_csr_write_address[11] ),
    .B(_06313_),
    .C(_06314_),
    .D(_06316_),
    .X(_06319_));
 sky130_fd_sc_hd__buf_1 _21591_ (.A(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__buf_1 _21592_ (.A(_06320_),
    .X(_06321_));
 sky130_fd_sc_hd__and2_2 _21593_ (.A(_06317_),
    .B(\csr.io_inst_retired ),
    .X(_06322_));
 sky130_fd_sc_hd__buf_1 _21594_ (.A(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__a211oi_2 _21595_ (.A1(\csr._mcycle_T_2[0] ),
    .A2(_06321_),
    .B1(_06323_),
    .C1(\csr.minstret[0] ),
    .Y(_06324_));
 sky130_fd_sc_hd__a311oi_2 _21596_ (.A1(\csr.minstret[0] ),
    .A2(_06317_),
    .A3(\csr.io_inst_retired ),
    .B1(_06318_),
    .C1(_06324_),
    .Y(_01117_));
 sky130_fd_sc_hd__buf_1 _21597_ (.A(_06320_),
    .X(_06325_));
 sky130_fd_sc_hd__a221oi_2 _21598_ (.A1(\csr._mcycle_T_2[1] ),
    .A2(_06325_),
    .B1(_06323_),
    .B2(\csr.minstret[0] ),
    .C1(\csr.minstret[1] ),
    .Y(_06326_));
 sky130_fd_sc_hd__buf_1 _21599_ (.A(_10576_),
    .X(_06327_));
 sky130_fd_sc_hd__a311oi_2 _21600_ (.A1(\csr.minstret[0] ),
    .A2(\csr.minstret[1] ),
    .A3(_06323_),
    .B1(_06326_),
    .C1(_06327_),
    .Y(_01118_));
 sky130_fd_sc_hd__and3_2 _21601_ (.A(\csr.minstret[0] ),
    .B(\csr.minstret[1] ),
    .C(_06323_),
    .X(_06328_));
 sky130_fd_sc_hd__buf_1 _21602_ (.A(_06320_),
    .X(_06329_));
 sky130_fd_sc_hd__a211oi_2 _21603_ (.A1(\csr._mcycle_T_2[2] ),
    .A2(_06329_),
    .B1(_06328_),
    .C1(\csr.minstret[2] ),
    .Y(_06330_));
 sky130_fd_sc_hd__buf_1 _21604_ (.A(_03579_),
    .X(_06331_));
 sky130_fd_sc_hd__a211oi_2 _21605_ (.A1(\csr.minstret[2] ),
    .A2(_06328_),
    .B1(_06330_),
    .C1(_06331_),
    .Y(_01119_));
 sky130_fd_sc_hd__and4_2 _21606_ (.A(\csr.minstret[0] ),
    .B(\csr.minstret[1] ),
    .C(\csr.minstret[2] ),
    .D(\csr.minstret[3] ),
    .X(_06332_));
 sky130_fd_sc_hd__buf_1 _21607_ (.A(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__a221oi_2 _21608_ (.A1(\csr._mcycle_T_2[3] ),
    .A2(_06325_),
    .B1(_06328_),
    .B2(\csr.minstret[2] ),
    .C1(\csr.minstret[3] ),
    .Y(_06334_));
 sky130_fd_sc_hd__a211oi_2 _21609_ (.A1(_06323_),
    .A2(_06333_),
    .B1(_06334_),
    .C1(_06331_),
    .Y(_01120_));
 sky130_fd_sc_hd__a221oi_2 _21610_ (.A1(\csr._mcycle_T_2[4] ),
    .A2(_06325_),
    .B1(_06323_),
    .B2(_06333_),
    .C1(_05613_),
    .Y(_06335_));
 sky130_fd_sc_hd__buf_1 _21611_ (.A(_10576_),
    .X(_06336_));
 sky130_fd_sc_hd__a311oi_2 _21612_ (.A1(_05613_),
    .A2(_06323_),
    .A3(_06333_),
    .B1(_06335_),
    .C1(_06336_),
    .Y(_01121_));
 sky130_fd_sc_hd__and3_2 _21613_ (.A(_06317_),
    .B(_06333_),
    .C(\csr.io_inst_retired ),
    .X(_06337_));
 sky130_fd_sc_hd__buf_1 _21614_ (.A(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__a221oi_2 _21615_ (.A1(\csr._mcycle_T_2[5] ),
    .A2(_06325_),
    .B1(_06338_),
    .B2(_05613_),
    .C1(\csr.minstret[5] ),
    .Y(_06339_));
 sky130_fd_sc_hd__a311oi_2 _21616_ (.A1(_05613_),
    .A2(\csr.minstret[5] ),
    .A3(_06338_),
    .B1(_06339_),
    .C1(_06336_),
    .Y(_01122_));
 sky130_fd_sc_hd__and3_2 _21617_ (.A(_05613_),
    .B(\csr.minstret[5] ),
    .C(_06338_),
    .X(_06340_));
 sky130_fd_sc_hd__a211oi_2 _21618_ (.A1(\csr._mcycle_T_2[6] ),
    .A2(_06329_),
    .B1(_06340_),
    .C1(\csr.minstret[6] ),
    .Y(_06341_));
 sky130_fd_sc_hd__a211oi_2 _21619_ (.A1(\csr.minstret[6] ),
    .A2(_06340_),
    .B1(_06341_),
    .C1(_06331_),
    .Y(_01123_));
 sky130_fd_sc_hd__and4_2 _21620_ (.A(_05613_),
    .B(\csr.minstret[5] ),
    .C(\csr.io_inst_retired ),
    .D(_06333_),
    .X(_06342_));
 sky130_fd_sc_hd__a21oi_2 _21621_ (.A1(\csr.minstret[6] ),
    .A2(_06342_),
    .B1(\csr.minstret[7] ),
    .Y(_06343_));
 sky130_fd_sc_hd__and3_2 _21622_ (.A(\csr.minstret[6] ),
    .B(\csr.minstret[7] ),
    .C(_06342_),
    .X(_06344_));
 sky130_fd_sc_hd__o21ai_2 _21623_ (.A1(_06343_),
    .A2(_06344_),
    .B1(_06317_),
    .Y(_06345_));
 sky130_fd_sc_hd__o311a_2 _21624_ (.A1(\csr._mcycle_T_2[7] ),
    .A2(_06317_),
    .A3(\csr.minstret[7] ),
    .B1(_05856_),
    .C1(_06345_),
    .X(_01124_));
 sky130_fd_sc_hd__and4_2 _21625_ (.A(_06317_),
    .B(_06342_),
    .C(\csr.minstret[6] ),
    .D(\csr.minstret[7] ),
    .X(_06346_));
 sky130_fd_sc_hd__a211oi_2 _21626_ (.A1(\csr._mcycle_T_2[8] ),
    .A2(_06329_),
    .B1(_06346_),
    .C1(\csr.minstret[8] ),
    .Y(_06347_));
 sky130_fd_sc_hd__a211oi_2 _21627_ (.A1(\csr.minstret[8] ),
    .A2(_06346_),
    .B1(_06347_),
    .C1(_06331_),
    .Y(_01125_));
 sky130_fd_sc_hd__a221oi_2 _21628_ (.A1(\csr._mcycle_T_2[9] ),
    .A2(_06321_),
    .B1(_06346_),
    .B2(\csr.minstret[8] ),
    .C1(\csr.minstret[9] ),
    .Y(_06348_));
 sky130_fd_sc_hd__and4_2 _21629_ (.A(\csr.minstret[6] ),
    .B(\csr.minstret[7] ),
    .C(\csr.minstret[8] ),
    .D(\csr.minstret[9] ),
    .X(_06349_));
 sky130_fd_sc_hd__and4_2 _21630_ (.A(_05613_),
    .B(\csr.minstret[5] ),
    .C(_06338_),
    .D(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__nor3_2 _21631_ (.A(_03580_),
    .B(_06348_),
    .C(_06350_),
    .Y(_01126_));
 sky130_fd_sc_hd__a221oi_2 _21632_ (.A1(\csr._mcycle_T_2[10] ),
    .A2(_06325_),
    .B1(_06340_),
    .B2(_06349_),
    .C1(\csr.minstret[10] ),
    .Y(_06351_));
 sky130_fd_sc_hd__buf_1 _21633_ (.A(_03579_),
    .X(_06352_));
 sky130_fd_sc_hd__a211oi_2 _21634_ (.A1(\csr.minstret[10] ),
    .A2(_06350_),
    .B1(_06351_),
    .C1(_06352_),
    .Y(_01127_));
 sky130_fd_sc_hd__a221oi_2 _21635_ (.A1(\csr._mcycle_T_2[11] ),
    .A2(_06325_),
    .B1(_06350_),
    .B2(\csr.minstret[10] ),
    .C1(\csr.minstret[11] ),
    .Y(_06353_));
 sky130_fd_sc_hd__a311oi_2 _21636_ (.A1(\csr.minstret[10] ),
    .A2(\csr.minstret[11] ),
    .A3(_06350_),
    .B1(_06353_),
    .C1(_06336_),
    .Y(_01128_));
 sky130_fd_sc_hd__and3_2 _21637_ (.A(_05613_),
    .B(\csr.minstret[5] ),
    .C(\csr.minstret[10] ),
    .X(_06354_));
 sky130_fd_sc_hd__and3_2 _21638_ (.A(\csr.minstret[11] ),
    .B(_06349_),
    .C(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__a221oi_2 _21639_ (.A1(\csr._mcycle_T_2[12] ),
    .A2(_06325_),
    .B1(_06338_),
    .B2(_06355_),
    .C1(\csr.minstret[12] ),
    .Y(_06356_));
 sky130_fd_sc_hd__a311oi_2 _21640_ (.A1(\csr.minstret[12] ),
    .A2(_06338_),
    .A3(_06355_),
    .B1(_06356_),
    .C1(_06336_),
    .Y(_01129_));
 sky130_fd_sc_hd__a32o_2 _21641_ (.A1(\csr.minstret[12] ),
    .A2(_06338_),
    .A3(_06355_),
    .B1(_06329_),
    .B2(\csr._mcycle_T_2[13] ),
    .X(_06357_));
 sky130_fd_sc_hd__and3_2 _21642_ (.A(\csr.minstret[12] ),
    .B(_06338_),
    .C(_06355_),
    .X(_06358_));
 sky130_fd_sc_hd__nand2_2 _21643_ (.A(\csr.minstret[13] ),
    .B(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__o211a_2 _21644_ (.A1(\csr.minstret[13] ),
    .A2(_06357_),
    .B1(_06359_),
    .C1(_10546_),
    .X(_01130_));
 sky130_fd_sc_hd__and2_2 _21645_ (.A(\csr.minstret[12] ),
    .B(\csr.minstret[13] ),
    .X(_06360_));
 sky130_fd_sc_hd__and4_2 _21646_ (.A(\csr.minstret[10] ),
    .B(\csr.minstret[11] ),
    .C(_06349_),
    .D(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__and4_2 _21647_ (.A(\csr.minstret[4] ),
    .B(\csr.minstret[5] ),
    .C(\csr.minstret[14] ),
    .D(_06333_),
    .X(_06362_));
 sky130_fd_sc_hd__and3_2 _21648_ (.A(_06317_),
    .B(_06361_),
    .C(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__a221oi_2 _21649_ (.A1(\csr._mcycle_T_2[14] ),
    .A2(_06325_),
    .B1(_06358_),
    .B2(\csr.minstret[13] ),
    .C1(\csr.minstret[14] ),
    .Y(_06364_));
 sky130_fd_sc_hd__a211oi_2 _21650_ (.A1(\csr.io_inst_retired ),
    .A2(_06363_),
    .B1(_06364_),
    .C1(_06352_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand4_2 _21651_ (.A(\csr.minstret[14] ),
    .B(_06333_),
    .C(_06355_),
    .D(_06360_),
    .Y(_06365_));
 sky130_fd_sc_hd__nor3b_2 _21652_ (.A(_06320_),
    .B(_06365_),
    .C_N(\csr.io_inst_retired ),
    .Y(_06366_));
 sky130_fd_sc_hd__a211oi_2 _21653_ (.A1(\csr._mcycle_T_2[15] ),
    .A2(_06329_),
    .B1(_06366_),
    .C1(_05691_),
    .Y(_06367_));
 sky130_fd_sc_hd__a211oi_2 _21654_ (.A1(_05691_),
    .A2(_06366_),
    .B1(_06367_),
    .C1(_06352_),
    .Y(_01132_));
 sky130_fd_sc_hd__a221oi_2 _21655_ (.A1(\csr._mcycle_T_2[16] ),
    .A2(_06321_),
    .B1(_06366_),
    .B2(_05691_),
    .C1(\csr.minstret[16] ),
    .Y(_06368_));
 sky130_fd_sc_hd__and3_2 _21656_ (.A(_05691_),
    .B(\csr.minstret[16] ),
    .C(_06366_),
    .X(_06369_));
 sky130_fd_sc_hd__nor3_2 _21657_ (.A(_03580_),
    .B(_06368_),
    .C(_06369_),
    .Y(_01133_));
 sky130_fd_sc_hd__and4_2 _21658_ (.A(_05691_),
    .B(\csr.minstret[16] ),
    .C(\csr.io_inst_retired ),
    .D(_06363_),
    .X(_06370_));
 sky130_fd_sc_hd__a211o_2 _21659_ (.A1(\csr._mcycle_T_2[17] ),
    .A2(_06325_),
    .B1(_06370_),
    .C1(\csr.minstret[17] ),
    .X(_06371_));
 sky130_fd_sc_hd__nand2_2 _21660_ (.A(\csr.minstret[17] ),
    .B(_06370_),
    .Y(_06372_));
 sky130_fd_sc_hd__and3_2 _21661_ (.A(_10019_),
    .B(_06371_),
    .C(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__buf_1 _21662_ (.A(_06373_),
    .X(_01134_));
 sky130_fd_sc_hd__a21oi_2 _21663_ (.A1(\csr._mcycle_T_2[18] ),
    .A2(_06329_),
    .B1(\csr.minstret[18] ),
    .Y(_06374_));
 sky130_fd_sc_hd__and3_2 _21664_ (.A(\csr.minstret[17] ),
    .B(\csr.minstret[18] ),
    .C(_06370_),
    .X(_06375_));
 sky130_fd_sc_hd__a211oi_2 _21665_ (.A1(_06374_),
    .A2(_06372_),
    .B1(_06327_),
    .C1(_06375_),
    .Y(_01135_));
 sky130_fd_sc_hd__a211oi_2 _21666_ (.A1(\csr._mcycle_T_2[19] ),
    .A2(_06321_),
    .B1(_06375_),
    .C1(\csr.minstret[19] ),
    .Y(_06376_));
 sky130_fd_sc_hd__a211oi_2 _21667_ (.A1(\csr.minstret[19] ),
    .A2(_06375_),
    .B1(_06376_),
    .C1(_06352_),
    .Y(_01136_));
 sky130_fd_sc_hd__buf_1 _21668_ (.A(_03579_),
    .X(_06377_));
 sky130_fd_sc_hd__and4_2 _21669_ (.A(\csr.minstret[17] ),
    .B(\csr.minstret[18] ),
    .C(\csr.minstret[19] ),
    .D(_06369_),
    .X(_06378_));
 sky130_fd_sc_hd__a211oi_2 _21670_ (.A1(\csr._mcycle_T_2[20] ),
    .A2(_06329_),
    .B1(_06378_),
    .C1(\csr.minstret[20] ),
    .Y(_06379_));
 sky130_fd_sc_hd__and4_2 _21671_ (.A(\csr.minstret[17] ),
    .B(\csr.minstret[18] ),
    .C(\csr.minstret[19] ),
    .D(\csr.minstret[20] ),
    .X(_06380_));
 sky130_fd_sc_hd__and4_2 _21672_ (.A(_05691_),
    .B(\csr.minstret[16] ),
    .C(_06366_),
    .D(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__nor3_2 _21673_ (.A(_06377_),
    .B(_06379_),
    .C(_06381_),
    .Y(_01137_));
 sky130_fd_sc_hd__a211o_2 _21674_ (.A1(\csr._mcycle_T_2[21] ),
    .A2(_06320_),
    .B1(_06381_),
    .C1(\csr.minstret[21] ),
    .X(_06382_));
 sky130_fd_sc_hd__and3_2 _21675_ (.A(\csr.minstret[19] ),
    .B(\csr.minstret[20] ),
    .C(_06375_),
    .X(_06383_));
 sky130_fd_sc_hd__nand2_2 _21676_ (.A(\csr.minstret[21] ),
    .B(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__and3_2 _21677_ (.A(_10019_),
    .B(_06382_),
    .C(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__buf_1 _21678_ (.A(_06385_),
    .X(_01138_));
 sky130_fd_sc_hd__a21oi_2 _21679_ (.A1(\csr._mcycle_T_2[22] ),
    .A2(_06329_),
    .B1(\csr.minstret[22] ),
    .Y(_06386_));
 sky130_fd_sc_hd__and3_2 _21680_ (.A(\csr.minstret[21] ),
    .B(\csr.minstret[22] ),
    .C(_06381_),
    .X(_06387_));
 sky130_fd_sc_hd__a211oi_2 _21681_ (.A1(_06384_),
    .A2(_06386_),
    .B1(_06387_),
    .C1(_06352_),
    .Y(_01139_));
 sky130_fd_sc_hd__a211oi_2 _21682_ (.A1(\csr._mcycle_T_2[23] ),
    .A2(_06321_),
    .B1(_06387_),
    .C1(\csr.minstret[23] ),
    .Y(_06388_));
 sky130_fd_sc_hd__a211oi_2 _21683_ (.A1(\csr.minstret[23] ),
    .A2(_06387_),
    .B1(_06388_),
    .C1(_06352_),
    .Y(_01140_));
 sky130_fd_sc_hd__and4_2 _21684_ (.A(\csr.minstret[21] ),
    .B(\csr.minstret[22] ),
    .C(\csr.minstret[23] ),
    .D(_06383_),
    .X(_06389_));
 sky130_fd_sc_hd__a211oi_2 _21685_ (.A1(\csr._mcycle_T_2[24] ),
    .A2(_06329_),
    .B1(_06389_),
    .C1(\csr.minstret[24] ),
    .Y(_06390_));
 sky130_fd_sc_hd__and4_2 _21686_ (.A(\csr.minstret[21] ),
    .B(\csr.minstret[22] ),
    .C(\csr.minstret[23] ),
    .D(\csr.minstret[24] ),
    .X(_06391_));
 sky130_fd_sc_hd__and3_2 _21687_ (.A(_06369_),
    .B(_06380_),
    .C(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__nor3_2 _21688_ (.A(_06377_),
    .B(_06390_),
    .C(_06392_),
    .Y(_01141_));
 sky130_fd_sc_hd__a211oi_2 _21689_ (.A1(\csr._mcycle_T_2[25] ),
    .A2(_06321_),
    .B1(_06392_),
    .C1(\csr.minstret[25] ),
    .Y(_06393_));
 sky130_fd_sc_hd__a211oi_2 _21690_ (.A1(\csr.minstret[25] ),
    .A2(_06392_),
    .B1(_06393_),
    .C1(_06352_),
    .Y(_01142_));
 sky130_fd_sc_hd__a21o_2 _21691_ (.A1(\csr._mcycle_T_2[26] ),
    .A2(_06329_),
    .B1(\csr.minstret[26] ),
    .X(_06394_));
 sky130_fd_sc_hd__and3_2 _21692_ (.A(\csr.minstret[25] ),
    .B(_06381_),
    .C(_06391_),
    .X(_06395_));
 sky130_fd_sc_hd__buf_1 _21693_ (.A(_03449_),
    .X(_06396_));
 sky130_fd_sc_hd__and3_2 _21694_ (.A(_05691_),
    .B(\csr.minstret[16] ),
    .C(_06391_),
    .X(_06397_));
 sky130_fd_sc_hd__and4_2 _21695_ (.A(\csr.minstret[25] ),
    .B(\csr.minstret[26] ),
    .C(\csr.io_inst_retired ),
    .D(_06380_),
    .X(_06398_));
 sky130_fd_sc_hd__or4bb_2 _21696_ (.A(_06320_),
    .B(_06365_),
    .C_N(_06397_),
    .D_N(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__o211a_2 _21697_ (.A1(_06394_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06399_),
    .X(_01143_));
 sky130_fd_sc_hd__and3_2 _21698_ (.A(\csr.minstret[22] ),
    .B(\csr.minstret[23] ),
    .C(\csr.minstret[24] ),
    .X(_06400_));
 sky130_fd_sc_hd__and4_2 _21699_ (.A(\csr.minstret[16] ),
    .B(\csr.minstret[19] ),
    .C(\csr.minstret[20] ),
    .D(\csr.minstret[21] ),
    .X(_06401_));
 sky130_fd_sc_hd__and4_2 _21700_ (.A(\csr.minstret[17] ),
    .B(\csr.minstret[18] ),
    .C(_06400_),
    .D(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__and4_2 _21701_ (.A(\csr.minstret[15] ),
    .B(\csr.minstret[25] ),
    .C(\csr.minstret[26] ),
    .D(\csr.io_inst_retired ),
    .X(_06403_));
 sky130_fd_sc_hd__and3_2 _21702_ (.A(_06363_),
    .B(_06402_),
    .C(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__and3_2 _21703_ (.A(\csr.minstret[25] ),
    .B(\csr.minstret[26] ),
    .C(_06392_),
    .X(_06405_));
 sky130_fd_sc_hd__a211oi_2 _21704_ (.A1(\csr._mcycle_T_2[27] ),
    .A2(_06321_),
    .B1(_06405_),
    .C1(\csr.minstret[27] ),
    .Y(_06406_));
 sky130_fd_sc_hd__a211oi_2 _21705_ (.A1(\csr.minstret[27] ),
    .A2(_06404_),
    .B1(_06406_),
    .C1(_06352_),
    .Y(_01144_));
 sky130_fd_sc_hd__and4_2 _21706_ (.A(\csr.minstret[14] ),
    .B(_06333_),
    .C(_06355_),
    .D(_06360_),
    .X(_06407_));
 sky130_fd_sc_hd__and4_2 _21707_ (.A(_05691_),
    .B(\csr.minstret[16] ),
    .C(\csr.minstret[17] ),
    .D(\csr.minstret[18] ),
    .X(_06408_));
 sky130_fd_sc_hd__and4_2 _21708_ (.A(\csr.minstret[19] ),
    .B(\csr.minstret[26] ),
    .C(\csr.io_inst_retired ),
    .D(_06408_),
    .X(_06409_));
 sky130_fd_sc_hd__and3_2 _21709_ (.A(\csr.minstret[25] ),
    .B(_06407_),
    .C(_06409_),
    .X(_06410_));
 sky130_fd_sc_hd__and3_2 _21710_ (.A(\csr.minstret[20] ),
    .B(\csr.minstret[21] ),
    .C(\csr.minstret[22] ),
    .X(_06411_));
 sky130_fd_sc_hd__and3_2 _21711_ (.A(\csr.minstret[23] ),
    .B(\csr.minstret[24] ),
    .C(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__and4_2 _21712_ (.A(\csr.minstret[27] ),
    .B(_06410_),
    .C(_06317_),
    .D(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__a211oi_2 _21713_ (.A1(\csr._mcycle_T_2[28] ),
    .A2(_06321_),
    .B1(_06413_),
    .C1(\csr.minstret[28] ),
    .Y(_06414_));
 sky130_fd_sc_hd__a211oi_2 _21714_ (.A1(\csr.minstret[28] ),
    .A2(_06413_),
    .B1(_06414_),
    .C1(_06352_),
    .Y(_01145_));
 sky130_fd_sc_hd__and3_2 _21715_ (.A(\csr.minstret[27] ),
    .B(\csr.minstret[28] ),
    .C(_06404_),
    .X(_06415_));
 sky130_fd_sc_hd__a221oi_2 _21716_ (.A1(\csr._mcycle_T_2[29] ),
    .A2(_06325_),
    .B1(_06413_),
    .B2(\csr.minstret[28] ),
    .C1(\csr.minstret[29] ),
    .Y(_06416_));
 sky130_fd_sc_hd__a211oi_2 _21717_ (.A1(\csr.minstret[29] ),
    .A2(_06415_),
    .B1(_06416_),
    .C1(_06352_),
    .Y(_01146_));
 sky130_fd_sc_hd__and3_2 _21718_ (.A(\csr.minstret[28] ),
    .B(\csr.minstret[29] ),
    .C(_06413_),
    .X(_06417_));
 sky130_fd_sc_hd__a211oi_2 _21719_ (.A1(\csr._mcycle_T_2[30] ),
    .A2(_06321_),
    .B1(_06417_),
    .C1(\csr.minstret[30] ),
    .Y(_06418_));
 sky130_fd_sc_hd__buf_1 _21720_ (.A(_03579_),
    .X(_06419_));
 sky130_fd_sc_hd__a211oi_2 _21721_ (.A1(\csr.minstret[30] ),
    .A2(_06417_),
    .B1(_06418_),
    .C1(_06419_),
    .Y(_01147_));
 sky130_fd_sc_hd__and3_2 _21722_ (.A(\csr.minstret[29] ),
    .B(\csr.minstret[30] ),
    .C(_06415_),
    .X(_06420_));
 sky130_fd_sc_hd__a211oi_2 _21723_ (.A1(\csr._mcycle_T_2[31] ),
    .A2(_06321_),
    .B1(_06420_),
    .C1(\csr.minstret[31] ),
    .Y(_06421_));
 sky130_fd_sc_hd__a211oi_2 _21724_ (.A1(\csr.minstret[31] ),
    .A2(_06420_),
    .B1(_06421_),
    .C1(_06419_),
    .Y(_01148_));
 sky130_fd_sc_hd__buf_1 _21725_ (.A(_10576_),
    .X(_06422_));
 sky130_fd_sc_hd__a311oi_2 _21726_ (.A1(\csr.msie ),
    .A2(\csr.msip ),
    .A3(\csr.ie ),
    .B1(\execute.exception_out_reg ),
    .C1(_06031_),
    .Y(_06423_));
 sky130_fd_sc_hd__a31o_2 _21727_ (.A1(\csr.mtie ),
    .A2(\csr.ie ),
    .A3(\csr.mtip ),
    .B1(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__and4bb_2 _21728_ (.A_N(_06422_),
    .B_N(_09923_),
    .C(_06025_),
    .D(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__buf_1 _21729_ (.A(_06425_),
    .X(_01149_));
 sky130_fd_sc_hd__and3_2 _21730_ (.A(_09885_),
    .B(_09892_),
    .C(_09916_),
    .X(_06426_));
 sky130_fd_sc_hd__buf_1 _21731_ (.A(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__buf_1 _21732_ (.A(_06427_),
    .X(_06428_));
 sky130_fd_sc_hd__mux2_2 _21733_ (.A0(\fetch.bht.bhtTable_tag[4][0] ),
    .A1(_10820_),
    .S(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__buf_1 _21734_ (.A(_06429_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_2 _21735_ (.A0(\fetch.bht.bhtTable_tag[4][1] ),
    .A1(_10821_),
    .S(_06428_),
    .X(_06430_));
 sky130_fd_sc_hd__buf_1 _21736_ (.A(_06430_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_2 _21737_ (.A0(\fetch.bht.bhtTable_tag[4][2] ),
    .A1(_10881_),
    .S(_06428_),
    .X(_06431_));
 sky130_fd_sc_hd__buf_1 _21738_ (.A(_06431_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_2 _21739_ (.A0(\fetch.bht.bhtTable_tag[4][3] ),
    .A1(_10817_),
    .S(_06428_),
    .X(_06432_));
 sky130_fd_sc_hd__buf_1 _21740_ (.A(_06432_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_2 _21741_ (.A0(\fetch.bht.bhtTable_tag[4][4] ),
    .A1(_10878_),
    .S(_06428_),
    .X(_06433_));
 sky130_fd_sc_hd__buf_1 _21742_ (.A(_06433_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_2 _21743_ (.A0(\fetch.bht.bhtTable_tag[4][5] ),
    .A1(_10812_),
    .S(_06428_),
    .X(_06434_));
 sky130_fd_sc_hd__buf_1 _21744_ (.A(_06434_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_2 _21745_ (.A0(\fetch.bht.bhtTable_tag[4][6] ),
    .A1(\csr.io_mem_pc[12] ),
    .S(_06428_),
    .X(_06435_));
 sky130_fd_sc_hd__buf_1 _21746_ (.A(_06435_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_2 _21747_ (.A0(\fetch.bht.bhtTable_tag[4][7] ),
    .A1(_10871_),
    .S(_06428_),
    .X(_06436_));
 sky130_fd_sc_hd__buf_1 _21748_ (.A(_06436_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_2 _21749_ (.A0(\fetch.bht.bhtTable_tag[4][8] ),
    .A1(_10872_),
    .S(_06428_),
    .X(_06437_));
 sky130_fd_sc_hd__buf_1 _21750_ (.A(_06437_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_2 _21751_ (.A0(\fetch.bht.bhtTable_tag[4][9] ),
    .A1(_10807_),
    .S(_06428_),
    .X(_06438_));
 sky130_fd_sc_hd__buf_1 _21752_ (.A(_06438_),
    .X(_01159_));
 sky130_fd_sc_hd__buf_1 _21753_ (.A(_06427_),
    .X(_06439_));
 sky130_fd_sc_hd__mux2_2 _21754_ (.A0(\fetch.bht.bhtTable_tag[4][10] ),
    .A1(_10868_),
    .S(_06439_),
    .X(_06440_));
 sky130_fd_sc_hd__buf_1 _21755_ (.A(_06440_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_2 _21756_ (.A0(\fetch.bht.bhtTable_tag[4][11] ),
    .A1(_10803_),
    .S(_06439_),
    .X(_06441_));
 sky130_fd_sc_hd__buf_1 _21757_ (.A(_06441_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_2 _21758_ (.A0(\fetch.bht.bhtTable_tag[4][12] ),
    .A1(\csr.io_mem_pc[18] ),
    .S(_06439_),
    .X(_06442_));
 sky130_fd_sc_hd__buf_1 _21759_ (.A(_06442_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_2 _21760_ (.A0(\fetch.bht.bhtTable_tag[4][13] ),
    .A1(_10800_),
    .S(_06439_),
    .X(_06443_));
 sky130_fd_sc_hd__buf_1 _21761_ (.A(_06443_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_2 _21762_ (.A0(\fetch.bht.bhtTable_tag[4][14] ),
    .A1(_10795_),
    .S(_06439_),
    .X(_06444_));
 sky130_fd_sc_hd__buf_1 _21763_ (.A(_06444_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_2 _21764_ (.A0(\fetch.bht.bhtTable_tag[4][15] ),
    .A1(\csr.io_mem_pc[21] ),
    .S(_06439_),
    .X(_06445_));
 sky130_fd_sc_hd__buf_1 _21765_ (.A(_06445_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_2 _21766_ (.A0(\fetch.bht.bhtTable_tag[4][16] ),
    .A1(_10787_),
    .S(_06439_),
    .X(_06446_));
 sky130_fd_sc_hd__buf_1 _21767_ (.A(_06446_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_2 _21768_ (.A0(\fetch.bht.bhtTable_tag[4][17] ),
    .A1(\csr.io_mem_pc[23] ),
    .S(_06439_),
    .X(_06447_));
 sky130_fd_sc_hd__buf_1 _21769_ (.A(_06447_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_2 _21770_ (.A0(\fetch.bht.bhtTable_tag[4][18] ),
    .A1(_10772_),
    .S(_06439_),
    .X(_06448_));
 sky130_fd_sc_hd__buf_1 _21771_ (.A(_06448_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_2 _21772_ (.A0(\fetch.bht.bhtTable_tag[4][19] ),
    .A1(_10773_),
    .S(_06439_),
    .X(_06449_));
 sky130_fd_sc_hd__buf_1 _21773_ (.A(_06449_),
    .X(_01169_));
 sky130_fd_sc_hd__buf_1 _21774_ (.A(_06426_),
    .X(_06450_));
 sky130_fd_sc_hd__mux2_2 _21775_ (.A0(\fetch.bht.bhtTable_tag[4][20] ),
    .A1(_10760_),
    .S(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__buf_1 _21776_ (.A(_06451_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_2 _21777_ (.A0(\fetch.bht.bhtTable_tag[4][21] ),
    .A1(_10759_),
    .S(_06450_),
    .X(_06452_));
 sky130_fd_sc_hd__buf_1 _21778_ (.A(_06452_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_2 _21779_ (.A0(\fetch.bht.bhtTable_tag[4][22] ),
    .A1(_10771_),
    .S(_06450_),
    .X(_06453_));
 sky130_fd_sc_hd__buf_1 _21780_ (.A(_06453_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_2 _21781_ (.A0(\fetch.bht.bhtTable_tag[4][23] ),
    .A1(\csr.io_mem_pc[29] ),
    .S(_06450_),
    .X(_06454_));
 sky130_fd_sc_hd__buf_1 _21782_ (.A(_06454_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_2 _21783_ (.A0(\fetch.bht.bhtTable_tag[4][24] ),
    .A1(_10777_),
    .S(_06450_),
    .X(_06455_));
 sky130_fd_sc_hd__buf_1 _21784_ (.A(_06455_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_2 _21785_ (.A0(\fetch.bht.bhtTable_tag[4][25] ),
    .A1(\csr.io_mem_pc[31] ),
    .S(_06450_),
    .X(_06456_));
 sky130_fd_sc_hd__buf_1 _21786_ (.A(_06456_),
    .X(_01175_));
 sky130_fd_sc_hd__buf_1 _21787_ (.A(\csr.io_csr_write_address[0] ),
    .X(_06457_));
 sky130_fd_sc_hd__and4bb_2 _21788_ (.A_N(\csr.io_csr_write_address[10] ),
    .B_N(\csr.io_csr_write_address[11] ),
    .C(\csr.io_csr_write_address[9] ),
    .D(\csr.io_csr_write_address[8] ),
    .X(_06458_));
 sky130_fd_sc_hd__nor2_2 _21789_ (.A(\csr.io_csr_write_address[1] ),
    .B(_06315_),
    .Y(_06459_));
 sky130_fd_sc_hd__nand4b_2 _21790_ (.A_N(_06457_),
    .B(_06313_),
    .C(_06458_),
    .D(_06459_),
    .Y(_06460_));
 sky130_fd_sc_hd__inv_2 _21791_ (.A(_06037_),
    .Y(_06461_));
 sky130_fd_sc_hd__and2_2 _21792_ (.A(_06461_),
    .B(_10970_),
    .X(_06462_));
 sky130_fd_sc_hd__buf_1 _21793_ (.A(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__and4b_2 _21794_ (.A_N(_06457_),
    .B(_06313_),
    .C(_06458_),
    .D(_06459_),
    .X(_06464_));
 sky130_fd_sc_hd__a221o_2 _21795_ (.A1(\csr.ie ),
    .A2(_05857_),
    .B1(_06463_),
    .B2(\csr.pie ),
    .C1(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__o211a_2 _21796_ (.A1(_06460_),
    .A2(\csr._mcycle_T_2[3] ),
    .B1(_06396_),
    .C1(_06465_),
    .X(_01177_));
 sky130_fd_sc_hd__and4bb_2 _21797_ (.A_N(\csr.io_csr_write_address[1] ),
    .B_N(\csr.io_csr_write_address[3] ),
    .C(\csr.io_csr_write_address[2] ),
    .D(\csr.io_csr_write_enable ),
    .X(_06466_));
 sky130_fd_sc_hd__and4b_2 _21798_ (.A_N(_06457_),
    .B(_06313_),
    .C(_06458_),
    .D(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__or2b_2 _21799_ (.A(\csr._mcycle_T_2[7] ),
    .B_N(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__o211a_2 _21800_ (.A1(\csr.mtie ),
    .A2(_06467_),
    .B1(_06468_),
    .C1(_10546_),
    .X(_01178_));
 sky130_fd_sc_hd__nor3_2 _21801_ (.A(\csr.io_csr_write_address[5] ),
    .B(\csr.io_csr_write_address[4] ),
    .C(\csr.io_csr_write_address[7] ),
    .Y(_06469_));
 sky130_fd_sc_hd__and3_2 _21802_ (.A(\csr.io_csr_write_address[6] ),
    .B(_06469_),
    .C(_06458_),
    .X(_06470_));
 sky130_fd_sc_hd__and3b_2 _21803_ (.A_N(_06457_),
    .B(_06466_),
    .C(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__and3_2 _21804_ (.A(\csr.io_csr_write_address[6] ),
    .B(_06469_),
    .C(_06458_),
    .X(_06472_));
 sky130_fd_sc_hd__or4bb_2 _21805_ (.A(\csr._mcycle_T_2[3] ),
    .B(_06457_),
    .C_N(_06466_),
    .D_N(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__o211a_2 _21806_ (.A1(\csr.msip ),
    .A2(_06471_),
    .B1(_06473_),
    .C1(_10546_),
    .X(_01179_));
 sky130_fd_sc_hd__or2b_2 _21807_ (.A(\csr._mcycle_T_2[3] ),
    .B_N(_06467_),
    .X(_06474_));
 sky130_fd_sc_hd__o211a_2 _21808_ (.A1(\csr.msie ),
    .A2(_06467_),
    .B1(_06474_),
    .C1(_10546_),
    .X(_01180_));
 sky130_fd_sc_hd__or2b_2 _21809_ (.A(\csr._mcycle_T_2[11] ),
    .B_N(_06467_),
    .X(_06475_));
 sky130_fd_sc_hd__o211a_2 _21810_ (.A1(\csr.meie ),
    .A2(_06467_),
    .B1(_06475_),
    .C1(_10546_),
    .X(_01181_));
 sky130_fd_sc_hd__o22a_2 _21811_ (.A1(_06461_),
    .A2(\csr.ie ),
    .B1(\csr.pie ),
    .B2(_06032_),
    .X(_06476_));
 sky130_fd_sc_hd__mux2_2 _21812_ (.A0(\csr._mcycle_T_2[7] ),
    .A1(_06476_),
    .S(_06460_),
    .X(_06477_));
 sky130_fd_sc_hd__and2_2 _21813_ (.A(_06477_),
    .B(_10019_),
    .X(_06478_));
 sky130_fd_sc_hd__buf_1 _21814_ (.A(_06478_),
    .X(_01182_));
 sky130_fd_sc_hd__nand2_2 _21815_ (.A(_06316_),
    .B(_06472_),
    .Y(_06479_));
 sky130_fd_sc_hd__buf_1 _21816_ (.A(_06461_),
    .X(_06480_));
 sky130_fd_sc_hd__buf_1 _21817_ (.A(_06038_),
    .X(_06481_));
 sky130_fd_sc_hd__a22o_2 _21818_ (.A1(_06481_),
    .A2(\csr.io_interrupt ),
    .B1(_06316_),
    .B2(_06470_),
    .X(_06482_));
 sky130_fd_sc_hd__a21o_2 _21819_ (.A1(_06480_),
    .A2(\csr._csr_read_data_T_9[31] ),
    .B1(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__o211a_2 _21820_ (.A1(_06479_),
    .A2(\csr._mcycle_T_2[31] ),
    .B1(_06396_),
    .C1(_06483_),
    .X(_01183_));
 sky130_fd_sc_hd__a22o_2 _21821_ (.A1(_06481_),
    .A2(\csr.io_ecause[0] ),
    .B1(_06316_),
    .B2(_06470_),
    .X(_06484_));
 sky130_fd_sc_hd__a21o_2 _21822_ (.A1(_06480_),
    .A2(\csr._csr_read_data_T_9[0] ),
    .B1(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__o211a_2 _21823_ (.A1(_06479_),
    .A2(\csr._mcycle_T_2[0] ),
    .B1(_06396_),
    .C1(_06485_),
    .X(_01184_));
 sky130_fd_sc_hd__a22o_2 _21824_ (.A1(_06481_),
    .A2(\csr.io_ecause[1] ),
    .B1(_06316_),
    .B2(_06470_),
    .X(_06486_));
 sky130_fd_sc_hd__a21o_2 _21825_ (.A1(_06480_),
    .A2(\csr._csr_read_data_T_9[1] ),
    .B1(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__o211a_2 _21826_ (.A1(_06479_),
    .A2(\csr._mcycle_T_2[1] ),
    .B1(_06396_),
    .C1(_06487_),
    .X(_01185_));
 sky130_fd_sc_hd__a22o_2 _21827_ (.A1(_06481_),
    .A2(\csr.io_ecause[2] ),
    .B1(_06316_),
    .B2(_06470_),
    .X(_06488_));
 sky130_fd_sc_hd__a21o_2 _21828_ (.A1(_06480_),
    .A2(\csr._csr_read_data_T_9[2] ),
    .B1(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__o211a_2 _21829_ (.A1(_06479_),
    .A2(\csr._mcycle_T_2[2] ),
    .B1(_06396_),
    .C1(_06489_),
    .X(_01186_));
 sky130_fd_sc_hd__a22o_2 _21830_ (.A1(_06480_),
    .A2(\csr._csr_read_data_T_9[3] ),
    .B1(_06316_),
    .B2(_06472_),
    .X(_06490_));
 sky130_fd_sc_hd__o211a_2 _21831_ (.A1(_06479_),
    .A2(\csr._mcycle_T_2[3] ),
    .B1(_06396_),
    .C1(_06490_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_2 _21832_ (.A0(\csr.io_mret_vector[0] ),
    .A1(\csr.io_mem_pc[0] ),
    .S(_06040_),
    .X(_06491_));
 sky130_fd_sc_hd__and3_2 _21833_ (.A(_06457_),
    .B(_06459_),
    .C(_06472_),
    .X(_06492_));
 sky130_fd_sc_hd__buf_1 _21834_ (.A(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__buf_1 _21835_ (.A(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__buf_1 _21836_ (.A(_03449_),
    .X(_06495_));
 sky130_fd_sc_hd__or4bb_2 _21837_ (.A(_06315_),
    .B(\csr.io_csr_write_address[1] ),
    .C_N(\csr.io_csr_write_address[0] ),
    .D_N(_06472_),
    .X(_06496_));
 sky130_fd_sc_hd__buf_1 _21838_ (.A(_06496_),
    .X(_06497_));
 sky130_fd_sc_hd__or2_2 _21839_ (.A(\csr._mcycle_T_2[0] ),
    .B(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__o211a_2 _21840_ (.A1(_06491_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06498_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_2 _21841_ (.A0(\csr.io_mret_vector[1] ),
    .A1(\csr.io_mem_pc[1] ),
    .S(_06040_),
    .X(_06499_));
 sky130_fd_sc_hd__or2_2 _21842_ (.A(\csr._mcycle_T_2[1] ),
    .B(_06497_),
    .X(_06500_));
 sky130_fd_sc_hd__o211a_2 _21843_ (.A1(_06499_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06500_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_2 _21844_ (.A0(\csr.io_mret_vector[2] ),
    .A1(_10556_),
    .S(_06040_),
    .X(_06501_));
 sky130_fd_sc_hd__or2_2 _21845_ (.A(\csr._mcycle_T_2[2] ),
    .B(_06497_),
    .X(_06502_));
 sky130_fd_sc_hd__o211a_2 _21846_ (.A1(_06501_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06502_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_2 _21847_ (.A0(\csr.io_mret_vector[3] ),
    .A1(_10557_),
    .S(_06040_),
    .X(_06503_));
 sky130_fd_sc_hd__or2_2 _21848_ (.A(\csr._mcycle_T_2[3] ),
    .B(_06497_),
    .X(_06504_));
 sky130_fd_sc_hd__o211a_2 _21849_ (.A1(_06503_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06504_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_2 _21850_ (.A0(\csr.io_mret_vector[4] ),
    .A1(_09881_),
    .S(_06040_),
    .X(_06505_));
 sky130_fd_sc_hd__or2_2 _21851_ (.A(\csr._mcycle_T_2[4] ),
    .B(_06497_),
    .X(_06506_));
 sky130_fd_sc_hd__o211a_2 _21852_ (.A1(_06505_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06506_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_2 _21853_ (.A0(\csr.io_mret_vector[5] ),
    .A1(_09884_),
    .S(_06040_),
    .X(_06507_));
 sky130_fd_sc_hd__or2_2 _21854_ (.A(\csr._mcycle_T_2[5] ),
    .B(_06497_),
    .X(_06508_));
 sky130_fd_sc_hd__o211a_2 _21855_ (.A1(_06507_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06508_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_2 _21856_ (.A0(\csr.io_mret_vector[6] ),
    .A1(_10820_),
    .S(_06040_),
    .X(_06509_));
 sky130_fd_sc_hd__or2_2 _21857_ (.A(\csr._mcycle_T_2[6] ),
    .B(_06497_),
    .X(_06510_));
 sky130_fd_sc_hd__o211a_2 _21858_ (.A1(_06509_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06510_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_2 _21859_ (.A0(\csr.io_mret_vector[7] ),
    .A1(_10821_),
    .S(_06040_),
    .X(_06511_));
 sky130_fd_sc_hd__or2_2 _21860_ (.A(\csr._mcycle_T_2[7] ),
    .B(_06497_),
    .X(_06512_));
 sky130_fd_sc_hd__o211a_2 _21861_ (.A1(_06511_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06512_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_2 _21862_ (.A0(\csr.io_mret_vector[8] ),
    .A1(_10881_),
    .S(_06040_),
    .X(_06513_));
 sky130_fd_sc_hd__or2_2 _21863_ (.A(\csr._mcycle_T_2[8] ),
    .B(_06497_),
    .X(_06514_));
 sky130_fd_sc_hd__o211a_2 _21864_ (.A1(_06513_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06514_),
    .X(_01196_));
 sky130_fd_sc_hd__buf_1 _21865_ (.A(_06039_),
    .X(_06515_));
 sky130_fd_sc_hd__mux2_2 _21866_ (.A0(\csr.io_mret_vector[9] ),
    .A1(_10817_),
    .S(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__or2_2 _21867_ (.A(\csr._mcycle_T_2[9] ),
    .B(_06497_),
    .X(_06517_));
 sky130_fd_sc_hd__o211a_2 _21868_ (.A1(_06516_),
    .A2(_06494_),
    .B1(_06495_),
    .C1(_06517_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_2 _21869_ (.A0(\csr.io_mret_vector[10] ),
    .A1(_10878_),
    .S(_06515_),
    .X(_06518_));
 sky130_fd_sc_hd__buf_1 _21870_ (.A(_06493_),
    .X(_06519_));
 sky130_fd_sc_hd__buf_1 _21871_ (.A(_03449_),
    .X(_06520_));
 sky130_fd_sc_hd__buf_1 _21872_ (.A(_06496_),
    .X(_06521_));
 sky130_fd_sc_hd__or2_2 _21873_ (.A(\csr._mcycle_T_2[10] ),
    .B(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__o211a_2 _21874_ (.A1(_06518_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06522_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_2 _21875_ (.A0(\csr.io_mret_vector[11] ),
    .A1(_10812_),
    .S(_06515_),
    .X(_06523_));
 sky130_fd_sc_hd__or2_2 _21876_ (.A(\csr._mcycle_T_2[11] ),
    .B(_06521_),
    .X(_06524_));
 sky130_fd_sc_hd__o211a_2 _21877_ (.A1(_06523_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06524_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_2 _21878_ (.A0(\csr.io_mret_vector[12] ),
    .A1(\csr.io_mem_pc[12] ),
    .S(_06515_),
    .X(_06525_));
 sky130_fd_sc_hd__or2_2 _21879_ (.A(\csr._mcycle_T_2[12] ),
    .B(_06521_),
    .X(_06526_));
 sky130_fd_sc_hd__o211a_2 _21880_ (.A1(_06525_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06526_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_2 _21881_ (.A0(\csr.io_mret_vector[13] ),
    .A1(_10871_),
    .S(_06515_),
    .X(_06527_));
 sky130_fd_sc_hd__or2_2 _21882_ (.A(\csr._mcycle_T_2[13] ),
    .B(_06521_),
    .X(_06528_));
 sky130_fd_sc_hd__o211a_2 _21883_ (.A1(_06527_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06528_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_2 _21884_ (.A0(\csr.io_mret_vector[14] ),
    .A1(_10872_),
    .S(_06515_),
    .X(_06529_));
 sky130_fd_sc_hd__or2_2 _21885_ (.A(\csr._mcycle_T_2[14] ),
    .B(_06521_),
    .X(_06530_));
 sky130_fd_sc_hd__o211a_2 _21886_ (.A1(_06529_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06530_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_2 _21887_ (.A0(\csr.io_mret_vector[15] ),
    .A1(_10807_),
    .S(_06515_),
    .X(_06531_));
 sky130_fd_sc_hd__or2_2 _21888_ (.A(\csr._mcycle_T_2[15] ),
    .B(_06521_),
    .X(_06532_));
 sky130_fd_sc_hd__o211a_2 _21889_ (.A1(_06531_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06532_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_2 _21890_ (.A0(\csr.io_mret_vector[16] ),
    .A1(_10868_),
    .S(_06515_),
    .X(_06533_));
 sky130_fd_sc_hd__or2_2 _21891_ (.A(\csr._mcycle_T_2[16] ),
    .B(_06521_),
    .X(_06534_));
 sky130_fd_sc_hd__o211a_2 _21892_ (.A1(_06533_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06534_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_2 _21893_ (.A0(\csr.io_mret_vector[17] ),
    .A1(_10803_),
    .S(_06515_),
    .X(_06535_));
 sky130_fd_sc_hd__or2_2 _21894_ (.A(\csr._mcycle_T_2[17] ),
    .B(_06521_),
    .X(_06536_));
 sky130_fd_sc_hd__o211a_2 _21895_ (.A1(_06535_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06536_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_2 _21896_ (.A0(\csr.io_mret_vector[18] ),
    .A1(\csr.io_mem_pc[18] ),
    .S(_06515_),
    .X(_06537_));
 sky130_fd_sc_hd__or2_2 _21897_ (.A(\csr._mcycle_T_2[18] ),
    .B(_06521_),
    .X(_06538_));
 sky130_fd_sc_hd__o211a_2 _21898_ (.A1(_06537_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06538_),
    .X(_01206_));
 sky130_fd_sc_hd__buf_1 _21899_ (.A(_06039_),
    .X(_06539_));
 sky130_fd_sc_hd__mux2_2 _21900_ (.A0(\csr.io_mret_vector[19] ),
    .A1(_10800_),
    .S(_06539_),
    .X(_06540_));
 sky130_fd_sc_hd__or2_2 _21901_ (.A(\csr._mcycle_T_2[19] ),
    .B(_06521_),
    .X(_06541_));
 sky130_fd_sc_hd__o211a_2 _21902_ (.A1(_06540_),
    .A2(_06519_),
    .B1(_06520_),
    .C1(_06541_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_2 _21903_ (.A0(\csr.io_mret_vector[20] ),
    .A1(_10795_),
    .S(_06539_),
    .X(_06542_));
 sky130_fd_sc_hd__buf_1 _21904_ (.A(_06493_),
    .X(_06543_));
 sky130_fd_sc_hd__buf_1 _21905_ (.A(_03449_),
    .X(_06544_));
 sky130_fd_sc_hd__buf_1 _21906_ (.A(_06496_),
    .X(_06545_));
 sky130_fd_sc_hd__or2_2 _21907_ (.A(\csr._mcycle_T_2[20] ),
    .B(_06545_),
    .X(_06546_));
 sky130_fd_sc_hd__o211a_2 _21908_ (.A1(_06542_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06546_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_2 _21909_ (.A0(\csr.io_mret_vector[21] ),
    .A1(\csr.io_mem_pc[21] ),
    .S(_06539_),
    .X(_06547_));
 sky130_fd_sc_hd__or2_2 _21910_ (.A(\csr._mcycle_T_2[21] ),
    .B(_06545_),
    .X(_06548_));
 sky130_fd_sc_hd__o211a_2 _21911_ (.A1(_06547_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06548_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_2 _21912_ (.A0(\csr.io_mret_vector[22] ),
    .A1(_10787_),
    .S(_06539_),
    .X(_06549_));
 sky130_fd_sc_hd__or2_2 _21913_ (.A(\csr._mcycle_T_2[22] ),
    .B(_06545_),
    .X(_06550_));
 sky130_fd_sc_hd__o211a_2 _21914_ (.A1(_06549_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06550_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_2 _21915_ (.A0(\csr.io_mret_vector[23] ),
    .A1(\csr.io_mem_pc[23] ),
    .S(_06539_),
    .X(_06551_));
 sky130_fd_sc_hd__or2_2 _21916_ (.A(\csr._mcycle_T_2[23] ),
    .B(_06545_),
    .X(_06552_));
 sky130_fd_sc_hd__o211a_2 _21917_ (.A1(_06551_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06552_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_2 _21918_ (.A0(\csr.io_mret_vector[24] ),
    .A1(_10772_),
    .S(_06539_),
    .X(_06553_));
 sky130_fd_sc_hd__or2_2 _21919_ (.A(\csr._mcycle_T_2[24] ),
    .B(_06545_),
    .X(_06554_));
 sky130_fd_sc_hd__o211a_2 _21920_ (.A1(_06553_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06554_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_2 _21921_ (.A0(\csr.io_mret_vector[25] ),
    .A1(_10773_),
    .S(_06539_),
    .X(_06555_));
 sky130_fd_sc_hd__or2_2 _21922_ (.A(\csr._mcycle_T_2[25] ),
    .B(_06545_),
    .X(_06556_));
 sky130_fd_sc_hd__o211a_2 _21923_ (.A1(_06555_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06556_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_2 _21924_ (.A0(\csr.io_mret_vector[26] ),
    .A1(_10760_),
    .S(_06539_),
    .X(_06557_));
 sky130_fd_sc_hd__or2_2 _21925_ (.A(\csr._mcycle_T_2[26] ),
    .B(_06545_),
    .X(_06558_));
 sky130_fd_sc_hd__o211a_2 _21926_ (.A1(_06557_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06558_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_2 _21927_ (.A0(\csr.io_mret_vector[27] ),
    .A1(_10759_),
    .S(_06539_),
    .X(_06559_));
 sky130_fd_sc_hd__or2_2 _21928_ (.A(\csr._mcycle_T_2[27] ),
    .B(_06545_),
    .X(_06560_));
 sky130_fd_sc_hd__o211a_2 _21929_ (.A1(_06559_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06560_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_2 _21930_ (.A0(\csr.io_mret_vector[28] ),
    .A1(_10771_),
    .S(_06539_),
    .X(_06561_));
 sky130_fd_sc_hd__or2_2 _21931_ (.A(\csr._mcycle_T_2[28] ),
    .B(_06545_),
    .X(_06562_));
 sky130_fd_sc_hd__o211a_2 _21932_ (.A1(_06561_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06562_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_2 _21933_ (.A0(\csr.io_mret_vector[29] ),
    .A1(\csr.io_mem_pc[29] ),
    .S(_06481_),
    .X(_06563_));
 sky130_fd_sc_hd__or2_2 _21934_ (.A(\csr._mcycle_T_2[29] ),
    .B(_06545_),
    .X(_06564_));
 sky130_fd_sc_hd__o211a_2 _21935_ (.A1(_06563_),
    .A2(_06543_),
    .B1(_06544_),
    .C1(_06564_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_2 _21936_ (.A0(\csr.io_mret_vector[30] ),
    .A1(_10777_),
    .S(_06481_),
    .X(_06565_));
 sky130_fd_sc_hd__buf_1 _21937_ (.A(_03449_),
    .X(_06566_));
 sky130_fd_sc_hd__or2_2 _21938_ (.A(\csr._mcycle_T_2[30] ),
    .B(_06496_),
    .X(_06567_));
 sky130_fd_sc_hd__o211a_2 _21939_ (.A1(_06565_),
    .A2(_06493_),
    .B1(_06566_),
    .C1(_06567_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_2 _21940_ (.A0(\csr.io_mret_vector[31] ),
    .A1(\csr.io_mem_pc[31] ),
    .S(_06481_),
    .X(_06568_));
 sky130_fd_sc_hd__or2_2 _21941_ (.A(\csr._mcycle_T_2[31] ),
    .B(_06496_),
    .X(_06569_));
 sky130_fd_sc_hd__o211a_2 _21942_ (.A1(_06568_),
    .A2(_06493_),
    .B1(_06566_),
    .C1(_06569_),
    .X(_01219_));
 sky130_fd_sc_hd__or4b_2 _21943_ (.A(\csr.io_csr_write_address[1] ),
    .B(_06457_),
    .C(_06315_),
    .D_N(_06470_),
    .X(_06570_));
 sky130_fd_sc_hd__buf_1 _21944_ (.A(_06570_),
    .X(_06571_));
 sky130_fd_sc_hd__buf_1 _21945_ (.A(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__and3b_2 _21946_ (.A_N(_06457_),
    .B(_06459_),
    .C(_06470_),
    .X(_06573_));
 sky130_fd_sc_hd__buf_1 _21947_ (.A(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__or2_2 _21948_ (.A(\csr.mscratch[0] ),
    .B(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__o211a_2 _21949_ (.A1(\csr._mcycle_T_2[0] ),
    .A2(_06572_),
    .B1(_06575_),
    .C1(_10546_),
    .X(_01220_));
 sky130_fd_sc_hd__or2_2 _21950_ (.A(\csr.mscratch[1] ),
    .B(_06574_),
    .X(_06576_));
 sky130_fd_sc_hd__o211a_2 _21951_ (.A1(\csr._mcycle_T_2[1] ),
    .A2(_06572_),
    .B1(_06576_),
    .C1(_10546_),
    .X(_01221_));
 sky130_fd_sc_hd__or2_2 _21952_ (.A(\csr.mscratch[2] ),
    .B(_06574_),
    .X(_06577_));
 sky130_fd_sc_hd__buf_1 _21953_ (.A(_10130_),
    .X(_06578_));
 sky130_fd_sc_hd__buf_1 _21954_ (.A(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__o211a_2 _21955_ (.A1(\csr._mcycle_T_2[2] ),
    .A2(_06572_),
    .B1(_06577_),
    .C1(_06579_),
    .X(_01222_));
 sky130_fd_sc_hd__or2_2 _21956_ (.A(\csr.mscratch[3] ),
    .B(_06574_),
    .X(_06580_));
 sky130_fd_sc_hd__o211a_2 _21957_ (.A1(\csr._mcycle_T_2[3] ),
    .A2(_06572_),
    .B1(_06580_),
    .C1(_06579_),
    .X(_01223_));
 sky130_fd_sc_hd__or2_2 _21958_ (.A(\csr.mscratch[4] ),
    .B(_06574_),
    .X(_06581_));
 sky130_fd_sc_hd__o211a_2 _21959_ (.A1(\csr._mcycle_T_2[4] ),
    .A2(_06572_),
    .B1(_06581_),
    .C1(_06579_),
    .X(_01224_));
 sky130_fd_sc_hd__or2_2 _21960_ (.A(\csr.mscratch[5] ),
    .B(_06574_),
    .X(_06582_));
 sky130_fd_sc_hd__o211a_2 _21961_ (.A1(\csr._mcycle_T_2[5] ),
    .A2(_06572_),
    .B1(_06582_),
    .C1(_06579_),
    .X(_01225_));
 sky130_fd_sc_hd__or2_2 _21962_ (.A(\csr.mscratch[6] ),
    .B(_06574_),
    .X(_06583_));
 sky130_fd_sc_hd__o211a_2 _21963_ (.A1(\csr._mcycle_T_2[6] ),
    .A2(_06572_),
    .B1(_06583_),
    .C1(_06579_),
    .X(_01226_));
 sky130_fd_sc_hd__or2_2 _21964_ (.A(\csr.mscratch[7] ),
    .B(_06574_),
    .X(_06584_));
 sky130_fd_sc_hd__o211a_2 _21965_ (.A1(\csr._mcycle_T_2[7] ),
    .A2(_06572_),
    .B1(_06584_),
    .C1(_06579_),
    .X(_01227_));
 sky130_fd_sc_hd__or2_2 _21966_ (.A(\csr.mscratch[8] ),
    .B(_06574_),
    .X(_06585_));
 sky130_fd_sc_hd__o211a_2 _21967_ (.A1(\csr._mcycle_T_2[8] ),
    .A2(_06572_),
    .B1(_06585_),
    .C1(_06579_),
    .X(_01228_));
 sky130_fd_sc_hd__or2_2 _21968_ (.A(\csr.mscratch[9] ),
    .B(_06574_),
    .X(_06586_));
 sky130_fd_sc_hd__o211a_2 _21969_ (.A1(\csr._mcycle_T_2[9] ),
    .A2(_06572_),
    .B1(_06586_),
    .C1(_06579_),
    .X(_01229_));
 sky130_fd_sc_hd__buf_1 _21970_ (.A(_06571_),
    .X(_06587_));
 sky130_fd_sc_hd__buf_1 _21971_ (.A(_06573_),
    .X(_06588_));
 sky130_fd_sc_hd__or2_2 _21972_ (.A(\csr.mscratch[10] ),
    .B(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__o211a_2 _21973_ (.A1(\csr._mcycle_T_2[10] ),
    .A2(_06587_),
    .B1(_06589_),
    .C1(_06579_),
    .X(_01230_));
 sky130_fd_sc_hd__or2_2 _21974_ (.A(\csr.mscratch[11] ),
    .B(_06588_),
    .X(_06590_));
 sky130_fd_sc_hd__o211a_2 _21975_ (.A1(\csr._mcycle_T_2[11] ),
    .A2(_06587_),
    .B1(_06590_),
    .C1(_06579_),
    .X(_01231_));
 sky130_fd_sc_hd__or2_2 _21976_ (.A(\csr.mscratch[12] ),
    .B(_06588_),
    .X(_06591_));
 sky130_fd_sc_hd__buf_1 _21977_ (.A(_06578_),
    .X(_06592_));
 sky130_fd_sc_hd__o211a_2 _21978_ (.A1(\csr._mcycle_T_2[12] ),
    .A2(_06587_),
    .B1(_06591_),
    .C1(_06592_),
    .X(_01232_));
 sky130_fd_sc_hd__or2_2 _21979_ (.A(\csr.mscratch[13] ),
    .B(_06588_),
    .X(_06593_));
 sky130_fd_sc_hd__o211a_2 _21980_ (.A1(\csr._mcycle_T_2[13] ),
    .A2(_06587_),
    .B1(_06593_),
    .C1(_06592_),
    .X(_01233_));
 sky130_fd_sc_hd__or2_2 _21981_ (.A(\csr.mscratch[14] ),
    .B(_06588_),
    .X(_06594_));
 sky130_fd_sc_hd__o211a_2 _21982_ (.A1(\csr._mcycle_T_2[14] ),
    .A2(_06587_),
    .B1(_06594_),
    .C1(_06592_),
    .X(_01234_));
 sky130_fd_sc_hd__or2_2 _21983_ (.A(\csr.mscratch[15] ),
    .B(_06588_),
    .X(_06595_));
 sky130_fd_sc_hd__o211a_2 _21984_ (.A1(\csr._mcycle_T_2[15] ),
    .A2(_06587_),
    .B1(_06595_),
    .C1(_06592_),
    .X(_01235_));
 sky130_fd_sc_hd__or2_2 _21985_ (.A(\csr.mscratch[16] ),
    .B(_06588_),
    .X(_06596_));
 sky130_fd_sc_hd__o211a_2 _21986_ (.A1(\csr._mcycle_T_2[16] ),
    .A2(_06587_),
    .B1(_06596_),
    .C1(_06592_),
    .X(_01236_));
 sky130_fd_sc_hd__or2_2 _21987_ (.A(\csr.mscratch[17] ),
    .B(_06588_),
    .X(_06597_));
 sky130_fd_sc_hd__o211a_2 _21988_ (.A1(\csr._mcycle_T_2[17] ),
    .A2(_06587_),
    .B1(_06597_),
    .C1(_06592_),
    .X(_01237_));
 sky130_fd_sc_hd__or2_2 _21989_ (.A(\csr.mscratch[18] ),
    .B(_06588_),
    .X(_06598_));
 sky130_fd_sc_hd__o211a_2 _21990_ (.A1(\csr._mcycle_T_2[18] ),
    .A2(_06587_),
    .B1(_06598_),
    .C1(_06592_),
    .X(_01238_));
 sky130_fd_sc_hd__or2_2 _21991_ (.A(\csr.mscratch[19] ),
    .B(_06588_),
    .X(_06599_));
 sky130_fd_sc_hd__o211a_2 _21992_ (.A1(\csr._mcycle_T_2[19] ),
    .A2(_06587_),
    .B1(_06599_),
    .C1(_06592_),
    .X(_01239_));
 sky130_fd_sc_hd__buf_1 _21993_ (.A(_06571_),
    .X(_06600_));
 sky130_fd_sc_hd__buf_1 _21994_ (.A(_06573_),
    .X(_06601_));
 sky130_fd_sc_hd__or2_2 _21995_ (.A(\csr.mscratch[20] ),
    .B(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__o211a_2 _21996_ (.A1(\csr._mcycle_T_2[20] ),
    .A2(_06600_),
    .B1(_06602_),
    .C1(_06592_),
    .X(_01240_));
 sky130_fd_sc_hd__or2_2 _21997_ (.A(\csr.mscratch[21] ),
    .B(_06601_),
    .X(_06603_));
 sky130_fd_sc_hd__o211a_2 _21998_ (.A1(\csr._mcycle_T_2[21] ),
    .A2(_06600_),
    .B1(_06603_),
    .C1(_06592_),
    .X(_01241_));
 sky130_fd_sc_hd__or2_2 _21999_ (.A(\csr.mscratch[22] ),
    .B(_06601_),
    .X(_06604_));
 sky130_fd_sc_hd__buf_1 _22000_ (.A(_06578_),
    .X(_06605_));
 sky130_fd_sc_hd__o211a_2 _22001_ (.A1(\csr._mcycle_T_2[22] ),
    .A2(_06600_),
    .B1(_06604_),
    .C1(_06605_),
    .X(_01242_));
 sky130_fd_sc_hd__or2_2 _22002_ (.A(\csr.mscratch[23] ),
    .B(_06601_),
    .X(_06606_));
 sky130_fd_sc_hd__o211a_2 _22003_ (.A1(\csr._mcycle_T_2[23] ),
    .A2(_06600_),
    .B1(_06606_),
    .C1(_06605_),
    .X(_01243_));
 sky130_fd_sc_hd__or2_2 _22004_ (.A(\csr.mscratch[24] ),
    .B(_06601_),
    .X(_06607_));
 sky130_fd_sc_hd__o211a_2 _22005_ (.A1(\csr._mcycle_T_2[24] ),
    .A2(_06600_),
    .B1(_06607_),
    .C1(_06605_),
    .X(_01244_));
 sky130_fd_sc_hd__or2_2 _22006_ (.A(\csr.mscratch[25] ),
    .B(_06601_),
    .X(_06608_));
 sky130_fd_sc_hd__o211a_2 _22007_ (.A1(\csr._mcycle_T_2[25] ),
    .A2(_06600_),
    .B1(_06608_),
    .C1(_06605_),
    .X(_01245_));
 sky130_fd_sc_hd__or2_2 _22008_ (.A(\csr.mscratch[26] ),
    .B(_06601_),
    .X(_06609_));
 sky130_fd_sc_hd__o211a_2 _22009_ (.A1(\csr._mcycle_T_2[26] ),
    .A2(_06600_),
    .B1(_06609_),
    .C1(_06605_),
    .X(_01246_));
 sky130_fd_sc_hd__or2_2 _22010_ (.A(\csr.mscratch[27] ),
    .B(_06601_),
    .X(_06610_));
 sky130_fd_sc_hd__o211a_2 _22011_ (.A1(\csr._mcycle_T_2[27] ),
    .A2(_06600_),
    .B1(_06610_),
    .C1(_06605_),
    .X(_01247_));
 sky130_fd_sc_hd__or2_2 _22012_ (.A(\csr.mscratch[28] ),
    .B(_06601_),
    .X(_06611_));
 sky130_fd_sc_hd__o211a_2 _22013_ (.A1(\csr._mcycle_T_2[28] ),
    .A2(_06600_),
    .B1(_06611_),
    .C1(_06605_),
    .X(_01248_));
 sky130_fd_sc_hd__or2_2 _22014_ (.A(\csr.mscratch[29] ),
    .B(_06601_),
    .X(_06612_));
 sky130_fd_sc_hd__o211a_2 _22015_ (.A1(\csr._mcycle_T_2[29] ),
    .A2(_06600_),
    .B1(_06612_),
    .C1(_06605_),
    .X(_01249_));
 sky130_fd_sc_hd__or2_2 _22016_ (.A(\csr.mscratch[30] ),
    .B(_06573_),
    .X(_06613_));
 sky130_fd_sc_hd__o211a_2 _22017_ (.A1(\csr._mcycle_T_2[30] ),
    .A2(_06571_),
    .B1(_06613_),
    .C1(_06605_),
    .X(_01250_));
 sky130_fd_sc_hd__or2_2 _22018_ (.A(\csr.mscratch[31] ),
    .B(_06573_),
    .X(_06614_));
 sky130_fd_sc_hd__o211a_2 _22019_ (.A1(\csr._mcycle_T_2[31] ),
    .A2(_06571_),
    .B1(_06614_),
    .C1(_06605_),
    .X(_01251_));
 sky130_fd_sc_hd__buf_1 _22020_ (.A(_00000_),
    .X(_06615_));
 sky130_fd_sc_hd__buf_1 _22021_ (.A(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__buf_1 _22022_ (.A(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__buf_1 _22023_ (.A(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__buf_1 _22024_ (.A(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__buf_1 _22025_ (.A(_00001_),
    .X(_06620_));
 sky130_fd_sc_hd__buf_1 _22026_ (.A(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__buf_1 _22027_ (.A(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__buf_1 _22028_ (.A(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__buf_1 _22029_ (.A(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__mux4_2 _22030_ (.A0(\fetch.bht.bhtTable_tag[8][22] ),
    .A1(\fetch.bht.bhtTable_tag[9][22] ),
    .A2(\fetch.bht.bhtTable_tag[10][22] ),
    .A3(\fetch.bht.bhtTable_tag[11][22] ),
    .S0(_06619_),
    .S1(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__inv_2 _22031_ (.A(_00002_),
    .Y(_06626_));
 sky130_fd_sc_hd__buf_1 _22032_ (.A(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__buf_1 _22033_ (.A(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__buf_1 _22034_ (.A(_06628_),
    .X(_06629_));
 sky130_fd_sc_hd__and2_2 _22035_ (.A(_06625_),
    .B(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__buf_1 _22036_ (.A(_00002_),
    .X(_06631_));
 sky130_fd_sc_hd__buf_1 _22037_ (.A(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__buf_1 _22038_ (.A(_06632_),
    .X(_06633_));
 sky130_fd_sc_hd__mux4_2 _22039_ (.A0(\fetch.bht.bhtTable_tag[12][22] ),
    .A1(\fetch.bht.bhtTable_tag[13][22] ),
    .A2(\fetch.bht.bhtTable_tag[14][22] ),
    .A3(\fetch.bht.bhtTable_tag[15][22] ),
    .S0(_06619_),
    .S1(_06624_),
    .X(_06634_));
 sky130_fd_sc_hd__inv_2 _22040_ (.A(_00003_),
    .Y(_06635_));
 sky130_fd_sc_hd__buf_1 _22041_ (.A(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__buf_1 _22042_ (.A(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__a21o_2 _22043_ (.A1(_06633_),
    .A2(_06634_),
    .B1(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__mux4_2 _22044_ (.A0(\fetch.bht.bhtTable_tag[0][22] ),
    .A1(\fetch.bht.bhtTable_tag[1][22] ),
    .A2(\fetch.bht.bhtTable_tag[2][22] ),
    .A3(\fetch.bht.bhtTable_tag[3][22] ),
    .S0(_06619_),
    .S1(_06624_),
    .X(_06639_));
 sky130_fd_sc_hd__buf_1 _22045_ (.A(_00003_),
    .X(_06640_));
 sky130_fd_sc_hd__buf_1 _22046_ (.A(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__buf_1 _22047_ (.A(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__buf_1 _22048_ (.A(_06615_),
    .X(_06643_));
 sky130_fd_sc_hd__buf_1 _22049_ (.A(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__buf_1 _22050_ (.A(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__buf_1 _22051_ (.A(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__mux2_2 _22052_ (.A0(\fetch.bht.bhtTable_tag[4][22] ),
    .A1(\fetch.bht.bhtTable_tag[5][22] ),
    .S(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__mux2_2 _22053_ (.A0(\fetch.bht.bhtTable_tag[6][22] ),
    .A1(\fetch.bht.bhtTable_tag[7][22] ),
    .S(_06645_),
    .X(_06648_));
 sky130_fd_sc_hd__buf_1 _22054_ (.A(_00001_),
    .X(_06649_));
 sky130_fd_sc_hd__buf_1 _22055_ (.A(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__buf_1 _22056_ (.A(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__buf_1 _22057_ (.A(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__or2b_2 _22058_ (.A(_06648_),
    .B_N(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__o211a_2 _22059_ (.A1(_06624_),
    .A2(_06647_),
    .B1(_06632_),
    .C1(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__a211o_2 _22060_ (.A1(_06639_),
    .A2(_06629_),
    .B1(_06642_),
    .C1(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__o21ai_2 _22061_ (.A1(_06630_),
    .A2(_06638_),
    .B1(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__mux4_2 _22062_ (.A0(\fetch.bht.bhtTable_tag[0][18] ),
    .A1(\fetch.bht.bhtTable_tag[1][18] ),
    .A2(\fetch.bht.bhtTable_tag[2][18] ),
    .A3(\fetch.bht.bhtTable_tag[3][18] ),
    .S0(_06646_),
    .S1(_06652_),
    .X(_06657_));
 sky130_fd_sc_hd__a21o_2 _22063_ (.A1(_06657_),
    .A2(_06629_),
    .B1(_06642_),
    .X(_06658_));
 sky130_fd_sc_hd__and2b_2 _22064_ (.A_N(_06619_),
    .B(\fetch.bht.bhtTable_tag[6][18] ),
    .X(_06659_));
 sky130_fd_sc_hd__a21bo_2 _22065_ (.A1(_06619_),
    .A2(\fetch.bht.bhtTable_tag[7][18] ),
    .B1_N(_06652_),
    .X(_06660_));
 sky130_fd_sc_hd__buf_1 _22066_ (.A(_06652_),
    .X(_06661_));
 sky130_fd_sc_hd__mux2_2 _22067_ (.A0(\fetch.bht.bhtTable_tag[4][18] ),
    .A1(\fetch.bht.bhtTable_tag[5][18] ),
    .S(_06646_),
    .X(_06662_));
 sky130_fd_sc_hd__o221a_2 _22068_ (.A1(_06659_),
    .A2(_06660_),
    .B1(_06661_),
    .B2(_06662_),
    .C1(_06633_),
    .X(_06663_));
 sky130_fd_sc_hd__mux4_2 _22069_ (.A0(\fetch.bht.bhtTable_tag[8][18] ),
    .A1(\fetch.bht.bhtTable_tag[9][18] ),
    .A2(\fetch.bht.bhtTable_tag[10][18] ),
    .A3(\fetch.bht.bhtTable_tag[11][18] ),
    .S0(_06646_),
    .S1(_06624_),
    .X(_06664_));
 sky130_fd_sc_hd__a21oi_2 _22070_ (.A1(_06664_),
    .A2(_06629_),
    .B1(_06637_),
    .Y(_06665_));
 sky130_fd_sc_hd__mux2_2 _22071_ (.A0(\fetch.bht.bhtTable_tag[12][18] ),
    .A1(\fetch.bht.bhtTable_tag[13][18] ),
    .S(_06619_),
    .X(_06666_));
 sky130_fd_sc_hd__mux2_2 _22072_ (.A0(\fetch.bht.bhtTable_tag[14][18] ),
    .A1(\fetch.bht.bhtTable_tag[15][18] ),
    .S(_06618_),
    .X(_06667_));
 sky130_fd_sc_hd__or2b_2 _22073_ (.A(_06667_),
    .B_N(_06624_),
    .X(_06668_));
 sky130_fd_sc_hd__o211ai_2 _22074_ (.A1(_06661_),
    .A2(_06666_),
    .B1(_06633_),
    .C1(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__a2bb2o_2 _22075_ (.A1_N(_06658_),
    .A2_N(_06663_),
    .B1(_06665_),
    .B2(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__a2bb2o_2 _22076_ (.A1_N(io_fetch_address[28]),
    .A2_N(_06656_),
    .B1(_06670_),
    .B2(io_fetch_address[24]),
    .X(_06671_));
 sky130_fd_sc_hd__buf_1 _22077_ (.A(_00002_),
    .X(_06672_));
 sky130_fd_sc_hd__buf_1 _22078_ (.A(_06672_),
    .X(_06673_));
 sky130_fd_sc_hd__buf_1 _22079_ (.A(_06643_),
    .X(_06674_));
 sky130_fd_sc_hd__buf_1 _22080_ (.A(_06649_),
    .X(_06675_));
 sky130_fd_sc_hd__mux4_2 _22081_ (.A0(\fetch.bht.bhtTable_tag[0][7] ),
    .A1(\fetch.bht.bhtTable_tag[1][7] ),
    .A2(\fetch.bht.bhtTable_tag[2][7] ),
    .A3(\fetch.bht.bhtTable_tag[3][7] ),
    .S0(_06674_),
    .S1(_06675_),
    .X(_06676_));
 sky130_fd_sc_hd__buf_1 _22082_ (.A(_06620_),
    .X(_06677_));
 sky130_fd_sc_hd__buf_1 _22083_ (.A(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__buf_1 _22084_ (.A(_06615_),
    .X(_06679_));
 sky130_fd_sc_hd__buf_1 _22085_ (.A(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__mux2_2 _22086_ (.A0(\fetch.bht.bhtTable_tag[4][7] ),
    .A1(\fetch.bht.bhtTable_tag[5][7] ),
    .S(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__and2b_2 _22087_ (.A_N(_06678_),
    .B(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__mux2_2 _22088_ (.A0(\fetch.bht.bhtTable_tag[6][7] ),
    .A1(\fetch.bht.bhtTable_tag[7][7] ),
    .S(_06644_),
    .X(_06683_));
 sky130_fd_sc_hd__buf_1 _22089_ (.A(_00001_),
    .X(_06684_));
 sky130_fd_sc_hd__buf_1 _22090_ (.A(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__buf_1 _22091_ (.A(_06626_),
    .X(_06686_));
 sky130_fd_sc_hd__buf_1 _22092_ (.A(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__a21o_2 _22093_ (.A1(_06683_),
    .A2(_06685_),
    .B1(_06687_),
    .X(_06688_));
 sky130_fd_sc_hd__o22a_2 _22094_ (.A1(_06673_),
    .A2(_06676_),
    .B1(_06682_),
    .B2(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__buf_1 _22095_ (.A(_06621_),
    .X(_06690_));
 sky130_fd_sc_hd__buf_1 _22096_ (.A(_06679_),
    .X(_06691_));
 sky130_fd_sc_hd__mux2_2 _22097_ (.A0(\fetch.bht.bhtTable_tag[12][7] ),
    .A1(\fetch.bht.bhtTable_tag[13][7] ),
    .S(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__and2b_2 _22098_ (.A_N(_06690_),
    .B(_06692_),
    .X(_06693_));
 sky130_fd_sc_hd__mux2_2 _22099_ (.A0(\fetch.bht.bhtTable_tag[14][7] ),
    .A1(\fetch.bht.bhtTable_tag[15][7] ),
    .S(_06680_),
    .X(_06694_));
 sky130_fd_sc_hd__a21o_2 _22100_ (.A1(_06694_),
    .A2(_06690_),
    .B1(_06627_),
    .X(_06695_));
 sky130_fd_sc_hd__mux4_2 _22101_ (.A0(\fetch.bht.bhtTable_tag[8][7] ),
    .A1(\fetch.bht.bhtTable_tag[9][7] ),
    .A2(\fetch.bht.bhtTable_tag[10][7] ),
    .A3(\fetch.bht.bhtTable_tag[11][7] ),
    .S0(_06674_),
    .S1(_06675_),
    .X(_06696_));
 sky130_fd_sc_hd__o221a_2 _22102_ (.A1(_06693_),
    .A2(_06695_),
    .B1(_06696_),
    .B2(_06673_),
    .C1(_06641_),
    .X(_06697_));
 sky130_fd_sc_hd__a21oi_2 _22103_ (.A1(_06636_),
    .A2(_06689_),
    .B1(_06697_),
    .Y(_06698_));
 sky130_fd_sc_hd__buf_1 _22104_ (.A(_06640_),
    .X(_06699_));
 sky130_fd_sc_hd__buf_1 _22105_ (.A(_06691_),
    .X(_06700_));
 sky130_fd_sc_hd__mux2_2 _22106_ (.A0(\fetch.bht.bhtTable_tag[2][3] ),
    .A1(\fetch.bht.bhtTable_tag[3][3] ),
    .S(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__mux2_2 _22107_ (.A0(\fetch.bht.bhtTable_tag[0][3] ),
    .A1(\fetch.bht.bhtTable_tag[1][3] ),
    .S(_06680_),
    .X(_06702_));
 sky130_fd_sc_hd__and2b_2 _22108_ (.A_N(_06678_),
    .B(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__a211oi_2 _22109_ (.A1(_06701_),
    .A2(_06623_),
    .B1(_06673_),
    .C1(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__mux2_2 _22110_ (.A0(\fetch.bht.bhtTable_tag[6][3] ),
    .A1(\fetch.bht.bhtTable_tag[7][3] ),
    .S(_06700_),
    .X(_06705_));
 sky130_fd_sc_hd__buf_1 _22111_ (.A(_06615_),
    .X(_06706_));
 sky130_fd_sc_hd__buf_1 _22112_ (.A(_06706_),
    .X(_06707_));
 sky130_fd_sc_hd__mux2_2 _22113_ (.A0(\fetch.bht.bhtTable_tag[4][3] ),
    .A1(\fetch.bht.bhtTable_tag[5][3] ),
    .S(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__and2b_2 _22114_ (.A_N(_06685_),
    .B(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__a211oi_2 _22115_ (.A1(_06623_),
    .A2(_06705_),
    .B1(_06628_),
    .C1(_06709_),
    .Y(_06710_));
 sky130_fd_sc_hd__mux4_2 _22116_ (.A0(\fetch.bht.bhtTable_tag[8][3] ),
    .A1(\fetch.bht.bhtTable_tag[9][3] ),
    .A2(\fetch.bht.bhtTable_tag[10][3] ),
    .A3(\fetch.bht.bhtTable_tag[11][3] ),
    .S0(_06617_),
    .S1(_06690_),
    .X(_06711_));
 sky130_fd_sc_hd__mux2_2 _22117_ (.A0(\fetch.bht.bhtTable_tag[12][3] ),
    .A1(\fetch.bht.bhtTable_tag[13][3] ),
    .S(_06644_),
    .X(_06712_));
 sky130_fd_sc_hd__and2b_2 _22118_ (.A_N(_06685_),
    .B(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__mux2_2 _22119_ (.A0(\fetch.bht.bhtTable_tag[14][3] ),
    .A1(\fetch.bht.bhtTable_tag[15][3] ),
    .S(_06674_),
    .X(_06714_));
 sky130_fd_sc_hd__a21o_2 _22120_ (.A1(_06714_),
    .A2(_06651_),
    .B1(_06687_),
    .X(_06715_));
 sky130_fd_sc_hd__o221ai_2 _22121_ (.A1(_06632_),
    .A2(_06711_),
    .B1(_06713_),
    .B2(_06715_),
    .C1(_06699_),
    .Y(_06716_));
 sky130_fd_sc_hd__o31a_2 _22122_ (.A1(_06699_),
    .A2(_06704_),
    .A3(_06710_),
    .B1(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__buf_1 _22123_ (.A(io_fetch_address[9]),
    .X(_06718_));
 sky130_fd_sc_hd__o22ai_2 _22124_ (.A1(io_fetch_address[13]),
    .A2(_06698_),
    .B1(_06717_),
    .B2(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__or2_2 _22125_ (.A(_06671_),
    .B(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__mux2_2 _22126_ (.A0(\fetch.bht.bhtTable_tag[10][4] ),
    .A1(\fetch.bht.bhtTable_tag[11][4] ),
    .S(_06680_),
    .X(_06721_));
 sky130_fd_sc_hd__mux2_2 _22127_ (.A0(\fetch.bht.bhtTable_tag[8][4] ),
    .A1(\fetch.bht.bhtTable_tag[9][4] ),
    .S(_06706_),
    .X(_06722_));
 sky130_fd_sc_hd__and2b_2 _22128_ (.A_N(_06677_),
    .B(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__a211oi_2 _22129_ (.A1(_06721_),
    .A2(_06690_),
    .B1(_06672_),
    .C1(_06723_),
    .Y(_06724_));
 sky130_fd_sc_hd__mux2_2 _22130_ (.A0(\fetch.bht.bhtTable_tag[14][4] ),
    .A1(\fetch.bht.bhtTable_tag[15][4] ),
    .S(_06680_),
    .X(_06725_));
 sky130_fd_sc_hd__mux2_2 _22131_ (.A0(\fetch.bht.bhtTable_tag[12][4] ),
    .A1(\fetch.bht.bhtTable_tag[13][4] ),
    .S(_06706_),
    .X(_06726_));
 sky130_fd_sc_hd__and2b_2 _22132_ (.A_N(_06684_),
    .B(_06726_),
    .X(_06727_));
 sky130_fd_sc_hd__a211oi_2 _22133_ (.A1(_06685_),
    .A2(_06725_),
    .B1(_06627_),
    .C1(_06727_),
    .Y(_06728_));
 sky130_fd_sc_hd__mux2_2 _22134_ (.A0(\fetch.bht.bhtTable_tag[6][4] ),
    .A1(\fetch.bht.bhtTable_tag[7][4] ),
    .S(_06643_),
    .X(_06729_));
 sky130_fd_sc_hd__buf_1 _22135_ (.A(_06649_),
    .X(_06730_));
 sky130_fd_sc_hd__nand2_2 _22136_ (.A(_06729_),
    .B(_06730_),
    .Y(_06731_));
 sky130_fd_sc_hd__mux2_2 _22137_ (.A0(\fetch.bht.bhtTable_tag[4][4] ),
    .A1(\fetch.bht.bhtTable_tag[5][4] ),
    .S(_06679_),
    .X(_06732_));
 sky130_fd_sc_hd__or2b_2 _22138_ (.A(_06649_),
    .B_N(_06732_),
    .X(_06733_));
 sky130_fd_sc_hd__mux2_2 _22139_ (.A0(\fetch.bht.bhtTable_tag[2][4] ),
    .A1(\fetch.bht.bhtTable_tag[3][4] ),
    .S(_06706_),
    .X(_06734_));
 sky130_fd_sc_hd__mux2_2 _22140_ (.A0(\fetch.bht.bhtTable_tag[0][4] ),
    .A1(\fetch.bht.bhtTable_tag[1][4] ),
    .S(_06615_),
    .X(_06735_));
 sky130_fd_sc_hd__and2b_2 _22141_ (.A_N(_06620_),
    .B(_06735_),
    .X(_06736_));
 sky130_fd_sc_hd__a211oi_2 _22142_ (.A1(_06734_),
    .A2(_06677_),
    .B1(_00002_),
    .C1(_06736_),
    .Y(_06737_));
 sky130_fd_sc_hd__a311o_2 _22143_ (.A1(_06672_),
    .A2(_06731_),
    .A3(_06733_),
    .B1(_06737_),
    .C1(_06640_),
    .X(_06738_));
 sky130_fd_sc_hd__o31a_2 _22144_ (.A1(_06635_),
    .A2(_06724_),
    .A3(_06728_),
    .B1(_06738_),
    .X(_06739_));
 sky130_fd_sc_hd__buf_1 _22145_ (.A(_06642_),
    .X(_06740_));
 sky130_fd_sc_hd__mux4_2 _22146_ (.A0(\fetch.bht.bhtTable_tag[0][23] ),
    .A1(\fetch.bht.bhtTable_tag[1][23] ),
    .A2(\fetch.bht.bhtTable_tag[2][23] ),
    .A3(\fetch.bht.bhtTable_tag[3][23] ),
    .S0(_06618_),
    .S1(_06652_),
    .X(_06741_));
 sky130_fd_sc_hd__nor2_2 _22147_ (.A(_06632_),
    .B(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__mux2_2 _22148_ (.A0(\fetch.bht.bhtTable_tag[6][23] ),
    .A1(\fetch.bht.bhtTable_tag[7][23] ),
    .S(_06646_),
    .X(_06743_));
 sky130_fd_sc_hd__mux2_2 _22149_ (.A0(\fetch.bht.bhtTable_tag[4][23] ),
    .A1(\fetch.bht.bhtTable_tag[5][23] ),
    .S(_06618_),
    .X(_06744_));
 sky130_fd_sc_hd__and2b_2 _22150_ (.A_N(_06652_),
    .B(_06744_),
    .X(_06745_));
 sky130_fd_sc_hd__a211oi_2 _22151_ (.A1(_06661_),
    .A2(_06743_),
    .B1(_06629_),
    .C1(_06745_),
    .Y(_06746_));
 sky130_fd_sc_hd__mux4_2 _22152_ (.A0(\fetch.bht.bhtTable_tag[8][23] ),
    .A1(\fetch.bht.bhtTable_tag[9][23] ),
    .A2(\fetch.bht.bhtTable_tag[10][23] ),
    .A3(\fetch.bht.bhtTable_tag[11][23] ),
    .S0(_06618_),
    .S1(_06623_),
    .X(_06747_));
 sky130_fd_sc_hd__mux2_2 _22153_ (.A0(\fetch.bht.bhtTable_tag[12][23] ),
    .A1(\fetch.bht.bhtTable_tag[13][23] ),
    .S(_06618_),
    .X(_06748_));
 sky130_fd_sc_hd__and2b_2 _22154_ (.A_N(_06652_),
    .B(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__mux2_2 _22155_ (.A0(\fetch.bht.bhtTable_tag[14][23] ),
    .A1(\fetch.bht.bhtTable_tag[15][23] ),
    .S(_06618_),
    .X(_06750_));
 sky130_fd_sc_hd__a21o_2 _22156_ (.A1(_06750_),
    .A2(_06652_),
    .B1(_06629_),
    .X(_06751_));
 sky130_fd_sc_hd__o221ai_2 _22157_ (.A1(_06632_),
    .A2(_06747_),
    .B1(_06749_),
    .B2(_06751_),
    .C1(_06642_),
    .Y(_06752_));
 sky130_fd_sc_hd__o31a_2 _22158_ (.A1(_06740_),
    .A2(_06742_),
    .A3(_06746_),
    .B1(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__buf_1 _22159_ (.A(_06616_),
    .X(_06754_));
 sky130_fd_sc_hd__mux4_2 _22160_ (.A0(\fetch.bht.bhtTable_tag[0][13] ),
    .A1(\fetch.bht.bhtTable_tag[1][13] ),
    .A2(\fetch.bht.bhtTable_tag[2][13] ),
    .A3(\fetch.bht.bhtTable_tag[3][13] ),
    .S0(_06754_),
    .S1(_06622_),
    .X(_06755_));
 sky130_fd_sc_hd__mux2_2 _22161_ (.A0(\fetch.bht.bhtTable_tag[4][13] ),
    .A1(\fetch.bht.bhtTable_tag[5][13] ),
    .S(_06707_),
    .X(_06756_));
 sky130_fd_sc_hd__and2b_2 _22162_ (.A_N(_06678_),
    .B(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__mux2_2 _22163_ (.A0(\fetch.bht.bhtTable_tag[6][13] ),
    .A1(\fetch.bht.bhtTable_tag[7][13] ),
    .S(_06644_),
    .X(_06758_));
 sky130_fd_sc_hd__a21o_2 _22164_ (.A1(_06758_),
    .A2(_06685_),
    .B1(_06687_),
    .X(_06759_));
 sky130_fd_sc_hd__o22a_2 _22165_ (.A1(_06673_),
    .A2(_06755_),
    .B1(_06757_),
    .B2(_06759_),
    .X(_06760_));
 sky130_fd_sc_hd__mux2_2 _22166_ (.A0(\fetch.bht.bhtTable_tag[12][13] ),
    .A1(\fetch.bht.bhtTable_tag[13][13] ),
    .S(_06680_),
    .X(_06761_));
 sky130_fd_sc_hd__and2b_2 _22167_ (.A_N(_06690_),
    .B(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__mux2_2 _22168_ (.A0(\fetch.bht.bhtTable_tag[14][13] ),
    .A1(\fetch.bht.bhtTable_tag[15][13] ),
    .S(_06644_),
    .X(_06763_));
 sky130_fd_sc_hd__a21o_2 _22169_ (.A1(_06763_),
    .A2(_06678_),
    .B1(_06627_),
    .X(_06764_));
 sky130_fd_sc_hd__mux4_2 _22170_ (.A0(\fetch.bht.bhtTable_tag[8][13] ),
    .A1(\fetch.bht.bhtTable_tag[9][13] ),
    .A2(\fetch.bht.bhtTable_tag[10][13] ),
    .A3(\fetch.bht.bhtTable_tag[11][13] ),
    .S0(_06754_),
    .S1(_06622_),
    .X(_06765_));
 sky130_fd_sc_hd__o221a_2 _22171_ (.A1(_06762_),
    .A2(_06764_),
    .B1(_06765_),
    .B2(_06673_),
    .C1(_06699_),
    .X(_06766_));
 sky130_fd_sc_hd__a21oi_2 _22172_ (.A1(_06636_),
    .A2(_06760_),
    .B1(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__o22a_2 _22173_ (.A1(io_fetch_address[29]),
    .A2(_06753_),
    .B1(_06767_),
    .B2(io_fetch_address[19]),
    .X(_06768_));
 sky130_fd_sc_hd__o221ai_2 _22174_ (.A1(io_fetch_address[10]),
    .A2(_06739_),
    .B1(_06670_),
    .B2(io_fetch_address[24]),
    .C1(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__mux2_2 _22175_ (.A0(\fetch.bht.bhtTable_tag[6][25] ),
    .A1(\fetch.bht.bhtTable_tag[7][25] ),
    .S(_06619_),
    .X(_06770_));
 sky130_fd_sc_hd__mux2_2 _22176_ (.A0(\fetch.bht.bhtTable_tag[4][25] ),
    .A1(\fetch.bht.bhtTable_tag[5][25] ),
    .S(_06646_),
    .X(_06771_));
 sky130_fd_sc_hd__and2b_2 _22177_ (.A_N(_06624_),
    .B(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__a211oi_2 _22178_ (.A1(_06661_),
    .A2(_06770_),
    .B1(_06629_),
    .C1(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__mux2_2 _22179_ (.A0(\fetch.bht.bhtTable_tag[2][25] ),
    .A1(\fetch.bht.bhtTable_tag[3][25] ),
    .S(_06619_),
    .X(_06774_));
 sky130_fd_sc_hd__mux2_2 _22180_ (.A0(\fetch.bht.bhtTable_tag[0][25] ),
    .A1(\fetch.bht.bhtTable_tag[1][25] ),
    .S(_06646_),
    .X(_06775_));
 sky130_fd_sc_hd__and2b_2 _22181_ (.A_N(_06624_),
    .B(_06775_),
    .X(_06776_));
 sky130_fd_sc_hd__a211oi_2 _22182_ (.A1(_06774_),
    .A2(_06661_),
    .B1(_06633_),
    .C1(_06776_),
    .Y(_06777_));
 sky130_fd_sc_hd__mux4_2 _22183_ (.A0(\fetch.bht.bhtTable_tag[8][25] ),
    .A1(\fetch.bht.bhtTable_tag[9][25] ),
    .A2(\fetch.bht.bhtTable_tag[10][25] ),
    .A3(\fetch.bht.bhtTable_tag[11][25] ),
    .S0(_06619_),
    .S1(_06624_),
    .X(_06778_));
 sky130_fd_sc_hd__mux2_2 _22184_ (.A0(\fetch.bht.bhtTable_tag[12][25] ),
    .A1(\fetch.bht.bhtTable_tag[13][25] ),
    .S(_06646_),
    .X(_06779_));
 sky130_fd_sc_hd__and2b_2 _22185_ (.A_N(_06624_),
    .B(_06779_),
    .X(_06780_));
 sky130_fd_sc_hd__mux2_2 _22186_ (.A0(\fetch.bht.bhtTable_tag[14][25] ),
    .A1(\fetch.bht.bhtTable_tag[15][25] ),
    .S(_06646_),
    .X(_06781_));
 sky130_fd_sc_hd__a21o_2 _22187_ (.A1(_06781_),
    .A2(_06661_),
    .B1(_06629_),
    .X(_06782_));
 sky130_fd_sc_hd__o221ai_2 _22188_ (.A1(_06633_),
    .A2(_06778_),
    .B1(_06780_),
    .B2(_06782_),
    .C1(_06642_),
    .Y(_06783_));
 sky130_fd_sc_hd__o31a_2 _22189_ (.A1(_06740_),
    .A2(_06773_),
    .A3(_06777_),
    .B1(_06783_),
    .X(_06784_));
 sky130_fd_sc_hd__xnor2_2 _22190_ (.A(io_fetch_address[31]),
    .B(_06784_),
    .Y(_06785_));
 sky130_fd_sc_hd__mux4_2 _22191_ (.A0(\fetch.bht.bhtTable_tag[0][5] ),
    .A1(\fetch.bht.bhtTable_tag[1][5] ),
    .A2(\fetch.bht.bhtTable_tag[2][5] ),
    .A3(\fetch.bht.bhtTable_tag[3][5] ),
    .S0(_06700_),
    .S1(_06685_),
    .X(_06786_));
 sky130_fd_sc_hd__mux4_2 _22192_ (.A0(\fetch.bht.bhtTable_tag[4][5] ),
    .A1(\fetch.bht.bhtTable_tag[5][5] ),
    .A2(\fetch.bht.bhtTable_tag[6][5] ),
    .A3(\fetch.bht.bhtTable_tag[7][5] ),
    .S0(_06700_),
    .S1(_06685_),
    .X(_06787_));
 sky130_fd_sc_hd__mux2_2 _22193_ (.A0(_06786_),
    .A1(_06787_),
    .S(_06632_),
    .X(_06788_));
 sky130_fd_sc_hd__mux4_2 _22194_ (.A0(\fetch.bht.bhtTable_tag[12][5] ),
    .A1(\fetch.bht.bhtTable_tag[13][5] ),
    .A2(\fetch.bht.bhtTable_tag[14][5] ),
    .A3(\fetch.bht.bhtTable_tag[15][5] ),
    .S0(_06700_),
    .S1(_06651_),
    .X(_06789_));
 sky130_fd_sc_hd__buf_1 _22195_ (.A(_00002_),
    .X(_06790_));
 sky130_fd_sc_hd__mux4_2 _22196_ (.A0(\fetch.bht.bhtTable_tag[8][5] ),
    .A1(\fetch.bht.bhtTable_tag[9][5] ),
    .A2(\fetch.bht.bhtTable_tag[10][5] ),
    .A3(\fetch.bht.bhtTable_tag[11][5] ),
    .S0(_06644_),
    .S1(_06730_),
    .X(_06791_));
 sky130_fd_sc_hd__or2_2 _22197_ (.A(_06790_),
    .B(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__o211a_2 _22198_ (.A1(_06628_),
    .A2(_06789_),
    .B1(_06699_),
    .C1(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__a21oi_2 _22199_ (.A1(_06637_),
    .A2(_06788_),
    .B1(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__buf_1 _22200_ (.A(io_fetch_address[28]),
    .X(_06795_));
 sky130_fd_sc_hd__mux4_2 _22201_ (.A0(\fetch.bht.bhtTable_tag[0][24] ),
    .A1(\fetch.bht.bhtTable_tag[1][24] ),
    .A2(\fetch.bht.bhtTable_tag[2][24] ),
    .A3(\fetch.bht.bhtTable_tag[3][24] ),
    .S0(_06646_),
    .S1(_06652_),
    .X(_06796_));
 sky130_fd_sc_hd__mux2_2 _22202_ (.A0(\fetch.bht.bhtTable_tag[4][24] ),
    .A1(\fetch.bht.bhtTable_tag[5][24] ),
    .S(_06618_),
    .X(_06797_));
 sky130_fd_sc_hd__mux2_2 _22203_ (.A0(\fetch.bht.bhtTable_tag[6][24] ),
    .A1(\fetch.bht.bhtTable_tag[7][24] ),
    .S(_06700_),
    .X(_06798_));
 sky130_fd_sc_hd__or2b_2 _22204_ (.A(_06798_),
    .B_N(_06623_),
    .X(_06799_));
 sky130_fd_sc_hd__o211a_2 _22205_ (.A1(_06652_),
    .A2(_06797_),
    .B1(_06632_),
    .C1(_06799_),
    .X(_06800_));
 sky130_fd_sc_hd__a21oi_2 _22206_ (.A1(_06629_),
    .A2(_06796_),
    .B1(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__mux4_2 _22207_ (.A0(\fetch.bht.bhtTable_tag[12][24] ),
    .A1(\fetch.bht.bhtTable_tag[13][24] ),
    .A2(\fetch.bht.bhtTable_tag[14][24] ),
    .A3(\fetch.bht.bhtTable_tag[15][24] ),
    .S0(_06645_),
    .S1(_06651_),
    .X(_06802_));
 sky130_fd_sc_hd__mux4_2 _22208_ (.A0(\fetch.bht.bhtTable_tag[8][24] ),
    .A1(\fetch.bht.bhtTable_tag[9][24] ),
    .A2(\fetch.bht.bhtTable_tag[10][24] ),
    .A3(\fetch.bht.bhtTable_tag[11][24] ),
    .S0(_06645_),
    .S1(_06651_),
    .X(_06803_));
 sky130_fd_sc_hd__mux2_2 _22209_ (.A0(_06802_),
    .A1(_06803_),
    .S(_06628_),
    .X(_06804_));
 sky130_fd_sc_hd__nand2_2 _22210_ (.A(_06804_),
    .B(_06642_),
    .Y(_06805_));
 sky130_fd_sc_hd__o21a_2 _22211_ (.A1(_06642_),
    .A2(_06801_),
    .B1(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__xnor2_2 _22212_ (.A(io_fetch_address[30]),
    .B(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__a221oi_2 _22213_ (.A1(io_fetch_address[11]),
    .A2(_06794_),
    .B1(_06656_),
    .B2(_06795_),
    .C1(_06807_),
    .Y(_06808_));
 sky130_fd_sc_hd__buf_1 _22214_ (.A(_06615_),
    .X(_06809_));
 sky130_fd_sc_hd__mux4_2 _22215_ (.A0(\fetch.bht.bhtTable_tag[12][20] ),
    .A1(\fetch.bht.bhtTable_tag[13][20] ),
    .A2(\fetch.bht.bhtTable_tag[14][20] ),
    .A3(\fetch.bht.bhtTable_tag[15][20] ),
    .S0(_06809_),
    .S1(_06649_),
    .X(_06810_));
 sky130_fd_sc_hd__nand2_2 _22216_ (.A(_06631_),
    .B(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__a21bo_2 _22217_ (.A1(_06707_),
    .A2(\fetch.bht.bhtTable_tag[11][20] ),
    .B1_N(_06649_),
    .X(_06812_));
 sky130_fd_sc_hd__and2b_2 _22218_ (.A_N(_06691_),
    .B(\fetch.bht.bhtTable_tag[10][20] ),
    .X(_06813_));
 sky130_fd_sc_hd__mux2_2 _22219_ (.A0(\fetch.bht.bhtTable_tag[8][20] ),
    .A1(\fetch.bht.bhtTable_tag[9][20] ),
    .S(_06616_),
    .X(_06814_));
 sky130_fd_sc_hd__o221ai_2 _22220_ (.A1(_06812_),
    .A2(_06813_),
    .B1(_06675_),
    .B2(_06814_),
    .C1(_06627_),
    .Y(_06815_));
 sky130_fd_sc_hd__mux4_2 _22221_ (.A0(\fetch.bht.bhtTable_tag[4][20] ),
    .A1(\fetch.bht.bhtTable_tag[5][20] ),
    .A2(\fetch.bht.bhtTable_tag[6][20] ),
    .A3(\fetch.bht.bhtTable_tag[7][20] ),
    .S0(_06809_),
    .S1(_06649_),
    .X(_06816_));
 sky130_fd_sc_hd__mux4_2 _22222_ (.A0(\fetch.bht.bhtTable_tag[0][20] ),
    .A1(\fetch.bht.bhtTable_tag[1][20] ),
    .A2(\fetch.bht.bhtTable_tag[2][20] ),
    .A3(\fetch.bht.bhtTable_tag[3][20] ),
    .S0(_06615_),
    .S1(_06620_),
    .X(_06817_));
 sky130_fd_sc_hd__a21o_2 _22223_ (.A1(_06817_),
    .A2(_06686_),
    .B1(_00003_),
    .X(_06818_));
 sky130_fd_sc_hd__a21oi_2 _22224_ (.A1(_06672_),
    .A2(_06816_),
    .B1(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__a311o_2 _22225_ (.A1(_06740_),
    .A2(_06811_),
    .A3(_06815_),
    .B1(_06819_),
    .C1(io_fetch_address[26]),
    .X(_06820_));
 sky130_fd_sc_hd__nand2_2 _22226_ (.A(_06718_),
    .B(_06717_),
    .Y(_06821_));
 sky130_fd_sc_hd__nand4b_2 _22227_ (.A_N(_06785_),
    .B(_06808_),
    .C(_06820_),
    .D(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__mux4_2 _22228_ (.A0(\fetch.bht.bhtTable_tag[0][15] ),
    .A1(\fetch.bht.bhtTable_tag[1][15] ),
    .A2(\fetch.bht.bhtTable_tag[2][15] ),
    .A3(\fetch.bht.bhtTable_tag[3][15] ),
    .S0(_06617_),
    .S1(_06622_),
    .X(_06823_));
 sky130_fd_sc_hd__nand2_2 _22229_ (.A(_06823_),
    .B(_06628_),
    .Y(_06824_));
 sky130_fd_sc_hd__mux4_2 _22230_ (.A0(\fetch.bht.bhtTable_tag[4][15] ),
    .A1(\fetch.bht.bhtTable_tag[5][15] ),
    .A2(\fetch.bht.bhtTable_tag[6][15] ),
    .A3(\fetch.bht.bhtTable_tag[7][15] ),
    .S0(_06754_),
    .S1(_06622_),
    .X(_06825_));
 sky130_fd_sc_hd__nand2_2 _22231_ (.A(_06632_),
    .B(_06825_),
    .Y(_06826_));
 sky130_fd_sc_hd__mux2_2 _22232_ (.A0(\fetch.bht.bhtTable_tag[12][15] ),
    .A1(\fetch.bht.bhtTable_tag[13][15] ),
    .S(_06700_),
    .X(_06827_));
 sky130_fd_sc_hd__mux2_2 _22233_ (.A0(\fetch.bht.bhtTable_tag[14][15] ),
    .A1(\fetch.bht.bhtTable_tag[15][15] ),
    .S(_06680_),
    .X(_06828_));
 sky130_fd_sc_hd__or2b_2 _22234_ (.A(_06828_),
    .B_N(_06678_),
    .X(_06829_));
 sky130_fd_sc_hd__o211ai_2 _22235_ (.A1(_06623_),
    .A2(_06827_),
    .B1(_06673_),
    .C1(_06829_),
    .Y(_06830_));
 sky130_fd_sc_hd__mux4_2 _22236_ (.A0(\fetch.bht.bhtTable_tag[8][15] ),
    .A1(\fetch.bht.bhtTable_tag[9][15] ),
    .A2(\fetch.bht.bhtTable_tag[10][15] ),
    .A3(\fetch.bht.bhtTable_tag[11][15] ),
    .S0(_06754_),
    .S1(_06675_),
    .X(_06831_));
 sky130_fd_sc_hd__a21oi_2 _22237_ (.A1(_06831_),
    .A2(_06628_),
    .B1(_06635_),
    .Y(_06832_));
 sky130_fd_sc_hd__a32o_2 _22238_ (.A1(_06636_),
    .A2(_06824_),
    .A3(_06826_),
    .B1(_06830_),
    .B2(_06832_),
    .X(_06833_));
 sky130_fd_sc_hd__nor2_2 _22239_ (.A(io_fetch_address[21]),
    .B(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__mux2_2 _22240_ (.A0(\fetch.bht.bhtTable_tag[2][19] ),
    .A1(\fetch.bht.bhtTable_tag[3][19] ),
    .S(_06707_),
    .X(_06835_));
 sky130_fd_sc_hd__mux2_2 _22241_ (.A0(\fetch.bht.bhtTable_tag[0][19] ),
    .A1(\fetch.bht.bhtTable_tag[1][19] ),
    .S(_06706_),
    .X(_06836_));
 sky130_fd_sc_hd__and2b_2 _22242_ (.A_N(_06684_),
    .B(_06836_),
    .X(_06837_));
 sky130_fd_sc_hd__a211oi_2 _22243_ (.A1(_06835_),
    .A2(_06678_),
    .B1(_06672_),
    .C1(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__mux2_2 _22244_ (.A0(\fetch.bht.bhtTable_tag[6][19] ),
    .A1(\fetch.bht.bhtTable_tag[7][19] ),
    .S(_06707_),
    .X(_06839_));
 sky130_fd_sc_hd__mux2_2 _22245_ (.A0(\fetch.bht.bhtTable_tag[4][19] ),
    .A1(\fetch.bht.bhtTable_tag[5][19] ),
    .S(_06706_),
    .X(_06840_));
 sky130_fd_sc_hd__and2b_2 _22246_ (.A_N(_06684_),
    .B(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__a211oi_2 _22247_ (.A1(_06685_),
    .A2(_06839_),
    .B1(_06687_),
    .C1(_06841_),
    .Y(_06842_));
 sky130_fd_sc_hd__mux4_2 _22248_ (.A0(\fetch.bht.bhtTable_tag[8][19] ),
    .A1(\fetch.bht.bhtTable_tag[9][19] ),
    .A2(\fetch.bht.bhtTable_tag[10][19] ),
    .A3(\fetch.bht.bhtTable_tag[11][19] ),
    .S0(_06616_),
    .S1(_06621_),
    .X(_06843_));
 sky130_fd_sc_hd__mux2_2 _22249_ (.A0(\fetch.bht.bhtTable_tag[12][19] ),
    .A1(\fetch.bht.bhtTable_tag[13][19] ),
    .S(_06643_),
    .X(_06844_));
 sky130_fd_sc_hd__and2b_2 _22250_ (.A_N(_06684_),
    .B(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__mux2_2 _22251_ (.A0(\fetch.bht.bhtTable_tag[14][19] ),
    .A1(\fetch.bht.bhtTable_tag[15][19] ),
    .S(_06809_),
    .X(_06846_));
 sky130_fd_sc_hd__a21o_2 _22252_ (.A1(_06846_),
    .A2(_06730_),
    .B1(_06686_),
    .X(_06847_));
 sky130_fd_sc_hd__o221ai_2 _22253_ (.A1(_06631_),
    .A2(_06843_),
    .B1(_06845_),
    .B2(_06847_),
    .C1(_06640_),
    .Y(_06848_));
 sky130_fd_sc_hd__o311a_2 _22254_ (.A1(_06642_),
    .A2(_06838_),
    .A3(_06842_),
    .B1(_06848_),
    .C1(io_fetch_address[25]),
    .X(_06849_));
 sky130_fd_sc_hd__mux4_2 _22255_ (.A0(\fetch.bht.bhtTable_tag[0][17] ),
    .A1(\fetch.bht.bhtTable_tag[1][17] ),
    .A2(\fetch.bht.bhtTable_tag[2][17] ),
    .A3(\fetch.bht.bhtTable_tag[3][17] ),
    .S0(_06691_),
    .S1(_06677_),
    .X(_06850_));
 sky130_fd_sc_hd__mux2_2 _22256_ (.A0(\fetch.bht.bhtTable_tag[4][17] ),
    .A1(\fetch.bht.bhtTable_tag[5][17] ),
    .S(_06643_),
    .X(_06851_));
 sky130_fd_sc_hd__and2b_2 _22257_ (.A_N(_06650_),
    .B(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__mux2_2 _22258_ (.A0(\fetch.bht.bhtTable_tag[6][17] ),
    .A1(\fetch.bht.bhtTable_tag[7][17] ),
    .S(_06616_),
    .X(_06853_));
 sky130_fd_sc_hd__a21o_2 _22259_ (.A1(_06853_),
    .A2(_06650_),
    .B1(_06686_),
    .X(_06854_));
 sky130_fd_sc_hd__o22a_2 _22260_ (.A1(_06790_),
    .A2(_06850_),
    .B1(_06852_),
    .B2(_06854_),
    .X(_06855_));
 sky130_fd_sc_hd__mux2_2 _22261_ (.A0(\fetch.bht.bhtTable_tag[12][17] ),
    .A1(\fetch.bht.bhtTable_tag[13][17] ),
    .S(_06643_),
    .X(_06856_));
 sky130_fd_sc_hd__and2b_2 _22262_ (.A_N(_06730_),
    .B(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__mux2_2 _22263_ (.A0(\fetch.bht.bhtTable_tag[14][17] ),
    .A1(\fetch.bht.bhtTable_tag[15][17] ),
    .S(_06809_),
    .X(_06858_));
 sky130_fd_sc_hd__a21o_2 _22264_ (.A1(_06858_),
    .A2(_06650_),
    .B1(_06686_),
    .X(_06859_));
 sky130_fd_sc_hd__mux4_2 _22265_ (.A0(\fetch.bht.bhtTable_tag[8][17] ),
    .A1(\fetch.bht.bhtTable_tag[9][17] ),
    .A2(\fetch.bht.bhtTable_tag[10][17] ),
    .A3(\fetch.bht.bhtTable_tag[11][17] ),
    .S0(_06691_),
    .S1(_06677_),
    .X(_06860_));
 sky130_fd_sc_hd__o221a_2 _22266_ (.A1(_06857_),
    .A2(_06859_),
    .B1(_06860_),
    .B2(_06790_),
    .C1(_06641_),
    .X(_06861_));
 sky130_fd_sc_hd__a21oi_2 _22267_ (.A1(_06636_),
    .A2(_06855_),
    .B1(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__xnor2_2 _22268_ (.A(io_fetch_address[23]),
    .B(_06862_),
    .Y(_06863_));
 sky130_fd_sc_hd__or3_2 _22269_ (.A(_06834_),
    .B(_06849_),
    .C(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__mux2_2 _22270_ (.A0(\fetch.bht.bhtTable_tag[12][6] ),
    .A1(\fetch.bht.bhtTable_tag[13][6] ),
    .S(_06617_),
    .X(_06865_));
 sky130_fd_sc_hd__and2b_2 _22271_ (.A_N(_06651_),
    .B(_06865_),
    .X(_06866_));
 sky130_fd_sc_hd__mux2_2 _22272_ (.A0(\fetch.bht.bhtTable_tag[14][6] ),
    .A1(\fetch.bht.bhtTable_tag[15][6] ),
    .S(_06700_),
    .X(_06867_));
 sky130_fd_sc_hd__a21o_2 _22273_ (.A1(_06867_),
    .A2(_06623_),
    .B1(_06687_),
    .X(_06868_));
 sky130_fd_sc_hd__mux4_2 _22274_ (.A0(\fetch.bht.bhtTable_tag[8][6] ),
    .A1(\fetch.bht.bhtTable_tag[9][6] ),
    .A2(\fetch.bht.bhtTable_tag[10][6] ),
    .A3(\fetch.bht.bhtTable_tag[11][6] ),
    .S0(_06645_),
    .S1(_06651_),
    .X(_06869_));
 sky130_fd_sc_hd__o22a_2 _22275_ (.A1(_06866_),
    .A2(_06868_),
    .B1(_06869_),
    .B2(_06632_),
    .X(_06870_));
 sky130_fd_sc_hd__mux4_2 _22276_ (.A0(\fetch.bht.bhtTable_tag[0][6] ),
    .A1(\fetch.bht.bhtTable_tag[1][6] ),
    .A2(\fetch.bht.bhtTable_tag[2][6] ),
    .A3(\fetch.bht.bhtTable_tag[3][6] ),
    .S0(_06645_),
    .S1(_06651_),
    .X(_06871_));
 sky130_fd_sc_hd__mux2_2 _22277_ (.A0(\fetch.bht.bhtTable_tag[4][6] ),
    .A1(\fetch.bht.bhtTable_tag[5][6] ),
    .S(_06617_),
    .X(_06872_));
 sky130_fd_sc_hd__and2b_2 _22278_ (.A_N(_06651_),
    .B(_06872_),
    .X(_06873_));
 sky130_fd_sc_hd__mux2_2 _22279_ (.A0(\fetch.bht.bhtTable_tag[6][6] ),
    .A1(\fetch.bht.bhtTable_tag[7][6] ),
    .S(_06700_),
    .X(_06874_));
 sky130_fd_sc_hd__a21o_2 _22280_ (.A1(_06874_),
    .A2(_06623_),
    .B1(_06628_),
    .X(_06875_));
 sky130_fd_sc_hd__o221a_2 _22281_ (.A1(_06632_),
    .A2(_06871_),
    .B1(_06873_),
    .B2(_06875_),
    .C1(_06636_),
    .X(_06876_));
 sky130_fd_sc_hd__a21oi_2 _22282_ (.A1(_06642_),
    .A2(_06870_),
    .B1(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__buf_1 _22283_ (.A(_06679_),
    .X(_06878_));
 sky130_fd_sc_hd__mux4_2 _22284_ (.A0(\fetch.bht.bhtTable_tag[4][11] ),
    .A1(\fetch.bht.bhtTable_tag[5][11] ),
    .A2(\fetch.bht.bhtTable_tag[6][11] ),
    .A3(\fetch.bht.bhtTable_tag[7][11] ),
    .S0(_06878_),
    .S1(_06677_),
    .X(_06879_));
 sky130_fd_sc_hd__mux4_2 _22285_ (.A0(\fetch.bht.bhtTable_tag[0][11] ),
    .A1(\fetch.bht.bhtTable_tag[1][11] ),
    .A2(\fetch.bht.bhtTable_tag[2][11] ),
    .A3(\fetch.bht.bhtTable_tag[3][11] ),
    .S0(_06878_),
    .S1(_06621_),
    .X(_06880_));
 sky130_fd_sc_hd__mux2_2 _22286_ (.A0(_06879_),
    .A1(_06880_),
    .S(_06627_),
    .X(_06881_));
 sky130_fd_sc_hd__mux4_2 _22287_ (.A0(\fetch.bht.bhtTable_tag[8][11] ),
    .A1(\fetch.bht.bhtTable_tag[9][11] ),
    .A2(\fetch.bht.bhtTable_tag[10][11] ),
    .A3(\fetch.bht.bhtTable_tag[11][11] ),
    .S0(_06754_),
    .S1(_06675_),
    .X(_06882_));
 sky130_fd_sc_hd__nor2_2 _22288_ (.A(_06673_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__mux4_2 _22289_ (.A0(\fetch.bht.bhtTable_tag[12][11] ),
    .A1(\fetch.bht.bhtTable_tag[13][11] ),
    .A2(\fetch.bht.bhtTable_tag[14][11] ),
    .A3(\fetch.bht.bhtTable_tag[15][11] ),
    .S0(_06674_),
    .S1(_06650_),
    .X(_06884_));
 sky130_fd_sc_hd__o21ai_2 _22290_ (.A1(_06687_),
    .A2(_06884_),
    .B1(_06641_),
    .Y(_06885_));
 sky130_fd_sc_hd__o2bb2a_2 _22291_ (.A1_N(_06636_),
    .A2_N(_06881_),
    .B1(_06883_),
    .B2(_06885_),
    .X(_06886_));
 sky130_fd_sc_hd__buf_1 _22292_ (.A(io_fetch_address[17]),
    .X(_06887_));
 sky130_fd_sc_hd__a22o_2 _22293_ (.A1(io_fetch_address[12]),
    .A2(_06877_),
    .B1(_06886_),
    .B2(_06887_),
    .X(_06888_));
 sky130_fd_sc_hd__or2_2 _22294_ (.A(io_fetch_address[11]),
    .B(_06794_),
    .X(_06889_));
 sky130_fd_sc_hd__or2_2 _22295_ (.A(_06887_),
    .B(_06886_),
    .X(_06890_));
 sky130_fd_sc_hd__or4bb_2 _22296_ (.A(_06864_),
    .B(_06888_),
    .C_N(_06889_),
    .D_N(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__o31a_2 _22297_ (.A1(_06641_),
    .A2(_06838_),
    .A3(_06842_),
    .B1(_06848_),
    .X(_06892_));
 sky130_fd_sc_hd__a2bb2o_2 _22298_ (.A1_N(io_fetch_address[25]),
    .A2_N(_06892_),
    .B1(_06739_),
    .B2(io_fetch_address[10]),
    .X(_06893_));
 sky130_fd_sc_hd__o311a_2 _22299_ (.A1(_06642_),
    .A2(_06742_),
    .A3(_06746_),
    .B1(_06752_),
    .C1(io_fetch_address[29]),
    .X(_06894_));
 sky130_fd_sc_hd__a22o_2 _22300_ (.A1(io_fetch_address[21]),
    .A2(_06833_),
    .B1(_06698_),
    .B2(io_fetch_address[13]),
    .X(_06895_));
 sky130_fd_sc_hd__or2_2 _22301_ (.A(io_fetch_address[12]),
    .B(_06877_),
    .X(_06896_));
 sky130_fd_sc_hd__nand2_2 _22302_ (.A(io_fetch_address[19]),
    .B(_06767_),
    .Y(_06897_));
 sky130_fd_sc_hd__or4bb_2 _22303_ (.A(_06894_),
    .B(_06895_),
    .C_N(_06896_),
    .D_N(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__mux2_2 _22304_ (.A0(\fetch.bht.bhtTable_tag[4][0] ),
    .A1(\fetch.bht.bhtTable_tag[5][0] ),
    .S(_06878_),
    .X(_06899_));
 sky130_fd_sc_hd__and2b_2 _22305_ (.A_N(_06690_),
    .B(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__or2b_2 _22306_ (.A(\fetch.bht.bhtTable_tag[7][0] ),
    .B_N(_06674_),
    .X(_06901_));
 sky130_fd_sc_hd__o211a_2 _22307_ (.A1(_06645_),
    .A2(\fetch.bht.bhtTable_tag[6][0] ),
    .B1(_06690_),
    .C1(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__mux2_2 _22308_ (.A0(\fetch.bht.bhtTable_tag[2][0] ),
    .A1(\fetch.bht.bhtTable_tag[3][0] ),
    .S(_06644_),
    .X(_06903_));
 sky130_fd_sc_hd__mux2_2 _22309_ (.A0(\fetch.bht.bhtTable_tag[0][0] ),
    .A1(\fetch.bht.bhtTable_tag[1][0] ),
    .S(_06706_),
    .X(_06904_));
 sky130_fd_sc_hd__and2b_2 _22310_ (.A_N(_06684_),
    .B(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__a211o_2 _22311_ (.A1(_06903_),
    .A2(_06678_),
    .B1(_06631_),
    .C1(_06905_),
    .X(_06906_));
 sky130_fd_sc_hd__o311a_2 _22312_ (.A1(_06628_),
    .A2(_06900_),
    .A3(_06902_),
    .B1(_06906_),
    .C1(_06636_),
    .X(_06907_));
 sky130_fd_sc_hd__mux4_2 _22313_ (.A0(\fetch.bht.bhtTable_tag[12][0] ),
    .A1(\fetch.bht.bhtTable_tag[13][0] ),
    .A2(\fetch.bht.bhtTable_tag[14][0] ),
    .A3(\fetch.bht.bhtTable_tag[15][0] ),
    .S0(_06617_),
    .S1(_06622_),
    .X(_06908_));
 sky130_fd_sc_hd__mux2_2 _22314_ (.A0(\fetch.bht.bhtTable_tag[10][0] ),
    .A1(\fetch.bht.bhtTable_tag[11][0] ),
    .S(_06644_),
    .X(_06909_));
 sky130_fd_sc_hd__mux2_2 _22315_ (.A0(\fetch.bht.bhtTable_tag[8][0] ),
    .A1(\fetch.bht.bhtTable_tag[9][0] ),
    .S(_06643_),
    .X(_06910_));
 sky130_fd_sc_hd__and2b_2 _22316_ (.A_N(_06730_),
    .B(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__a211o_2 _22317_ (.A1(_06909_),
    .A2(_06685_),
    .B1(_06631_),
    .C1(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__o211a_2 _22318_ (.A1(_06628_),
    .A2(_06908_),
    .B1(_06699_),
    .C1(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__or3_2 _22319_ (.A(io_fetch_address[6]),
    .B(_06907_),
    .C(_06913_),
    .X(_06914_));
 sky130_fd_sc_hd__o21ai_2 _22320_ (.A1(_06907_),
    .A2(_06913_),
    .B1(io_fetch_address[6]),
    .Y(_06915_));
 sky130_fd_sc_hd__and2_2 _22321_ (.A(_06914_),
    .B(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__a21bo_2 _22322_ (.A1(_06707_),
    .A2(\fetch.bht.bhtTable_tag[11][8] ),
    .B1_N(_06649_),
    .X(_06917_));
 sky130_fd_sc_hd__and2b_2 _22323_ (.A_N(_06691_),
    .B(\fetch.bht.bhtTable_tag[10][8] ),
    .X(_06918_));
 sky130_fd_sc_hd__mux2_2 _22324_ (.A0(\fetch.bht.bhtTable_tag[8][8] ),
    .A1(\fetch.bht.bhtTable_tag[9][8] ),
    .S(_06616_),
    .X(_06919_));
 sky130_fd_sc_hd__o221a_2 _22325_ (.A1(_06917_),
    .A2(_06918_),
    .B1(_06675_),
    .B2(_06919_),
    .C1(_06686_),
    .X(_06920_));
 sky130_fd_sc_hd__mux4_2 _22326_ (.A0(\fetch.bht.bhtTable_tag[12][8] ),
    .A1(\fetch.bht.bhtTable_tag[13][8] ),
    .A2(\fetch.bht.bhtTable_tag[14][8] ),
    .A3(\fetch.bht.bhtTable_tag[15][8] ),
    .S0(_06809_),
    .S1(_06649_),
    .X(_06921_));
 sky130_fd_sc_hd__a21o_2 _22327_ (.A1(_06672_),
    .A2(_06921_),
    .B1(_06635_),
    .X(_06922_));
 sky130_fd_sc_hd__mux4_2 _22328_ (.A0(\fetch.bht.bhtTable_tag[4][8] ),
    .A1(\fetch.bht.bhtTable_tag[5][8] ),
    .A2(\fetch.bht.bhtTable_tag[6][8] ),
    .A3(\fetch.bht.bhtTable_tag[7][8] ),
    .S0(_06878_),
    .S1(_06677_),
    .X(_06923_));
 sky130_fd_sc_hd__nand2_2 _22329_ (.A(_06790_),
    .B(_06923_),
    .Y(_06924_));
 sky130_fd_sc_hd__mux4_2 _22330_ (.A0(\fetch.bht.bhtTable_tag[0][8] ),
    .A1(\fetch.bht.bhtTable_tag[1][8] ),
    .A2(\fetch.bht.bhtTable_tag[2][8] ),
    .A3(\fetch.bht.bhtTable_tag[3][8] ),
    .S0(_06878_),
    .S1(_06621_),
    .X(_06925_));
 sky130_fd_sc_hd__a21oi_2 _22331_ (.A1(_06925_),
    .A2(_06687_),
    .B1(_06640_),
    .Y(_06926_));
 sky130_fd_sc_hd__a2bb2o_2 _22332_ (.A1_N(_06920_),
    .A2_N(_06922_),
    .B1(_06924_),
    .B2(_06926_),
    .X(_06927_));
 sky130_fd_sc_hd__xnor2_2 _22333_ (.A(io_fetch_address[14]),
    .B(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__mux2_2 _22334_ (.A0(\fetch.bht.bhtTable_tag[6][10] ),
    .A1(\fetch.bht.bhtTable_tag[7][10] ),
    .S(_06680_),
    .X(_06929_));
 sky130_fd_sc_hd__mux2_2 _22335_ (.A0(\fetch.bht.bhtTable_tag[4][10] ),
    .A1(\fetch.bht.bhtTable_tag[5][10] ),
    .S(_06706_),
    .X(_06930_));
 sky130_fd_sc_hd__and2b_2 _22336_ (.A_N(_06684_),
    .B(_06930_),
    .X(_06931_));
 sky130_fd_sc_hd__a211oi_2 _22337_ (.A1(_06685_),
    .A2(_06929_),
    .B1(_06627_),
    .C1(_06931_),
    .Y(_06932_));
 sky130_fd_sc_hd__mux2_2 _22338_ (.A0(\fetch.bht.bhtTable_tag[2][10] ),
    .A1(\fetch.bht.bhtTable_tag[3][10] ),
    .S(_06644_),
    .X(_06933_));
 sky130_fd_sc_hd__mux2_2 _22339_ (.A0(\fetch.bht.bhtTable_tag[0][10] ),
    .A1(\fetch.bht.bhtTable_tag[1][10] ),
    .S(_06643_),
    .X(_06934_));
 sky130_fd_sc_hd__and2b_2 _22340_ (.A_N(_06730_),
    .B(_06934_),
    .X(_06935_));
 sky130_fd_sc_hd__a211oi_2 _22341_ (.A1(_06933_),
    .A2(_06678_),
    .B1(_06631_),
    .C1(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__mux4_2 _22342_ (.A0(\fetch.bht.bhtTable_tag[8][10] ),
    .A1(\fetch.bht.bhtTable_tag[9][10] ),
    .A2(\fetch.bht.bhtTable_tag[10][10] ),
    .A3(\fetch.bht.bhtTable_tag[11][10] ),
    .S0(_06878_),
    .S1(_06621_),
    .X(_06937_));
 sky130_fd_sc_hd__mux2_2 _22343_ (.A0(\fetch.bht.bhtTable_tag[12][10] ),
    .A1(\fetch.bht.bhtTable_tag[13][10] ),
    .S(_06643_),
    .X(_06938_));
 sky130_fd_sc_hd__and2b_2 _22344_ (.A_N(_06730_),
    .B(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__mux2_2 _22345_ (.A0(\fetch.bht.bhtTable_tag[14][10] ),
    .A1(\fetch.bht.bhtTable_tag[15][10] ),
    .S(_06809_),
    .X(_06940_));
 sky130_fd_sc_hd__a21o_2 _22346_ (.A1(_06940_),
    .A2(_06650_),
    .B1(_06686_),
    .X(_06941_));
 sky130_fd_sc_hd__o221ai_2 _22347_ (.A1(_06790_),
    .A2(_06937_),
    .B1(_06939_),
    .B2(_06941_),
    .C1(_06640_),
    .Y(_06942_));
 sky130_fd_sc_hd__o31a_2 _22348_ (.A1(_06641_),
    .A2(_06932_),
    .A3(_06936_),
    .B1(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__xnor2_2 _22349_ (.A(io_fetch_address[16]),
    .B(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__mux4_2 _22350_ (.A0(\fetch.bht.bhtTable_tag[0][14] ),
    .A1(\fetch.bht.bhtTable_tag[1][14] ),
    .A2(\fetch.bht.bhtTable_tag[2][14] ),
    .A3(\fetch.bht.bhtTable_tag[3][14] ),
    .S0(_06616_),
    .S1(_06621_),
    .X(_06945_));
 sky130_fd_sc_hd__nor2_2 _22351_ (.A(_06672_),
    .B(_06945_),
    .Y(_06946_));
 sky130_fd_sc_hd__mux2_2 _22352_ (.A0(\fetch.bht.bhtTable_tag[4][14] ),
    .A1(\fetch.bht.bhtTable_tag[5][14] ),
    .S(_06615_),
    .X(_06947_));
 sky130_fd_sc_hd__or2b_2 _22353_ (.A(_06649_),
    .B_N(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__mux2_2 _22354_ (.A0(\fetch.bht.bhtTable_tag[6][14] ),
    .A1(\fetch.bht.bhtTable_tag[7][14] ),
    .S(_06706_),
    .X(_06949_));
 sky130_fd_sc_hd__nand2_2 _22355_ (.A(_06949_),
    .B(_06677_),
    .Y(_06950_));
 sky130_fd_sc_hd__a31o_2 _22356_ (.A1(_06948_),
    .A2(_06672_),
    .A3(_06950_),
    .B1(_06640_),
    .X(_06951_));
 sky130_fd_sc_hd__mux4_2 _22357_ (.A0(\fetch.bht.bhtTable_tag[8][14] ),
    .A1(\fetch.bht.bhtTable_tag[9][14] ),
    .A2(\fetch.bht.bhtTable_tag[10][14] ),
    .A3(\fetch.bht.bhtTable_tag[11][14] ),
    .S0(_06679_),
    .S1(_06620_),
    .X(_06952_));
 sky130_fd_sc_hd__mux4_2 _22358_ (.A0(\fetch.bht.bhtTable_tag[12][14] ),
    .A1(\fetch.bht.bhtTable_tag[13][14] ),
    .A2(\fetch.bht.bhtTable_tag[14][14] ),
    .A3(\fetch.bht.bhtTable_tag[15][14] ),
    .S0(_06679_),
    .S1(_06620_),
    .X(_06953_));
 sky130_fd_sc_hd__mux2_2 _22359_ (.A0(_06952_),
    .A1(_06953_),
    .S(_00002_),
    .X(_06954_));
 sky130_fd_sc_hd__a2bb2o_2 _22360_ (.A1_N(_06946_),
    .A2_N(_06951_),
    .B1(_06640_),
    .B2(_06954_),
    .X(_06955_));
 sky130_fd_sc_hd__xnor2_2 _22361_ (.A(io_fetch_address[20]),
    .B(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__mux4_2 _22362_ (.A0(\fetch.bht.bhtTable_tag[0][2] ),
    .A1(\fetch.bht.bhtTable_tag[1][2] ),
    .A2(\fetch.bht.bhtTable_tag[2][2] ),
    .A3(\fetch.bht.bhtTable_tag[3][2] ),
    .S0(_06679_),
    .S1(_06620_),
    .X(_06957_));
 sky130_fd_sc_hd__mux4_2 _22363_ (.A0(\fetch.bht.bhtTable_tag[4][2] ),
    .A1(\fetch.bht.bhtTable_tag[5][2] ),
    .A2(\fetch.bht.bhtTable_tag[6][2] ),
    .A3(\fetch.bht.bhtTable_tag[7][2] ),
    .S0(_06679_),
    .S1(_06620_),
    .X(_06958_));
 sky130_fd_sc_hd__mux2_2 _22364_ (.A0(_06957_),
    .A1(_06958_),
    .S(_00002_),
    .X(_06959_));
 sky130_fd_sc_hd__mux4_2 _22365_ (.A0(\fetch.bht.bhtTable_tag[12][2] ),
    .A1(\fetch.bht.bhtTable_tag[13][2] ),
    .A2(\fetch.bht.bhtTable_tag[14][2] ),
    .A3(\fetch.bht.bhtTable_tag[15][2] ),
    .S0(_06615_),
    .S1(_06620_),
    .X(_06960_));
 sky130_fd_sc_hd__mux4_2 _22366_ (.A0(\fetch.bht.bhtTable_tag[8][2] ),
    .A1(\fetch.bht.bhtTable_tag[9][2] ),
    .A2(\fetch.bht.bhtTable_tag[10][2] ),
    .A3(\fetch.bht.bhtTable_tag[11][2] ),
    .S0(_06615_),
    .S1(_06620_),
    .X(_06961_));
 sky130_fd_sc_hd__mux2_2 _22367_ (.A0(_06960_),
    .A1(_06961_),
    .S(_06626_),
    .X(_06962_));
 sky130_fd_sc_hd__mux2_2 _22368_ (.A0(_06959_),
    .A1(_06962_),
    .S(_06640_),
    .X(_06963_));
 sky130_fd_sc_hd__xnor2_2 _22369_ (.A(io_fetch_address[8]),
    .B(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__nand2_2 _22370_ (.A(_06956_),
    .B(_06964_),
    .Y(_06965_));
 sky130_fd_sc_hd__mux4_2 _22371_ (.A0(\fetch.bht.bhtTable_tag[0][16] ),
    .A1(\fetch.bht.bhtTable_tag[1][16] ),
    .A2(\fetch.bht.bhtTable_tag[2][16] ),
    .A3(\fetch.bht.bhtTable_tag[3][16] ),
    .S0(_06878_),
    .S1(_06621_),
    .X(_06966_));
 sky130_fd_sc_hd__mux4_2 _22372_ (.A0(\fetch.bht.bhtTable_tag[4][16] ),
    .A1(\fetch.bht.bhtTable_tag[5][16] ),
    .A2(\fetch.bht.bhtTable_tag[6][16] ),
    .A3(\fetch.bht.bhtTable_tag[7][16] ),
    .S0(_06878_),
    .S1(_06621_),
    .X(_06967_));
 sky130_fd_sc_hd__mux2_2 _22373_ (.A0(_06966_),
    .A1(_06967_),
    .S(_06631_),
    .X(_06968_));
 sky130_fd_sc_hd__mux2_2 _22374_ (.A0(\fetch.bht.bhtTable_tag[12][16] ),
    .A1(\fetch.bht.bhtTable_tag[13][16] ),
    .S(_06643_),
    .X(_06969_));
 sky130_fd_sc_hd__and2b_2 _22375_ (.A_N(_06730_),
    .B(_06969_),
    .X(_06970_));
 sky130_fd_sc_hd__mux2_2 _22376_ (.A0(\fetch.bht.bhtTable_tag[14][16] ),
    .A1(\fetch.bht.bhtTable_tag[15][16] ),
    .S(_06809_),
    .X(_06971_));
 sky130_fd_sc_hd__a21o_2 _22377_ (.A1(_06971_),
    .A2(_06730_),
    .B1(_06686_),
    .X(_06972_));
 sky130_fd_sc_hd__mux4_2 _22378_ (.A0(\fetch.bht.bhtTable_tag[8][16] ),
    .A1(\fetch.bht.bhtTable_tag[9][16] ),
    .A2(\fetch.bht.bhtTable_tag[10][16] ),
    .A3(\fetch.bht.bhtTable_tag[11][16] ),
    .S0(_06691_),
    .S1(_06677_),
    .X(_06973_));
 sky130_fd_sc_hd__o221a_2 _22379_ (.A1(_06970_),
    .A2(_06972_),
    .B1(_06973_),
    .B2(_06790_),
    .C1(_06641_),
    .X(_06974_));
 sky130_fd_sc_hd__a21oi_2 _22380_ (.A1(_06968_),
    .A2(_06636_),
    .B1(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__xnor2_2 _22381_ (.A(io_fetch_address[22]),
    .B(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__or4_2 _22382_ (.A(_06928_),
    .B(_06944_),
    .C(_06965_),
    .D(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__mux2_2 _22383_ (.A0(\fetch.bht.bhtTable_tag[6][9] ),
    .A1(\fetch.bht.bhtTable_tag[7][9] ),
    .S(_06617_),
    .X(_06978_));
 sky130_fd_sc_hd__mux2_2 _22384_ (.A0(\fetch.bht.bhtTable_tag[4][9] ),
    .A1(\fetch.bht.bhtTable_tag[5][9] ),
    .S(_06878_),
    .X(_06979_));
 sky130_fd_sc_hd__and2b_2 _22385_ (.A_N(_06622_),
    .B(_06979_),
    .X(_06980_));
 sky130_fd_sc_hd__a211oi_2 _22386_ (.A1(_06623_),
    .A2(_06978_),
    .B1(_06687_),
    .C1(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__mux4_2 _22387_ (.A0(\fetch.bht.bhtTable_tag[0][9] ),
    .A1(\fetch.bht.bhtTable_tag[1][9] ),
    .A2(\fetch.bht.bhtTable_tag[2][9] ),
    .A3(\fetch.bht.bhtTable_tag[3][9] ),
    .S0(_06754_),
    .S1(_06622_),
    .X(_06982_));
 sky130_fd_sc_hd__nor2_2 _22388_ (.A(_06673_),
    .B(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__mux4_2 _22389_ (.A0(\fetch.bht.bhtTable_tag[8][9] ),
    .A1(\fetch.bht.bhtTable_tag[9][9] ),
    .A2(\fetch.bht.bhtTable_tag[10][9] ),
    .A3(\fetch.bht.bhtTable_tag[11][9] ),
    .S0(_06754_),
    .S1(_06675_),
    .X(_06984_));
 sky130_fd_sc_hd__mux2_2 _22390_ (.A0(\fetch.bht.bhtTable_tag[14][9] ),
    .A1(\fetch.bht.bhtTable_tag[15][9] ),
    .S(_06707_),
    .X(_06985_));
 sky130_fd_sc_hd__mux2_2 _22391_ (.A0(\fetch.bht.bhtTable_tag[12][9] ),
    .A1(\fetch.bht.bhtTable_tag[13][9] ),
    .S(_06706_),
    .X(_06986_));
 sky130_fd_sc_hd__and2b_2 _22392_ (.A_N(_06684_),
    .B(_06986_),
    .X(_06987_));
 sky130_fd_sc_hd__a211o_2 _22393_ (.A1(_06678_),
    .A2(_06985_),
    .B1(_06627_),
    .C1(_06987_),
    .X(_06988_));
 sky130_fd_sc_hd__o211ai_2 _22394_ (.A1(_06673_),
    .A2(_06984_),
    .B1(_06641_),
    .C1(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__o31a_2 _22395_ (.A1(_06699_),
    .A2(_06981_),
    .A3(_06983_),
    .B1(_06989_),
    .X(_06990_));
 sky130_fd_sc_hd__xnor2_2 _22396_ (.A(io_fetch_address[15]),
    .B(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__mux4_2 _22397_ (.A0(\fetch.bht.bhtTable_tag[8][21] ),
    .A1(\fetch.bht.bhtTable_tag[9][21] ),
    .A2(\fetch.bht.bhtTable_tag[10][21] ),
    .A3(\fetch.bht.bhtTable_tag[11][21] ),
    .S0(_06707_),
    .S1(_06730_),
    .X(_06992_));
 sky130_fd_sc_hd__mux2_2 _22398_ (.A0(\fetch.bht.bhtTable_tag[12][21] ),
    .A1(\fetch.bht.bhtTable_tag[13][21] ),
    .S(_06809_),
    .X(_06993_));
 sky130_fd_sc_hd__and2b_2 _22399_ (.A_N(_06650_),
    .B(_06993_),
    .X(_06994_));
 sky130_fd_sc_hd__mux2_2 _22400_ (.A0(\fetch.bht.bhtTable_tag[14][21] ),
    .A1(\fetch.bht.bhtTable_tag[15][21] ),
    .S(_06616_),
    .X(_06995_));
 sky130_fd_sc_hd__a21o_2 _22401_ (.A1(_06995_),
    .A2(_06675_),
    .B1(_06686_),
    .X(_06996_));
 sky130_fd_sc_hd__o22a_2 _22402_ (.A1(_06790_),
    .A2(_06992_),
    .B1(_06994_),
    .B2(_06996_),
    .X(_06997_));
 sky130_fd_sc_hd__mux4_2 _22403_ (.A0(\fetch.bht.bhtTable_tag[0][21] ),
    .A1(\fetch.bht.bhtTable_tag[1][21] ),
    .A2(\fetch.bht.bhtTable_tag[2][21] ),
    .A3(\fetch.bht.bhtTable_tag[3][21] ),
    .S0(_06617_),
    .S1(_06622_),
    .X(_06998_));
 sky130_fd_sc_hd__nor2_2 _22404_ (.A(_06673_),
    .B(_06998_),
    .Y(_06999_));
 sky130_fd_sc_hd__mux2_2 _22405_ (.A0(\fetch.bht.bhtTable_tag[4][21] ),
    .A1(\fetch.bht.bhtTable_tag[5][21] ),
    .S(_06809_),
    .X(_07000_));
 sky130_fd_sc_hd__or2b_2 _22406_ (.A(_06650_),
    .B_N(_07000_),
    .X(_07001_));
 sky130_fd_sc_hd__mux2_2 _22407_ (.A0(\fetch.bht.bhtTable_tag[6][21] ),
    .A1(\fetch.bht.bhtTable_tag[7][21] ),
    .S(_06707_),
    .X(_07002_));
 sky130_fd_sc_hd__nand2_2 _22408_ (.A(_07002_),
    .B(_06678_),
    .Y(_07003_));
 sky130_fd_sc_hd__a31o_2 _22409_ (.A1(_07001_),
    .A2(_07003_),
    .A3(_06790_),
    .B1(_06640_),
    .X(_07004_));
 sky130_fd_sc_hd__o2bb2a_2 _22410_ (.A1_N(_06699_),
    .A2_N(_06997_),
    .B1(_06999_),
    .B2(_07004_),
    .X(_07005_));
 sky130_fd_sc_hd__xor2_2 _22411_ (.A(io_fetch_address[27]),
    .B(_07005_),
    .X(_07006_));
 sky130_fd_sc_hd__or2b_2 _22412_ (.A(_06991_),
    .B_N(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__mux4_2 _22413_ (.A0(\fetch.bht.bhtTable_tag[0][1] ),
    .A1(\fetch.bht.bhtTable_tag[1][1] ),
    .A2(\fetch.bht.bhtTable_tag[2][1] ),
    .A3(\fetch.bht.bhtTable_tag[3][1] ),
    .S0(_06680_),
    .S1(_06684_),
    .X(_07008_));
 sky130_fd_sc_hd__mux4_2 _22414_ (.A0(\fetch.bht.bhtTable_tag[4][1] ),
    .A1(\fetch.bht.bhtTable_tag[5][1] ),
    .A2(\fetch.bht.bhtTable_tag[6][1] ),
    .A3(\fetch.bht.bhtTable_tag[7][1] ),
    .S0(_06680_),
    .S1(_06684_),
    .X(_07009_));
 sky130_fd_sc_hd__mux2_2 _22415_ (.A0(_07008_),
    .A1(_07009_),
    .S(_06790_),
    .X(_07010_));
 sky130_fd_sc_hd__mux4_2 _22416_ (.A0(\fetch.bht.bhtTable_tag[8][1] ),
    .A1(\fetch.bht.bhtTable_tag[9][1] ),
    .A2(\fetch.bht.bhtTable_tag[10][1] ),
    .A3(\fetch.bht.bhtTable_tag[11][1] ),
    .S0(_06674_),
    .S1(_06650_),
    .X(_07011_));
 sky130_fd_sc_hd__mux2_2 _22417_ (.A0(\fetch.bht.bhtTable_tag[12][1] ),
    .A1(\fetch.bht.bhtTable_tag[13][1] ),
    .S(_06691_),
    .X(_07012_));
 sky130_fd_sc_hd__mux2_2 _22418_ (.A0(\fetch.bht.bhtTable_tag[14][1] ),
    .A1(\fetch.bht.bhtTable_tag[15][1] ),
    .S(_06679_),
    .X(_07013_));
 sky130_fd_sc_hd__or2b_2 _22419_ (.A(_07013_),
    .B_N(_06677_),
    .X(_07014_));
 sky130_fd_sc_hd__o211a_2 _22420_ (.A1(_06690_),
    .A2(_07012_),
    .B1(_06672_),
    .C1(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__a211oi_2 _22421_ (.A1(_06628_),
    .A2(_07011_),
    .B1(_06635_),
    .C1(_07015_),
    .Y(_07016_));
 sky130_fd_sc_hd__o21ba_2 _22422_ (.A1(_06699_),
    .A2(_07010_),
    .B1_N(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__xor2_2 _22423_ (.A(io_fetch_address[7]),
    .B(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__mux4_2 _22424_ (.A0(\fetch.bht.bhtTable_tag[0][12] ),
    .A1(\fetch.bht.bhtTable_tag[1][12] ),
    .A2(\fetch.bht.bhtTable_tag[2][12] ),
    .A3(\fetch.bht.bhtTable_tag[3][12] ),
    .S0(_06644_),
    .S1(_06650_),
    .X(_07019_));
 sky130_fd_sc_hd__mux2_2 _22425_ (.A0(\fetch.bht.bhtTable_tag[4][12] ),
    .A1(\fetch.bht.bhtTable_tag[5][12] ),
    .S(_06878_),
    .X(_07020_));
 sky130_fd_sc_hd__and2b_2 _22426_ (.A_N(_06622_),
    .B(_07020_),
    .X(_07021_));
 sky130_fd_sc_hd__mux2_2 _22427_ (.A0(\fetch.bht.bhtTable_tag[6][12] ),
    .A1(\fetch.bht.bhtTable_tag[7][12] ),
    .S(_06691_),
    .X(_07022_));
 sky130_fd_sc_hd__a21o_2 _22428_ (.A1(_07022_),
    .A2(_06690_),
    .B1(_06627_),
    .X(_07023_));
 sky130_fd_sc_hd__o22a_2 _22429_ (.A1(_06790_),
    .A2(_07019_),
    .B1(_07021_),
    .B2(_07023_),
    .X(_07024_));
 sky130_fd_sc_hd__or2b_2 _22430_ (.A(\fetch.bht.bhtTable_tag[15][12] ),
    .B_N(_06707_),
    .X(_07025_));
 sky130_fd_sc_hd__o211a_2 _22431_ (.A1(_06700_),
    .A2(\fetch.bht.bhtTable_tag[14][12] ),
    .B1(_06675_),
    .C1(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__mux2_2 _22432_ (.A0(\fetch.bht.bhtTable_tag[12][12] ),
    .A1(\fetch.bht.bhtTable_tag[13][12] ),
    .S(_06616_),
    .X(_07027_));
 sky130_fd_sc_hd__and2b_2 _22433_ (.A_N(_06675_),
    .B(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__mux2_2 _22434_ (.A0(\fetch.bht.bhtTable_tag[10][12] ),
    .A1(\fetch.bht.bhtTable_tag[11][12] ),
    .S(_06691_),
    .X(_07029_));
 sky130_fd_sc_hd__mux2_2 _22435_ (.A0(\fetch.bht.bhtTable_tag[8][12] ),
    .A1(\fetch.bht.bhtTable_tag[9][12] ),
    .S(_06679_),
    .X(_07030_));
 sky130_fd_sc_hd__and2b_2 _22436_ (.A_N(_06621_),
    .B(_07030_),
    .X(_07031_));
 sky130_fd_sc_hd__a211o_2 _22437_ (.A1(_07029_),
    .A2(_06690_),
    .B1(_06672_),
    .C1(_07031_),
    .X(_07032_));
 sky130_fd_sc_hd__o311a_2 _22438_ (.A1(_06687_),
    .A2(_07026_),
    .A3(_07028_),
    .B1(_06641_),
    .C1(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__a21oi_2 _22439_ (.A1(_06636_),
    .A2(_07024_),
    .B1(_07033_),
    .Y(_07034_));
 sky130_fd_sc_hd__xor2_2 _22440_ (.A(io_fetch_address[18]),
    .B(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__a31oi_2 _22441_ (.A1(_06641_),
    .A2(_06811_),
    .A3(_06815_),
    .B1(_06819_),
    .Y(_07036_));
 sky130_fd_sc_hd__or2b_2 _22442_ (.A(_07036_),
    .B_N(io_fetch_address[26]),
    .X(_07037_));
 sky130_fd_sc_hd__and3b_2 _22443_ (.A_N(_06754_),
    .B(\fetch.btb.btbTable[10][1] ),
    .C(\fetch.bht.bhtTable_valid[10] ),
    .X(_07038_));
 sky130_fd_sc_hd__a311o_2 _22444_ (.A1(_06618_),
    .A2(\fetch.btb.btbTable[11][1] ),
    .A3(\fetch.bht.bhtTable_valid[11] ),
    .B1(_07038_),
    .C1(_06631_),
    .X(_07039_));
 sky130_fd_sc_hd__and3b_2 _22445_ (.A_N(_06617_),
    .B(\fetch.btb.btbTable[14][1] ),
    .C(\fetch.bht.bhtTable_valid[14] ),
    .X(_07040_));
 sky130_fd_sc_hd__a311o_2 _22446_ (.A1(_06645_),
    .A2(\fetch.btb.btbTable[15][1] ),
    .A3(\fetch.bht.bhtTable_valid[15] ),
    .B1(_06627_),
    .C1(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__and3b_2 _22447_ (.A_N(_06674_),
    .B(\fetch.btb.btbTable[6][1] ),
    .C(\fetch.bht.bhtTable_valid[6] ),
    .X(_07042_));
 sky130_fd_sc_hd__a31o_2 _22448_ (.A1(_06674_),
    .A2(\fetch.btb.btbTable[7][1] ),
    .A3(\fetch.bht.bhtTable_valid[7] ),
    .B1(_06626_),
    .X(_07043_));
 sky130_fd_sc_hd__o21ai_2 _22449_ (.A1(_07042_),
    .A2(_07043_),
    .B1(_06635_),
    .Y(_07044_));
 sky130_fd_sc_hd__and3b_2 _22450_ (.A_N(_06674_),
    .B(\fetch.btb.btbTable[2][1] ),
    .C(\fetch.bht.bhtTable_valid[2] ),
    .X(_07045_));
 sky130_fd_sc_hd__a311oi_2 _22451_ (.A1(_06645_),
    .A2(\fetch.btb.btbTable[3][1] ),
    .A3(\fetch.bht.bhtTable_valid[3] ),
    .B1(_07045_),
    .C1(_06631_),
    .Y(_07046_));
 sky130_fd_sc_hd__o21ai_2 _22452_ (.A1(_07044_),
    .A2(_07046_),
    .B1(_06623_),
    .Y(_07047_));
 sky130_fd_sc_hd__a31o_2 _22453_ (.A1(_06699_),
    .A2(_07039_),
    .A3(_07041_),
    .B1(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__and3b_2 _22454_ (.A_N(_06617_),
    .B(\fetch.btb.btbTable[12][1] ),
    .C(\fetch.bht.bhtTable_valid[12] ),
    .X(_07049_));
 sky130_fd_sc_hd__a311o_2 _22455_ (.A1(_06618_),
    .A2(\fetch.btb.btbTable[13][1] ),
    .A3(\fetch.bht.bhtTable_valid[13] ),
    .B1(_06687_),
    .C1(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__and3b_2 _22456_ (.A_N(_06754_),
    .B(\fetch.btb.btbTable[8][1] ),
    .C(\fetch.bht.bhtTable_valid[8] ),
    .X(_07051_));
 sky130_fd_sc_hd__a311o_2 _22457_ (.A1(_06645_),
    .A2(\fetch.btb.btbTable[9][1] ),
    .A3(\fetch.bht.bhtTable_valid[9] ),
    .B1(_07051_),
    .C1(_06631_),
    .X(_07052_));
 sky130_fd_sc_hd__and3b_2 _22458_ (.A_N(_06616_),
    .B(\fetch.btb.btbTable[4][1] ),
    .C(\fetch.bht.bhtTable_valid[4] ),
    .X(_07053_));
 sky130_fd_sc_hd__a311o_2 _22459_ (.A1(_06754_),
    .A2(\fetch.btb.btbTable[5][1] ),
    .A3(\fetch.bht.bhtTable_valid[5] ),
    .B1(_06686_),
    .C1(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__and3b_2 _22460_ (.A_N(_06809_),
    .B(\fetch.bht.bhtTable_valid[0] ),
    .C(\fetch.btb.btbTable[0][1] ),
    .X(_07055_));
 sky130_fd_sc_hd__a311o_2 _22461_ (.A1(\fetch.btb.btbTable[1][1] ),
    .A2(_06674_),
    .A3(\fetch.bht.bhtTable_valid[1] ),
    .B1(_07055_),
    .C1(_00002_),
    .X(_07056_));
 sky130_fd_sc_hd__a31o_2 _22462_ (.A1(_06635_),
    .A2(_07054_),
    .A3(_07056_),
    .B1(_06651_),
    .X(_07057_));
 sky130_fd_sc_hd__a31o_2 _22463_ (.A1(_06699_),
    .A2(_07050_),
    .A3(_07052_),
    .B1(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__and3_2 _22464_ (.A(_07037_),
    .B(_07048_),
    .C(_07058_),
    .X(_07059_));
 sky130_fd_sc_hd__and3b_2 _22465_ (.A_N(_07018_),
    .B(_07035_),
    .C(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__or4b_2 _22466_ (.A(_06916_),
    .B(_06977_),
    .C(_07007_),
    .D_N(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__or4_2 _22467_ (.A(_06891_),
    .B(_06893_),
    .C(_06898_),
    .D(_07061_),
    .X(_07062_));
 sky130_fd_sc_hd__o41a_2 _22468_ (.A1(_06720_),
    .A2(_06769_),
    .A3(_06822_),
    .A4(_07062_),
    .B1(_03591_),
    .X(_07063_));
 sky130_fd_sc_hd__buf_1 _22469_ (.A(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__a2bb2o_2 _22470_ (.A1_N(_10758_),
    .A2_N(_10914_),
    .B1(_07064_),
    .B2(_03590_),
    .X(_07065_));
 sky130_fd_sc_hd__buf_1 _22471_ (.A(_06619_),
    .X(_07066_));
 sky130_fd_sc_hd__buf_1 _22472_ (.A(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__buf_1 _22473_ (.A(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__buf_1 _22474_ (.A(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__buf_1 _22475_ (.A(_06661_),
    .X(_07070_));
 sky130_fd_sc_hd__buf_1 _22476_ (.A(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__buf_1 _22477_ (.A(_07071_),
    .X(_07072_));
 sky130_fd_sc_hd__mux4_2 _22478_ (.A0(\fetch.bht.bhtTable_target_pc[8][0] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][0] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][0] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][0] ),
    .S0(_07069_),
    .S1(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__mux4_2 _22479_ (.A0(\fetch.bht.bhtTable_target_pc[12][0] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][0] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][0] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][0] ),
    .S0(_07069_),
    .S1(_07072_),
    .X(_07074_));
 sky130_fd_sc_hd__buf_1 _22480_ (.A(_06633_),
    .X(_07075_));
 sky130_fd_sc_hd__buf_1 _22481_ (.A(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__mux2_2 _22482_ (.A0(_07073_),
    .A1(_07074_),
    .S(_07076_),
    .X(_07077_));
 sky130_fd_sc_hd__mux4_2 _22483_ (.A0(\fetch.bht.bhtTable_target_pc[4][0] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][0] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][0] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][0] ),
    .S0(_07069_),
    .S1(_07072_),
    .X(_07078_));
 sky130_fd_sc_hd__mux4_2 _22484_ (.A0(\fetch.bht.bhtTable_target_pc[0][0] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][0] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][0] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][0] ),
    .S0(_07069_),
    .S1(_07072_),
    .X(_07079_));
 sky130_fd_sc_hd__buf_1 _22485_ (.A(_06629_),
    .X(_07080_));
 sky130_fd_sc_hd__buf_1 _22486_ (.A(_07080_),
    .X(_07081_));
 sky130_fd_sc_hd__buf_1 _22487_ (.A(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__mux2_2 _22488_ (.A0(_07078_),
    .A1(_07079_),
    .S(_07082_),
    .X(_07083_));
 sky130_fd_sc_hd__buf_1 _22489_ (.A(_06637_),
    .X(_07084_));
 sky130_fd_sc_hd__buf_1 _22490_ (.A(_07084_),
    .X(_07085_));
 sky130_fd_sc_hd__mux2_2 _22491_ (.A0(_07077_),
    .A1(_07083_),
    .S(_07085_),
    .X(_07086_));
 sky130_fd_sc_hd__or4_2 _22492_ (.A(_06720_),
    .B(_06769_),
    .C(_06822_),
    .D(_07062_),
    .X(_07087_));
 sky130_fd_sc_hd__nor2_2 _22493_ (.A(_10757_),
    .B(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__buf_1 _22494_ (.A(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__buf_1 _22495_ (.A(_10757_),
    .X(_07090_));
 sky130_fd_sc_hd__buf_1 _22496_ (.A(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__a21o_2 _22497_ (.A1(\execute.io_target_pc[0] ),
    .A2(_07091_),
    .B1(_06041_),
    .X(_07092_));
 sky130_fd_sc_hd__a21oi_2 _22498_ (.A1(_07086_),
    .A2(_07089_),
    .B1(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__inv_2 _22499_ (.A(\csr.io_mret_vector[0] ),
    .Y(_07094_));
 sky130_fd_sc_hd__a211o_2 _22500_ (.A1(_06041_),
    .A2(_07094_),
    .B1(_06481_),
    .C1(_07065_),
    .X(_07095_));
 sky130_fd_sc_hd__o2bb2a_2 _22501_ (.A1_N(io_fetch_address[0]),
    .A2_N(_07065_),
    .B1(_07093_),
    .B2(_07095_),
    .X(_07096_));
 sky130_fd_sc_hd__nor2_2 _22502_ (.A(_03580_),
    .B(_07096_),
    .Y(_01252_));
 sky130_fd_sc_hd__buf_1 _22503_ (.A(_06740_),
    .X(_07097_));
 sky130_fd_sc_hd__buf_1 _22504_ (.A(_07066_),
    .X(_07098_));
 sky130_fd_sc_hd__buf_1 _22505_ (.A(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__buf_1 _22506_ (.A(_07070_),
    .X(_07100_));
 sky130_fd_sc_hd__buf_1 _22507_ (.A(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__mux4_2 _22508_ (.A0(\fetch.bht.bhtTable_target_pc[12][1] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][1] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][1] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][1] ),
    .S0(_07099_),
    .S1(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__buf_1 _22509_ (.A(_07100_),
    .X(_07103_));
 sky130_fd_sc_hd__mux4_2 _22510_ (.A0(\fetch.bht.bhtTable_target_pc[8][1] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][1] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][1] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][1] ),
    .S0(_07099_),
    .S1(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__mux2_2 _22511_ (.A0(_07102_),
    .A1(_07104_),
    .S(_07082_),
    .X(_07105_));
 sky130_fd_sc_hd__buf_1 _22512_ (.A(_07066_),
    .X(_07106_));
 sky130_fd_sc_hd__buf_1 _22513_ (.A(_07106_),
    .X(_07107_));
 sky130_fd_sc_hd__buf_1 _22514_ (.A(_07107_),
    .X(_07108_));
 sky130_fd_sc_hd__mux2_2 _22515_ (.A0(\fetch.bht.bhtTable_target_pc[2][1] ),
    .A1(\fetch.bht.bhtTable_target_pc[3][1] ),
    .S(_07108_),
    .X(_07109_));
 sky130_fd_sc_hd__buf_1 _22516_ (.A(_07070_),
    .X(_07110_));
 sky130_fd_sc_hd__buf_1 _22517_ (.A(_07110_),
    .X(_07111_));
 sky130_fd_sc_hd__buf_1 _22518_ (.A(_07111_),
    .X(_07112_));
 sky130_fd_sc_hd__buf_1 _22519_ (.A(_06661_),
    .X(_07113_));
 sky130_fd_sc_hd__buf_1 _22520_ (.A(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__buf_1 _22521_ (.A(_07114_),
    .X(_07115_));
 sky130_fd_sc_hd__mux2_2 _22522_ (.A0(\fetch.bht.bhtTable_target_pc[0][1] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][1] ),
    .S(_07099_),
    .X(_07116_));
 sky130_fd_sc_hd__and2b_2 _22523_ (.A_N(_07115_),
    .B(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__a211oi_2 _22524_ (.A1(_07109_),
    .A2(_07112_),
    .B1(_07076_),
    .C1(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__buf_1 _22525_ (.A(_07067_),
    .X(_07119_));
 sky130_fd_sc_hd__mux2_2 _22526_ (.A0(\fetch.bht.bhtTable_target_pc[4][1] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][1] ),
    .S(_07119_),
    .X(_07120_));
 sky130_fd_sc_hd__or2b_2 _22527_ (.A(_07072_),
    .B_N(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__buf_1 _22528_ (.A(_06633_),
    .X(_07122_));
 sky130_fd_sc_hd__buf_1 _22529_ (.A(_07068_),
    .X(_07123_));
 sky130_fd_sc_hd__mux2_2 _22530_ (.A0(\fetch.bht.bhtTable_target_pc[6][1] ),
    .A1(\fetch.bht.bhtTable_target_pc[7][1] ),
    .S(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__buf_1 _22531_ (.A(_07101_),
    .X(_07125_));
 sky130_fd_sc_hd__nand2_2 _22532_ (.A(_07124_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__buf_1 _22533_ (.A(_06740_),
    .X(_07127_));
 sky130_fd_sc_hd__a31o_2 _22534_ (.A1(_07121_),
    .A2(_07122_),
    .A3(_07126_),
    .B1(_07127_),
    .X(_07128_));
 sky130_fd_sc_hd__o2bb2a_2 _22535_ (.A1_N(_07097_),
    .A2_N(_07105_),
    .B1(_07118_),
    .B2(_07128_),
    .X(_07129_));
 sky130_fd_sc_hd__buf_1 _22536_ (.A(_07087_),
    .X(_07130_));
 sky130_fd_sc_hd__a21oi_2 _22537_ (.A1(\execute.io_target_pc[1] ),
    .A2(_07091_),
    .B1(_06041_),
    .Y(_07131_));
 sky130_fd_sc_hd__o31a_2 _22538_ (.A1(_07129_),
    .A2(_07091_),
    .A3(_07130_),
    .B1(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__inv_2 _22539_ (.A(\csr.io_mret_vector[1] ),
    .Y(_07133_));
 sky130_fd_sc_hd__a211o_2 _22540_ (.A1(_06041_),
    .A2(_07133_),
    .B1(_06481_),
    .C1(_07065_),
    .X(_07134_));
 sky130_fd_sc_hd__o2bb2a_2 _22541_ (.A1_N(io_fetch_address[1]),
    .A2_N(_07065_),
    .B1(_07132_),
    .B2(_07134_),
    .X(_07135_));
 sky130_fd_sc_hd__nor2_2 _22542_ (.A(_03580_),
    .B(_07135_),
    .Y(_01253_));
 sky130_fd_sc_hd__and3_2 _22543_ (.A(\csr.minstret[30] ),
    .B(\csr.minstret[31] ),
    .C(_06417_),
    .X(_07136_));
 sky130_fd_sc_hd__a31o_2 _22544_ (.A1(\csr._minstret_T_3[32] ),
    .A2(\csr.minstret[31] ),
    .A3(_06420_),
    .B1(_06422_),
    .X(_07137_));
 sky130_fd_sc_hd__o21ba_2 _22545_ (.A1(\csr._minstret_T_3[32] ),
    .A2(_07136_),
    .B1_N(_07137_),
    .X(_01254_));
 sky130_fd_sc_hd__a21oi_2 _22546_ (.A1(\csr._minstret_T_3[32] ),
    .A2(_07136_),
    .B1(\csr._minstret_T_3[33] ),
    .Y(_07138_));
 sky130_fd_sc_hd__and4_2 _22547_ (.A(\csr._minstret_T_3[33] ),
    .B(\csr._minstret_T_3[32] ),
    .C(\csr.minstret[31] ),
    .D(_06420_),
    .X(_07139_));
 sky130_fd_sc_hd__nor3_2 _22548_ (.A(_06377_),
    .B(_07138_),
    .C(_07139_),
    .Y(_01255_));
 sky130_fd_sc_hd__and4_2 _22549_ (.A(\csr._minstret_T_3[33] ),
    .B(\csr._minstret_T_3[32] ),
    .C(\csr.minstret[30] ),
    .D(\csr.minstret[31] ),
    .X(_07140_));
 sky130_fd_sc_hd__a31o_2 _22550_ (.A1(\csr._minstret_T_3[34] ),
    .A2(_06417_),
    .A3(_07140_),
    .B1(_06422_),
    .X(_07141_));
 sky130_fd_sc_hd__o21ba_2 _22551_ (.A1(\csr._minstret_T_3[34] ),
    .A2(_07139_),
    .B1_N(_07141_),
    .X(_01256_));
 sky130_fd_sc_hd__a21oi_2 _22552_ (.A1(\csr._minstret_T_3[34] ),
    .A2(_07139_),
    .B1(\csr._minstret_T_3[35] ),
    .Y(_07142_));
 sky130_fd_sc_hd__and3_2 _22553_ (.A(\csr._minstret_T_3[35] ),
    .B(\csr._minstret_T_3[34] ),
    .C(_07139_),
    .X(_07143_));
 sky130_fd_sc_hd__buf_1 _22554_ (.A(_07143_),
    .X(_07144_));
 sky130_fd_sc_hd__nor3_2 _22555_ (.A(_06377_),
    .B(_07142_),
    .C(_07144_),
    .Y(_01257_));
 sky130_fd_sc_hd__a21oi_2 _22556_ (.A1(\csr._minstret_T_3[36] ),
    .A2(_07144_),
    .B1(_06336_),
    .Y(_07145_));
 sky130_fd_sc_hd__o21a_2 _22557_ (.A1(\csr._minstret_T_3[36] ),
    .A2(_07144_),
    .B1(_07145_),
    .X(_01258_));
 sky130_fd_sc_hd__a21oi_2 _22558_ (.A1(\csr._minstret_T_3[36] ),
    .A2(_07144_),
    .B1(\csr._minstret_T_3[37] ),
    .Y(_07146_));
 sky130_fd_sc_hd__a311oi_2 _22559_ (.A1(\csr._minstret_T_3[37] ),
    .A2(\csr._minstret_T_3[36] ),
    .A3(_07144_),
    .B1(_07146_),
    .C1(_06336_),
    .Y(_01259_));
 sky130_fd_sc_hd__and3_2 _22560_ (.A(\csr._minstret_T_3[37] ),
    .B(\csr._minstret_T_3[36] ),
    .C(_07144_),
    .X(_07147_));
 sky130_fd_sc_hd__buf_1 _22561_ (.A(_10576_),
    .X(_07148_));
 sky130_fd_sc_hd__a41o_2 _22562_ (.A1(\csr._minstret_T_3[38] ),
    .A2(\csr._minstret_T_3[37] ),
    .A3(\csr._minstret_T_3[36] ),
    .A4(_07144_),
    .B1(_07148_),
    .X(_07149_));
 sky130_fd_sc_hd__o21ba_2 _22563_ (.A1(\csr._minstret_T_3[38] ),
    .A2(_07147_),
    .B1_N(_07149_),
    .X(_01260_));
 sky130_fd_sc_hd__a21oi_2 _22564_ (.A1(\csr._minstret_T_3[38] ),
    .A2(_07147_),
    .B1(\csr._minstret_T_3[39] ),
    .Y(_07150_));
 sky130_fd_sc_hd__and3_2 _22565_ (.A(\csr._minstret_T_3[39] ),
    .B(\csr._minstret_T_3[35] ),
    .C(\csr._minstret_T_3[34] ),
    .X(_07151_));
 sky130_fd_sc_hd__and4_2 _22566_ (.A(\csr._minstret_T_3[38] ),
    .B(\csr._minstret_T_3[37] ),
    .C(\csr._minstret_T_3[36] ),
    .D(_07151_),
    .X(_07152_));
 sky130_fd_sc_hd__and3_2 _22567_ (.A(_06417_),
    .B(_07140_),
    .C(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__nor3_2 _22568_ (.A(_06377_),
    .B(_07150_),
    .C(_07153_),
    .Y(_01261_));
 sky130_fd_sc_hd__a21oi_2 _22569_ (.A1(\csr._minstret_T_3[40] ),
    .A2(_07153_),
    .B1(_06336_),
    .Y(_07154_));
 sky130_fd_sc_hd__o21a_2 _22570_ (.A1(\csr._minstret_T_3[40] ),
    .A2(_07153_),
    .B1(_07154_),
    .X(_01262_));
 sky130_fd_sc_hd__inv_2 _22571_ (.A(\csr.minstret[27] ),
    .Y(_07155_));
 sky130_fd_sc_hd__nor2_2 _22572_ (.A(_07155_),
    .B(_06399_),
    .Y(_07156_));
 sky130_fd_sc_hd__and3_2 _22573_ (.A(\csr.minstret[28] ),
    .B(\csr.minstret[29] ),
    .C(_07156_),
    .X(_07157_));
 sky130_fd_sc_hd__and4_2 _22574_ (.A(\csr._minstret_T_3[33] ),
    .B(\csr.minstret[30] ),
    .C(\csr.minstret[31] ),
    .D(_07151_),
    .X(_07158_));
 sky130_fd_sc_hd__and4_2 _22575_ (.A(\csr._minstret_T_3[38] ),
    .B(\csr._minstret_T_3[37] ),
    .C(\csr._minstret_T_3[36] ),
    .D(_07158_),
    .X(_07159_));
 sky130_fd_sc_hd__and4_2 _22576_ (.A(\csr._minstret_T_3[40] ),
    .B(\csr._minstret_T_3[32] ),
    .C(_07157_),
    .D(_07159_),
    .X(_07160_));
 sky130_fd_sc_hd__and4_2 _22577_ (.A(\csr._minstret_T_3[33] ),
    .B(\csr._minstret_T_3[32] ),
    .C(\csr.minstret[31] ),
    .D(_07152_),
    .X(_07161_));
 sky130_fd_sc_hd__and3_2 _22578_ (.A(\csr._minstret_T_3[40] ),
    .B(_06420_),
    .C(_07161_),
    .X(_07162_));
 sky130_fd_sc_hd__nand2_2 _22579_ (.A(\csr._minstret_T_3[41] ),
    .B(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__buf_1 _22580_ (.A(_06578_),
    .X(_07164_));
 sky130_fd_sc_hd__o211a_2 _22581_ (.A1(\csr._minstret_T_3[41] ),
    .A2(_07160_),
    .B1(_07163_),
    .C1(_07164_),
    .X(_01263_));
 sky130_fd_sc_hd__a21oi_2 _22582_ (.A1(\csr._minstret_T_3[41] ),
    .A2(_07160_),
    .B1(\csr._minstret_T_3[42] ),
    .Y(_07165_));
 sky130_fd_sc_hd__and3_2 _22583_ (.A(\csr._minstret_T_3[42] ),
    .B(\csr._minstret_T_3[41] ),
    .C(_07162_),
    .X(_07166_));
 sky130_fd_sc_hd__nor3_2 _22584_ (.A(_06377_),
    .B(_07165_),
    .C(_07166_),
    .Y(_01264_));
 sky130_fd_sc_hd__a41o_2 _22585_ (.A1(\csr._minstret_T_3[43] ),
    .A2(\csr._minstret_T_3[42] ),
    .A3(\csr._minstret_T_3[41] ),
    .A4(_07162_),
    .B1(_07148_),
    .X(_07167_));
 sky130_fd_sc_hd__o21ba_2 _22586_ (.A1(\csr._minstret_T_3[43] ),
    .A2(_07166_),
    .B1_N(_07167_),
    .X(_01265_));
 sky130_fd_sc_hd__and4_2 _22587_ (.A(\csr._minstret_T_3[43] ),
    .B(\csr._minstret_T_3[42] ),
    .C(\csr._minstret_T_3[41] ),
    .D(_07160_),
    .X(_07168_));
 sky130_fd_sc_hd__a31o_2 _22588_ (.A1(\csr._minstret_T_3[44] ),
    .A2(\csr._minstret_T_3[43] ),
    .A3(_07166_),
    .B1(_06422_),
    .X(_07169_));
 sky130_fd_sc_hd__o21ba_2 _22589_ (.A1(\csr._minstret_T_3[44] ),
    .A2(_07168_),
    .B1_N(_07169_),
    .X(_01266_));
 sky130_fd_sc_hd__and3_2 _22590_ (.A(\csr._minstret_T_3[44] ),
    .B(\csr._minstret_T_3[43] ),
    .C(_07166_),
    .X(_07170_));
 sky130_fd_sc_hd__a41o_2 _22591_ (.A1(\csr._minstret_T_3[45] ),
    .A2(\csr._minstret_T_3[44] ),
    .A3(\csr._minstret_T_3[43] ),
    .A4(_07166_),
    .B1(_07148_),
    .X(_07171_));
 sky130_fd_sc_hd__o21ba_2 _22592_ (.A1(\csr._minstret_T_3[45] ),
    .A2(_07170_),
    .B1_N(_07171_),
    .X(_01267_));
 sky130_fd_sc_hd__and4_2 _22593_ (.A(\csr._minstret_T_3[45] ),
    .B(\csr._minstret_T_3[44] ),
    .C(\csr._minstret_T_3[43] ),
    .D(_07166_),
    .X(_07172_));
 sky130_fd_sc_hd__a31o_2 _22594_ (.A1(\csr._minstret_T_3[46] ),
    .A2(\csr._minstret_T_3[45] ),
    .A3(_07170_),
    .B1(_06422_),
    .X(_07173_));
 sky130_fd_sc_hd__o21ba_2 _22595_ (.A1(\csr._minstret_T_3[46] ),
    .A2(_07172_),
    .B1_N(_07173_),
    .X(_01268_));
 sky130_fd_sc_hd__and4_2 _22596_ (.A(\csr._minstret_T_3[46] ),
    .B(\csr._minstret_T_3[45] ),
    .C(\csr._minstret_T_3[44] ),
    .D(_07168_),
    .X(_07174_));
 sky130_fd_sc_hd__a31o_2 _22597_ (.A1(\csr._minstret_T_3[47] ),
    .A2(\csr._minstret_T_3[46] ),
    .A3(_07172_),
    .B1(_06422_),
    .X(_07175_));
 sky130_fd_sc_hd__o21ba_2 _22598_ (.A1(\csr._minstret_T_3[47] ),
    .A2(_07174_),
    .B1_N(_07175_),
    .X(_01269_));
 sky130_fd_sc_hd__a21oi_2 _22599_ (.A1(\csr._minstret_T_3[47] ),
    .A2(_07174_),
    .B1(\csr._minstret_T_3[48] ),
    .Y(_07176_));
 sky130_fd_sc_hd__and4_2 _22600_ (.A(\csr._minstret_T_3[48] ),
    .B(\csr._minstret_T_3[47] ),
    .C(\csr._minstret_T_3[46] ),
    .D(_07172_),
    .X(_07177_));
 sky130_fd_sc_hd__buf_1 _22601_ (.A(_07177_),
    .X(_07178_));
 sky130_fd_sc_hd__nor3_2 _22602_ (.A(_06377_),
    .B(_07176_),
    .C(_07178_),
    .Y(_01270_));
 sky130_fd_sc_hd__buf_1 _22603_ (.A(_10576_),
    .X(_07179_));
 sky130_fd_sc_hd__a21oi_2 _22604_ (.A1(\csr._minstret_T_3[49] ),
    .A2(_07178_),
    .B1(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__o21a_2 _22605_ (.A1(\csr._minstret_T_3[49] ),
    .A2(_07178_),
    .B1(_07180_),
    .X(_01271_));
 sky130_fd_sc_hd__and4_2 _22606_ (.A(\csr._minstret_T_3[49] ),
    .B(\csr._minstret_T_3[48] ),
    .C(\csr._minstret_T_3[47] ),
    .D(_07174_),
    .X(_07181_));
 sky130_fd_sc_hd__a31o_2 _22607_ (.A1(\csr._minstret_T_3[50] ),
    .A2(\csr._minstret_T_3[49] ),
    .A3(_07178_),
    .B1(_06422_),
    .X(_07182_));
 sky130_fd_sc_hd__o21ba_2 _22608_ (.A1(\csr._minstret_T_3[50] ),
    .A2(_07181_),
    .B1_N(_07182_),
    .X(_01272_));
 sky130_fd_sc_hd__a31oi_2 _22609_ (.A1(\csr._minstret_T_3[50] ),
    .A2(\csr._minstret_T_3[49] ),
    .A3(_07178_),
    .B1(\csr._minstret_T_3[51] ),
    .Y(_07183_));
 sky130_fd_sc_hd__and4_2 _22610_ (.A(\csr._minstret_T_3[51] ),
    .B(\csr._minstret_T_3[50] ),
    .C(\csr._minstret_T_3[49] ),
    .D(_07178_),
    .X(_07184_));
 sky130_fd_sc_hd__buf_1 _22611_ (.A(_07184_),
    .X(_07185_));
 sky130_fd_sc_hd__nor3_2 _22612_ (.A(_06377_),
    .B(_07183_),
    .C(_07185_),
    .Y(_01273_));
 sky130_fd_sc_hd__a21oi_2 _22613_ (.A1(\csr._minstret_T_3[52] ),
    .A2(_07185_),
    .B1(_07179_),
    .Y(_07186_));
 sky130_fd_sc_hd__o21a_2 _22614_ (.A1(\csr._minstret_T_3[52] ),
    .A2(_07185_),
    .B1(_07186_),
    .X(_01274_));
 sky130_fd_sc_hd__a21oi_2 _22615_ (.A1(\csr._minstret_T_3[52] ),
    .A2(_07185_),
    .B1(\csr._minstret_T_3[53] ),
    .Y(_07187_));
 sky130_fd_sc_hd__a311oi_2 _22616_ (.A1(\csr._minstret_T_3[53] ),
    .A2(\csr._minstret_T_3[52] ),
    .A3(_07185_),
    .B1(_07187_),
    .C1(_06336_),
    .Y(_01275_));
 sky130_fd_sc_hd__a31oi_2 _22617_ (.A1(\csr._minstret_T_3[53] ),
    .A2(\csr._minstret_T_3[52] ),
    .A3(_07185_),
    .B1(\csr._minstret_T_3[54] ),
    .Y(_07188_));
 sky130_fd_sc_hd__and4_2 _22618_ (.A(\csr._minstret_T_3[54] ),
    .B(\csr._minstret_T_3[53] ),
    .C(\csr._minstret_T_3[52] ),
    .D(_07185_),
    .X(_07189_));
 sky130_fd_sc_hd__buf_1 _22619_ (.A(_07189_),
    .X(_07190_));
 sky130_fd_sc_hd__nor3_2 _22620_ (.A(_06377_),
    .B(_07188_),
    .C(_07190_),
    .Y(_01276_));
 sky130_fd_sc_hd__a21oi_2 _22621_ (.A1(\csr._minstret_T_3[55] ),
    .A2(_07190_),
    .B1(_07179_),
    .Y(_07191_));
 sky130_fd_sc_hd__o21a_2 _22622_ (.A1(\csr._minstret_T_3[55] ),
    .A2(_07190_),
    .B1(_07191_),
    .X(_01277_));
 sky130_fd_sc_hd__a21oi_2 _22623_ (.A1(\csr._minstret_T_3[55] ),
    .A2(_07190_),
    .B1(\csr._minstret_T_3[56] ),
    .Y(_07192_));
 sky130_fd_sc_hd__a31o_2 _22624_ (.A1(\csr._minstret_T_3[56] ),
    .A2(\csr._minstret_T_3[55] ),
    .A3(_07190_),
    .B1(_07148_),
    .X(_07193_));
 sky130_fd_sc_hd__nor2_2 _22625_ (.A(_07192_),
    .B(_07193_),
    .Y(_01278_));
 sky130_fd_sc_hd__a31oi_2 _22626_ (.A1(\csr._minstret_T_3[56] ),
    .A2(\csr._minstret_T_3[55] ),
    .A3(_07190_),
    .B1(\csr._minstret_T_3[57] ),
    .Y(_07194_));
 sky130_fd_sc_hd__and4_2 _22627_ (.A(\csr._minstret_T_3[57] ),
    .B(\csr._minstret_T_3[56] ),
    .C(\csr._minstret_T_3[55] ),
    .D(_07190_),
    .X(_07195_));
 sky130_fd_sc_hd__buf_1 _22628_ (.A(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__nor3_2 _22629_ (.A(_06377_),
    .B(_07194_),
    .C(_07196_),
    .Y(_01279_));
 sky130_fd_sc_hd__a21oi_2 _22630_ (.A1(\csr._minstret_T_3[58] ),
    .A2(_07196_),
    .B1(_07179_),
    .Y(_07197_));
 sky130_fd_sc_hd__o21a_2 _22631_ (.A1(\csr._minstret_T_3[58] ),
    .A2(_07196_),
    .B1(_07197_),
    .X(_01280_));
 sky130_fd_sc_hd__a21oi_2 _22632_ (.A1(\csr._minstret_T_3[58] ),
    .A2(_07196_),
    .B1(\csr._minstret_T_3[59] ),
    .Y(_07198_));
 sky130_fd_sc_hd__a311oi_2 _22633_ (.A1(\csr._minstret_T_3[59] ),
    .A2(\csr._minstret_T_3[58] ),
    .A3(_07196_),
    .B1(_07198_),
    .C1(_06336_),
    .Y(_01281_));
 sky130_fd_sc_hd__buf_1 _22634_ (.A(_03579_),
    .X(_07199_));
 sky130_fd_sc_hd__a31oi_2 _22635_ (.A1(\csr._minstret_T_3[59] ),
    .A2(\csr._minstret_T_3[58] ),
    .A3(_07196_),
    .B1(\csr._minstret_T_3[60] ),
    .Y(_07200_));
 sky130_fd_sc_hd__and4_2 _22636_ (.A(\csr._minstret_T_3[60] ),
    .B(\csr._minstret_T_3[59] ),
    .C(\csr._minstret_T_3[58] ),
    .D(_07196_),
    .X(_07201_));
 sky130_fd_sc_hd__buf_1 _22637_ (.A(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__nor3_2 _22638_ (.A(_07199_),
    .B(_07200_),
    .C(_07202_),
    .Y(_01282_));
 sky130_fd_sc_hd__a21oi_2 _22639_ (.A1(\csr._minstret_T_3[61] ),
    .A2(_07202_),
    .B1(_07179_),
    .Y(_07203_));
 sky130_fd_sc_hd__o21a_2 _22640_ (.A1(\csr._minstret_T_3[61] ),
    .A2(_07202_),
    .B1(_07203_),
    .X(_01283_));
 sky130_fd_sc_hd__a21oi_2 _22641_ (.A1(\csr._minstret_T_3[61] ),
    .A2(_07202_),
    .B1(\csr._minstret_T_3[62] ),
    .Y(_07204_));
 sky130_fd_sc_hd__and3_2 _22642_ (.A(\csr._minstret_T_3[62] ),
    .B(\csr._minstret_T_3[61] ),
    .C(_07202_),
    .X(_07205_));
 sky130_fd_sc_hd__nor3_2 _22643_ (.A(_07199_),
    .B(_07204_),
    .C(_07205_),
    .Y(_01284_));
 sky130_fd_sc_hd__a41o_2 _22644_ (.A1(\csr._minstret_T_3[63] ),
    .A2(\csr._minstret_T_3[62] ),
    .A3(\csr._minstret_T_3[61] ),
    .A4(_07202_),
    .B1(_07148_),
    .X(_07206_));
 sky130_fd_sc_hd__o21ba_2 _22645_ (.A1(\csr._minstret_T_3[63] ),
    .A2(_07205_),
    .B1_N(_07206_),
    .X(_01285_));
 sky130_fd_sc_hd__and4_2 _22646_ (.A(_06457_),
    .B(_06313_),
    .C(_06458_),
    .D(_06466_),
    .X(_07207_));
 sky130_fd_sc_hd__buf_1 _22647_ (.A(_07207_),
    .X(_07208_));
 sky130_fd_sc_hd__nand4_2 _22648_ (.A(_06457_),
    .B(_06313_),
    .C(_06458_),
    .D(_06466_),
    .Y(_07209_));
 sky130_fd_sc_hd__buf_1 _22649_ (.A(_07209_),
    .X(_07210_));
 sky130_fd_sc_hd__or2_2 _22650_ (.A(\csr._mcycle_T_2[2] ),
    .B(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__o211a_2 _22651_ (.A1(\csr._csr_read_data_T_8[2] ),
    .A2(_07208_),
    .B1(_07211_),
    .C1(_07164_),
    .X(_01286_));
 sky130_fd_sc_hd__or2_2 _22652_ (.A(\csr._mcycle_T_2[3] ),
    .B(_07210_),
    .X(_07212_));
 sky130_fd_sc_hd__o211a_2 _22653_ (.A1(\csr._csr_read_data_T_8[3] ),
    .A2(_07208_),
    .B1(_07212_),
    .C1(_07164_),
    .X(_01287_));
 sky130_fd_sc_hd__or2_2 _22654_ (.A(\csr._mcycle_T_2[4] ),
    .B(_07210_),
    .X(_07213_));
 sky130_fd_sc_hd__o211a_2 _22655_ (.A1(\csr._csr_read_data_T_8[4] ),
    .A2(_07208_),
    .B1(_07213_),
    .C1(_07164_),
    .X(_01288_));
 sky130_fd_sc_hd__or2_2 _22656_ (.A(\csr._mcycle_T_2[5] ),
    .B(_07210_),
    .X(_07214_));
 sky130_fd_sc_hd__o211a_2 _22657_ (.A1(\csr._csr_read_data_T_8[5] ),
    .A2(_07208_),
    .B1(_07214_),
    .C1(_07164_),
    .X(_01289_));
 sky130_fd_sc_hd__or2_2 _22658_ (.A(\csr._mcycle_T_2[6] ),
    .B(_07210_),
    .X(_07215_));
 sky130_fd_sc_hd__o211a_2 _22659_ (.A1(\csr._csr_read_data_T_8[6] ),
    .A2(_07208_),
    .B1(_07215_),
    .C1(_07164_),
    .X(_01290_));
 sky130_fd_sc_hd__or2_2 _22660_ (.A(\csr._mcycle_T_2[7] ),
    .B(_07210_),
    .X(_07216_));
 sky130_fd_sc_hd__o211a_2 _22661_ (.A1(\csr._csr_read_data_T_8[7] ),
    .A2(_07208_),
    .B1(_07216_),
    .C1(_07164_),
    .X(_01291_));
 sky130_fd_sc_hd__or2_2 _22662_ (.A(\csr._mcycle_T_2[8] ),
    .B(_07210_),
    .X(_07217_));
 sky130_fd_sc_hd__o211a_2 _22663_ (.A1(\csr._csr_read_data_T_8[8] ),
    .A2(_07208_),
    .B1(_07217_),
    .C1(_07164_),
    .X(_01292_));
 sky130_fd_sc_hd__or2_2 _22664_ (.A(\csr._mcycle_T_2[9] ),
    .B(_07210_),
    .X(_07218_));
 sky130_fd_sc_hd__o211a_2 _22665_ (.A1(\csr._csr_read_data_T_8[9] ),
    .A2(_07208_),
    .B1(_07218_),
    .C1(_07164_),
    .X(_01293_));
 sky130_fd_sc_hd__or2_2 _22666_ (.A(\csr._mcycle_T_2[10] ),
    .B(_07210_),
    .X(_07219_));
 sky130_fd_sc_hd__o211a_2 _22667_ (.A1(\csr._csr_read_data_T_8[10] ),
    .A2(_07208_),
    .B1(_07219_),
    .C1(_07164_),
    .X(_01294_));
 sky130_fd_sc_hd__or2_2 _22668_ (.A(\csr._mcycle_T_2[11] ),
    .B(_07210_),
    .X(_07220_));
 sky130_fd_sc_hd__buf_1 _22669_ (.A(_06578_),
    .X(_07221_));
 sky130_fd_sc_hd__o211a_2 _22670_ (.A1(\csr._csr_read_data_T_8[11] ),
    .A2(_07208_),
    .B1(_07220_),
    .C1(_07221_),
    .X(_01295_));
 sky130_fd_sc_hd__buf_1 _22671_ (.A(_07207_),
    .X(_07222_));
 sky130_fd_sc_hd__buf_1 _22672_ (.A(_07209_),
    .X(_07223_));
 sky130_fd_sc_hd__or2_2 _22673_ (.A(\csr._mcycle_T_2[12] ),
    .B(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__o211a_2 _22674_ (.A1(\csr._csr_read_data_T_8[12] ),
    .A2(_07222_),
    .B1(_07224_),
    .C1(_07221_),
    .X(_01296_));
 sky130_fd_sc_hd__or2_2 _22675_ (.A(\csr._mcycle_T_2[13] ),
    .B(_07223_),
    .X(_07225_));
 sky130_fd_sc_hd__o211a_2 _22676_ (.A1(\csr._csr_read_data_T_8[13] ),
    .A2(_07222_),
    .B1(_07225_),
    .C1(_07221_),
    .X(_01297_));
 sky130_fd_sc_hd__or2_2 _22677_ (.A(\csr._mcycle_T_2[14] ),
    .B(_07223_),
    .X(_07226_));
 sky130_fd_sc_hd__o211a_2 _22678_ (.A1(\csr._csr_read_data_T_8[14] ),
    .A2(_07222_),
    .B1(_07226_),
    .C1(_07221_),
    .X(_01298_));
 sky130_fd_sc_hd__or2_2 _22679_ (.A(\csr._mcycle_T_2[15] ),
    .B(_07223_),
    .X(_07227_));
 sky130_fd_sc_hd__o211a_2 _22680_ (.A1(\csr._csr_read_data_T_8[15] ),
    .A2(_07222_),
    .B1(_07227_),
    .C1(_07221_),
    .X(_01299_));
 sky130_fd_sc_hd__or2_2 _22681_ (.A(\csr._mcycle_T_2[16] ),
    .B(_07223_),
    .X(_07228_));
 sky130_fd_sc_hd__o211a_2 _22682_ (.A1(\csr._csr_read_data_T_8[16] ),
    .A2(_07222_),
    .B1(_07228_),
    .C1(_07221_),
    .X(_01300_));
 sky130_fd_sc_hd__or2_2 _22683_ (.A(\csr._mcycle_T_2[17] ),
    .B(_07223_),
    .X(_07229_));
 sky130_fd_sc_hd__o211a_2 _22684_ (.A1(\csr._csr_read_data_T_8[17] ),
    .A2(_07222_),
    .B1(_07229_),
    .C1(_07221_),
    .X(_01301_));
 sky130_fd_sc_hd__or2_2 _22685_ (.A(\csr._mcycle_T_2[18] ),
    .B(_07223_),
    .X(_07230_));
 sky130_fd_sc_hd__o211a_2 _22686_ (.A1(\csr._csr_read_data_T_8[18] ),
    .A2(_07222_),
    .B1(_07230_),
    .C1(_07221_),
    .X(_01302_));
 sky130_fd_sc_hd__or2_2 _22687_ (.A(\csr._mcycle_T_2[19] ),
    .B(_07223_),
    .X(_07231_));
 sky130_fd_sc_hd__o211a_2 _22688_ (.A1(\csr._csr_read_data_T_8[19] ),
    .A2(_07222_),
    .B1(_07231_),
    .C1(_07221_),
    .X(_01303_));
 sky130_fd_sc_hd__or2_2 _22689_ (.A(\csr._mcycle_T_2[20] ),
    .B(_07223_),
    .X(_07232_));
 sky130_fd_sc_hd__o211a_2 _22690_ (.A1(\csr._csr_read_data_T_8[20] ),
    .A2(_07222_),
    .B1(_07232_),
    .C1(_07221_),
    .X(_01304_));
 sky130_fd_sc_hd__or2_2 _22691_ (.A(\csr._mcycle_T_2[21] ),
    .B(_07223_),
    .X(_07233_));
 sky130_fd_sc_hd__buf_1 _22692_ (.A(_06578_),
    .X(_07234_));
 sky130_fd_sc_hd__o211a_2 _22693_ (.A1(\csr._csr_read_data_T_8[21] ),
    .A2(_07222_),
    .B1(_07233_),
    .C1(_07234_),
    .X(_01305_));
 sky130_fd_sc_hd__buf_1 _22694_ (.A(_07207_),
    .X(_07235_));
 sky130_fd_sc_hd__buf_1 _22695_ (.A(_07209_),
    .X(_07236_));
 sky130_fd_sc_hd__or2_2 _22696_ (.A(\csr._mcycle_T_2[22] ),
    .B(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__o211a_2 _22697_ (.A1(\csr._csr_read_data_T_8[22] ),
    .A2(_07235_),
    .B1(_07237_),
    .C1(_07234_),
    .X(_01306_));
 sky130_fd_sc_hd__or2_2 _22698_ (.A(\csr._mcycle_T_2[23] ),
    .B(_07236_),
    .X(_07238_));
 sky130_fd_sc_hd__o211a_2 _22699_ (.A1(\csr._csr_read_data_T_8[23] ),
    .A2(_07235_),
    .B1(_07238_),
    .C1(_07234_),
    .X(_01307_));
 sky130_fd_sc_hd__or2_2 _22700_ (.A(\csr._mcycle_T_2[24] ),
    .B(_07236_),
    .X(_07239_));
 sky130_fd_sc_hd__o211a_2 _22701_ (.A1(\csr._csr_read_data_T_8[24] ),
    .A2(_07235_),
    .B1(_07239_),
    .C1(_07234_),
    .X(_01308_));
 sky130_fd_sc_hd__or2_2 _22702_ (.A(\csr._mcycle_T_2[25] ),
    .B(_07236_),
    .X(_07240_));
 sky130_fd_sc_hd__o211a_2 _22703_ (.A1(\csr._csr_read_data_T_8[25] ),
    .A2(_07235_),
    .B1(_07240_),
    .C1(_07234_),
    .X(_01309_));
 sky130_fd_sc_hd__or2_2 _22704_ (.A(\csr._mcycle_T_2[26] ),
    .B(_07236_),
    .X(_07241_));
 sky130_fd_sc_hd__o211a_2 _22705_ (.A1(\csr._csr_read_data_T_8[26] ),
    .A2(_07235_),
    .B1(_07241_),
    .C1(_07234_),
    .X(_01310_));
 sky130_fd_sc_hd__or2_2 _22706_ (.A(\csr._mcycle_T_2[27] ),
    .B(_07236_),
    .X(_07242_));
 sky130_fd_sc_hd__o211a_2 _22707_ (.A1(\csr._csr_read_data_T_8[27] ),
    .A2(_07235_),
    .B1(_07242_),
    .C1(_07234_),
    .X(_01311_));
 sky130_fd_sc_hd__or2_2 _22708_ (.A(\csr._mcycle_T_2[28] ),
    .B(_07236_),
    .X(_07243_));
 sky130_fd_sc_hd__o211a_2 _22709_ (.A1(\csr._csr_read_data_T_8[28] ),
    .A2(_07235_),
    .B1(_07243_),
    .C1(_07234_),
    .X(_01312_));
 sky130_fd_sc_hd__or2_2 _22710_ (.A(\csr._mcycle_T_2[29] ),
    .B(_07236_),
    .X(_07244_));
 sky130_fd_sc_hd__o211a_2 _22711_ (.A1(\csr._csr_read_data_T_8[29] ),
    .A2(_07235_),
    .B1(_07244_),
    .C1(_07234_),
    .X(_01313_));
 sky130_fd_sc_hd__or2_2 _22712_ (.A(\csr._mcycle_T_2[30] ),
    .B(_07236_),
    .X(_07245_));
 sky130_fd_sc_hd__o211a_2 _22713_ (.A1(\csr._csr_read_data_T_8[30] ),
    .A2(_07235_),
    .B1(_07245_),
    .C1(_07234_),
    .X(_01314_));
 sky130_fd_sc_hd__or2_2 _22714_ (.A(\csr._mcycle_T_2[31] ),
    .B(_07236_),
    .X(_07246_));
 sky130_fd_sc_hd__buf_1 _22715_ (.A(_06578_),
    .X(_07247_));
 sky130_fd_sc_hd__o211a_2 _22716_ (.A1(\csr._csr_read_data_T_8[31] ),
    .A2(_07235_),
    .B1(_07246_),
    .C1(_07247_),
    .X(_01315_));
 sky130_fd_sc_hd__or4b_2 _22717_ (.A(_10575_),
    .B(_11000_),
    .C(_11006_),
    .D_N(_10586_),
    .X(_07248_));
 sky130_fd_sc_hd__nand2_2 _22718_ (.A(_10943_),
    .B(_10941_),
    .Y(_07249_));
 sky130_fd_sc_hd__and3b_2 _22719_ (.A_N(\decode.control.io_funct3[0] ),
    .B(_10943_),
    .C(\decode.control.io_funct3[2] ),
    .X(_07250_));
 sky130_fd_sc_hd__o311a_2 _22720_ (.A1(_03524_),
    .A2(_03539_),
    .A3(_07250_),
    .B1(_03458_),
    .C1(\decode.control.io_opcode[5] ),
    .X(_07251_));
 sky130_fd_sc_hd__a41o_2 _22721_ (.A1(_10946_),
    .A2(_10964_),
    .A3(_10952_),
    .A4(_07249_),
    .B1(_07251_),
    .X(_07252_));
 sky130_fd_sc_hd__o21ai_2 _22722_ (.A1(_10946_),
    .A2(_03520_),
    .B1(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__nor4_2 _22723_ (.A(_03546_),
    .B(_07248_),
    .C(_07253_),
    .D(_03551_),
    .Y(_01316_));
 sky130_fd_sc_hd__and3_2 _22724_ (.A(_10941_),
    .B(_03458_),
    .C(_03541_),
    .X(_07254_));
 sky130_fd_sc_hd__and4bb_2 _22725_ (.A_N(_10913_),
    .B_N(_07248_),
    .C(_07254_),
    .D(_10916_),
    .X(_07255_));
 sky130_fd_sc_hd__buf_1 _22726_ (.A(_07255_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_2 _22727_ (.A0(_06101_),
    .A1(\fetch.bht.bhtTable_tag[10][0] ),
    .S(_09903_),
    .X(_07256_));
 sky130_fd_sc_hd__buf_1 _22728_ (.A(_07256_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_2 _22729_ (.A0(_06103_),
    .A1(\fetch.bht.bhtTable_tag[10][1] ),
    .S(_09903_),
    .X(_07257_));
 sky130_fd_sc_hd__buf_1 _22730_ (.A(_07257_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_2 _22731_ (.A0(_06105_),
    .A1(\fetch.bht.bhtTable_tag[10][2] ),
    .S(_09903_),
    .X(_07258_));
 sky130_fd_sc_hd__buf_1 _22732_ (.A(_07258_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_2 _22733_ (.A0(_06107_),
    .A1(\fetch.bht.bhtTable_tag[10][3] ),
    .S(_09903_),
    .X(_07259_));
 sky130_fd_sc_hd__buf_1 _22734_ (.A(_07259_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_2 _22735_ (.A0(_06109_),
    .A1(\fetch.bht.bhtTable_tag[10][4] ),
    .S(_09903_),
    .X(_07260_));
 sky130_fd_sc_hd__buf_1 _22736_ (.A(_07260_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_2 _22737_ (.A0(_06111_),
    .A1(\fetch.bht.bhtTable_tag[10][5] ),
    .S(_09903_),
    .X(_07261_));
 sky130_fd_sc_hd__buf_1 _22738_ (.A(_07261_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_2 _22739_ (.A0(_06113_),
    .A1(\fetch.bht.bhtTable_tag[10][6] ),
    .S(_09903_),
    .X(_07262_));
 sky130_fd_sc_hd__buf_1 _22740_ (.A(_07262_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_2 _22741_ (.A0(_06115_),
    .A1(\fetch.bht.bhtTable_tag[10][7] ),
    .S(_09903_),
    .X(_07263_));
 sky130_fd_sc_hd__buf_1 _22742_ (.A(_07263_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_2 _22743_ (.A0(_06117_),
    .A1(\fetch.bht.bhtTable_tag[10][8] ),
    .S(_09903_),
    .X(_07264_));
 sky130_fd_sc_hd__buf_1 _22744_ (.A(_07264_),
    .X(_01326_));
 sky130_fd_sc_hd__buf_1 _22745_ (.A(_09901_),
    .X(_07265_));
 sky130_fd_sc_hd__mux2_2 _22746_ (.A0(_06119_),
    .A1(\fetch.bht.bhtTable_tag[10][9] ),
    .S(_07265_),
    .X(_07266_));
 sky130_fd_sc_hd__buf_1 _22747_ (.A(_07266_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_2 _22748_ (.A0(_06122_),
    .A1(\fetch.bht.bhtTable_tag[10][10] ),
    .S(_07265_),
    .X(_07267_));
 sky130_fd_sc_hd__buf_1 _22749_ (.A(_07267_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_2 _22750_ (.A0(_06124_),
    .A1(\fetch.bht.bhtTable_tag[10][11] ),
    .S(_07265_),
    .X(_07268_));
 sky130_fd_sc_hd__buf_1 _22751_ (.A(_07268_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_2 _22752_ (.A0(_06126_),
    .A1(\fetch.bht.bhtTable_tag[10][12] ),
    .S(_07265_),
    .X(_07269_));
 sky130_fd_sc_hd__buf_1 _22753_ (.A(_07269_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_2 _22754_ (.A0(_06128_),
    .A1(\fetch.bht.bhtTable_tag[10][13] ),
    .S(_07265_),
    .X(_07270_));
 sky130_fd_sc_hd__buf_1 _22755_ (.A(_07270_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_2 _22756_ (.A0(_06130_),
    .A1(\fetch.bht.bhtTable_tag[10][14] ),
    .S(_07265_),
    .X(_07271_));
 sky130_fd_sc_hd__buf_1 _22757_ (.A(_07271_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_2 _22758_ (.A0(_06132_),
    .A1(\fetch.bht.bhtTable_tag[10][15] ),
    .S(_07265_),
    .X(_07272_));
 sky130_fd_sc_hd__buf_1 _22759_ (.A(_07272_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_2 _22760_ (.A0(_06134_),
    .A1(\fetch.bht.bhtTable_tag[10][16] ),
    .S(_07265_),
    .X(_07273_));
 sky130_fd_sc_hd__buf_1 _22761_ (.A(_07273_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_2 _22762_ (.A0(_06136_),
    .A1(\fetch.bht.bhtTable_tag[10][17] ),
    .S(_07265_),
    .X(_07274_));
 sky130_fd_sc_hd__buf_1 _22763_ (.A(_07274_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_2 _22764_ (.A0(_06138_),
    .A1(\fetch.bht.bhtTable_tag[10][18] ),
    .S(_07265_),
    .X(_07275_));
 sky130_fd_sc_hd__buf_1 _22765_ (.A(_07275_),
    .X(_01336_));
 sky130_fd_sc_hd__buf_1 _22766_ (.A(_09901_),
    .X(_07276_));
 sky130_fd_sc_hd__mux2_2 _22767_ (.A0(_06140_),
    .A1(\fetch.bht.bhtTable_tag[10][19] ),
    .S(_07276_),
    .X(_07277_));
 sky130_fd_sc_hd__buf_1 _22768_ (.A(_07277_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_2 _22769_ (.A0(_06143_),
    .A1(\fetch.bht.bhtTable_tag[10][20] ),
    .S(_07276_),
    .X(_07278_));
 sky130_fd_sc_hd__buf_1 _22770_ (.A(_07278_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_2 _22771_ (.A0(_06145_),
    .A1(\fetch.bht.bhtTable_tag[10][21] ),
    .S(_07276_),
    .X(_07279_));
 sky130_fd_sc_hd__buf_1 _22772_ (.A(_07279_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_2 _22773_ (.A0(_06147_),
    .A1(\fetch.bht.bhtTable_tag[10][22] ),
    .S(_07276_),
    .X(_07280_));
 sky130_fd_sc_hd__buf_1 _22774_ (.A(_07280_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_2 _22775_ (.A0(_06149_),
    .A1(\fetch.bht.bhtTable_tag[10][23] ),
    .S(_07276_),
    .X(_07281_));
 sky130_fd_sc_hd__buf_1 _22776_ (.A(_07281_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_2 _22777_ (.A0(_06151_),
    .A1(\fetch.bht.bhtTable_tag[10][24] ),
    .S(_07276_),
    .X(_07282_));
 sky130_fd_sc_hd__buf_1 _22778_ (.A(_07282_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_2 _22779_ (.A0(_06153_),
    .A1(\fetch.bht.bhtTable_tag[10][25] ),
    .S(_07276_),
    .X(_07283_));
 sky130_fd_sc_hd__buf_1 _22780_ (.A(_07283_),
    .X(_01343_));
 sky130_fd_sc_hd__and4_2 _22781_ (.A(_09880_),
    .B(_09882_),
    .C(_09885_),
    .D(_09892_),
    .X(_07284_));
 sky130_fd_sc_hd__buf_1 _22782_ (.A(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__buf_1 _22783_ (.A(_07285_),
    .X(_07286_));
 sky130_fd_sc_hd__mux2_2 _22784_ (.A0(\fetch.bht.bhtTable_tag[12][0] ),
    .A1(_10820_),
    .S(_07286_),
    .X(_07287_));
 sky130_fd_sc_hd__buf_1 _22785_ (.A(_07287_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_2 _22786_ (.A0(\fetch.bht.bhtTable_tag[12][1] ),
    .A1(_10821_),
    .S(_07286_),
    .X(_07288_));
 sky130_fd_sc_hd__buf_1 _22787_ (.A(_07288_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_2 _22788_ (.A0(\fetch.bht.bhtTable_tag[12][2] ),
    .A1(_10881_),
    .S(_07286_),
    .X(_07289_));
 sky130_fd_sc_hd__buf_1 _22789_ (.A(_07289_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_2 _22790_ (.A0(\fetch.bht.bhtTable_tag[12][3] ),
    .A1(_10817_),
    .S(_07286_),
    .X(_07290_));
 sky130_fd_sc_hd__buf_1 _22791_ (.A(_07290_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_2 _22792_ (.A0(\fetch.bht.bhtTable_tag[12][4] ),
    .A1(_10878_),
    .S(_07286_),
    .X(_07291_));
 sky130_fd_sc_hd__buf_1 _22793_ (.A(_07291_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_2 _22794_ (.A0(\fetch.bht.bhtTable_tag[12][5] ),
    .A1(_10812_),
    .S(_07286_),
    .X(_07292_));
 sky130_fd_sc_hd__buf_1 _22795_ (.A(_07292_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_2 _22796_ (.A0(\fetch.bht.bhtTable_tag[12][6] ),
    .A1(\csr.io_mem_pc[12] ),
    .S(_07286_),
    .X(_07293_));
 sky130_fd_sc_hd__buf_1 _22797_ (.A(_07293_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_2 _22798_ (.A0(\fetch.bht.bhtTable_tag[12][7] ),
    .A1(_10871_),
    .S(_07286_),
    .X(_07294_));
 sky130_fd_sc_hd__buf_1 _22799_ (.A(_07294_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_2 _22800_ (.A0(\fetch.bht.bhtTable_tag[12][8] ),
    .A1(_10872_),
    .S(_07286_),
    .X(_07295_));
 sky130_fd_sc_hd__buf_1 _22801_ (.A(_07295_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_2 _22802_ (.A0(\fetch.bht.bhtTable_tag[12][9] ),
    .A1(_10807_),
    .S(_07286_),
    .X(_07296_));
 sky130_fd_sc_hd__buf_1 _22803_ (.A(_07296_),
    .X(_01353_));
 sky130_fd_sc_hd__buf_1 _22804_ (.A(_07285_),
    .X(_07297_));
 sky130_fd_sc_hd__mux2_2 _22805_ (.A0(\fetch.bht.bhtTable_tag[12][10] ),
    .A1(_10868_),
    .S(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__buf_1 _22806_ (.A(_07298_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_2 _22807_ (.A0(\fetch.bht.bhtTable_tag[12][11] ),
    .A1(_10803_),
    .S(_07297_),
    .X(_07299_));
 sky130_fd_sc_hd__buf_1 _22808_ (.A(_07299_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_2 _22809_ (.A0(\fetch.bht.bhtTable_tag[12][12] ),
    .A1(\csr.io_mem_pc[18] ),
    .S(_07297_),
    .X(_07300_));
 sky130_fd_sc_hd__buf_1 _22810_ (.A(_07300_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_2 _22811_ (.A0(\fetch.bht.bhtTable_tag[12][13] ),
    .A1(_10800_),
    .S(_07297_),
    .X(_07301_));
 sky130_fd_sc_hd__buf_1 _22812_ (.A(_07301_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_2 _22813_ (.A0(\fetch.bht.bhtTable_tag[12][14] ),
    .A1(_10795_),
    .S(_07297_),
    .X(_07302_));
 sky130_fd_sc_hd__buf_1 _22814_ (.A(_07302_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_2 _22815_ (.A0(\fetch.bht.bhtTable_tag[12][15] ),
    .A1(\csr.io_mem_pc[21] ),
    .S(_07297_),
    .X(_07303_));
 sky130_fd_sc_hd__buf_1 _22816_ (.A(_07303_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_2 _22817_ (.A0(\fetch.bht.bhtTable_tag[12][16] ),
    .A1(_10787_),
    .S(_07297_),
    .X(_07304_));
 sky130_fd_sc_hd__buf_1 _22818_ (.A(_07304_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_2 _22819_ (.A0(\fetch.bht.bhtTable_tag[12][17] ),
    .A1(\csr.io_mem_pc[23] ),
    .S(_07297_),
    .X(_07305_));
 sky130_fd_sc_hd__buf_1 _22820_ (.A(_07305_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_2 _22821_ (.A0(\fetch.bht.bhtTable_tag[12][18] ),
    .A1(_10772_),
    .S(_07297_),
    .X(_07306_));
 sky130_fd_sc_hd__buf_1 _22822_ (.A(_07306_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_2 _22823_ (.A0(\fetch.bht.bhtTable_tag[12][19] ),
    .A1(_10773_),
    .S(_07297_),
    .X(_07307_));
 sky130_fd_sc_hd__buf_1 _22824_ (.A(_07307_),
    .X(_01363_));
 sky130_fd_sc_hd__buf_1 _22825_ (.A(_07284_),
    .X(_07308_));
 sky130_fd_sc_hd__mux2_2 _22826_ (.A0(\fetch.bht.bhtTable_tag[12][20] ),
    .A1(_10760_),
    .S(_07308_),
    .X(_07309_));
 sky130_fd_sc_hd__buf_1 _22827_ (.A(_07309_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_2 _22828_ (.A0(\fetch.bht.bhtTable_tag[12][21] ),
    .A1(_10759_),
    .S(_07308_),
    .X(_07310_));
 sky130_fd_sc_hd__buf_1 _22829_ (.A(_07310_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_2 _22830_ (.A0(\fetch.bht.bhtTable_tag[12][22] ),
    .A1(_10771_),
    .S(_07308_),
    .X(_07311_));
 sky130_fd_sc_hd__buf_1 _22831_ (.A(_07311_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_2 _22832_ (.A0(\fetch.bht.bhtTable_tag[12][23] ),
    .A1(\csr.io_mem_pc[29] ),
    .S(_07308_),
    .X(_07312_));
 sky130_fd_sc_hd__buf_1 _22833_ (.A(_07312_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_2 _22834_ (.A0(\fetch.bht.bhtTable_tag[12][24] ),
    .A1(_10777_),
    .S(_07308_),
    .X(_07313_));
 sky130_fd_sc_hd__buf_1 _22835_ (.A(_07313_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_2 _22836_ (.A0(\fetch.bht.bhtTable_tag[12][25] ),
    .A1(\csr.io_mem_pc[31] ),
    .S(_07308_),
    .X(_07314_));
 sky130_fd_sc_hd__buf_1 _22837_ (.A(_07314_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_2 _22838_ (.A0(\fetch.bht.bhtTable_tag[11][0] ),
    .A1(_10820_),
    .S(_09898_),
    .X(_07315_));
 sky130_fd_sc_hd__buf_1 _22839_ (.A(_07315_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_2 _22840_ (.A0(\fetch.bht.bhtTable_tag[11][1] ),
    .A1(_10821_),
    .S(_09898_),
    .X(_07316_));
 sky130_fd_sc_hd__buf_1 _22841_ (.A(_07316_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_2 _22842_ (.A0(\fetch.bht.bhtTable_tag[11][2] ),
    .A1(_10881_),
    .S(_09898_),
    .X(_07317_));
 sky130_fd_sc_hd__buf_1 _22843_ (.A(_07317_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_2 _22844_ (.A0(\fetch.bht.bhtTable_tag[11][3] ),
    .A1(_10817_),
    .S(_09898_),
    .X(_07318_));
 sky130_fd_sc_hd__buf_1 _22845_ (.A(_07318_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_2 _22846_ (.A0(\fetch.bht.bhtTable_tag[11][4] ),
    .A1(_10878_),
    .S(_09898_),
    .X(_07319_));
 sky130_fd_sc_hd__buf_1 _22847_ (.A(_07319_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_2 _22848_ (.A0(\fetch.bht.bhtTable_tag[11][5] ),
    .A1(_10812_),
    .S(_09898_),
    .X(_07320_));
 sky130_fd_sc_hd__buf_1 _22849_ (.A(_07320_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_2 _22850_ (.A0(\fetch.bht.bhtTable_tag[11][6] ),
    .A1(\csr.io_mem_pc[12] ),
    .S(_09898_),
    .X(_07321_));
 sky130_fd_sc_hd__buf_1 _22851_ (.A(_07321_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_2 _22852_ (.A0(\fetch.bht.bhtTable_tag[11][7] ),
    .A1(_10871_),
    .S(_09898_),
    .X(_07322_));
 sky130_fd_sc_hd__buf_1 _22853_ (.A(_07322_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_2 _22854_ (.A0(\fetch.bht.bhtTable_tag[11][8] ),
    .A1(_10872_),
    .S(_09898_),
    .X(_07323_));
 sky130_fd_sc_hd__buf_1 _22855_ (.A(_07323_),
    .X(_01378_));
 sky130_fd_sc_hd__buf_1 _22856_ (.A(_09896_),
    .X(_07324_));
 sky130_fd_sc_hd__mux2_2 _22857_ (.A0(\fetch.bht.bhtTable_tag[11][9] ),
    .A1(_10807_),
    .S(_07324_),
    .X(_07325_));
 sky130_fd_sc_hd__buf_1 _22858_ (.A(_07325_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_2 _22859_ (.A0(\fetch.bht.bhtTable_tag[11][10] ),
    .A1(_10868_),
    .S(_07324_),
    .X(_07326_));
 sky130_fd_sc_hd__buf_1 _22860_ (.A(_07326_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_2 _22861_ (.A0(\fetch.bht.bhtTable_tag[11][11] ),
    .A1(_10803_),
    .S(_07324_),
    .X(_07327_));
 sky130_fd_sc_hd__buf_1 _22862_ (.A(_07327_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_2 _22863_ (.A0(\fetch.bht.bhtTable_tag[11][12] ),
    .A1(\csr.io_mem_pc[18] ),
    .S(_07324_),
    .X(_07328_));
 sky130_fd_sc_hd__buf_1 _22864_ (.A(_07328_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_2 _22865_ (.A0(\fetch.bht.bhtTable_tag[11][13] ),
    .A1(_10800_),
    .S(_07324_),
    .X(_07329_));
 sky130_fd_sc_hd__buf_1 _22866_ (.A(_07329_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_2 _22867_ (.A0(\fetch.bht.bhtTable_tag[11][14] ),
    .A1(_10795_),
    .S(_07324_),
    .X(_07330_));
 sky130_fd_sc_hd__buf_1 _22868_ (.A(_07330_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_2 _22869_ (.A0(\fetch.bht.bhtTable_tag[11][15] ),
    .A1(\csr.io_mem_pc[21] ),
    .S(_07324_),
    .X(_07331_));
 sky130_fd_sc_hd__buf_1 _22870_ (.A(_07331_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_2 _22871_ (.A0(\fetch.bht.bhtTable_tag[11][16] ),
    .A1(_10787_),
    .S(_07324_),
    .X(_07332_));
 sky130_fd_sc_hd__buf_1 _22872_ (.A(_07332_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_2 _22873_ (.A0(\fetch.bht.bhtTable_tag[11][17] ),
    .A1(\csr.io_mem_pc[23] ),
    .S(_07324_),
    .X(_07333_));
 sky130_fd_sc_hd__buf_1 _22874_ (.A(_07333_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_2 _22875_ (.A0(\fetch.bht.bhtTable_tag[11][18] ),
    .A1(_10772_),
    .S(_07324_),
    .X(_07334_));
 sky130_fd_sc_hd__buf_1 _22876_ (.A(_07334_),
    .X(_01388_));
 sky130_fd_sc_hd__buf_1 _22877_ (.A(_09896_),
    .X(_07335_));
 sky130_fd_sc_hd__mux2_2 _22878_ (.A0(\fetch.bht.bhtTable_tag[11][19] ),
    .A1(_10773_),
    .S(_07335_),
    .X(_07336_));
 sky130_fd_sc_hd__buf_1 _22879_ (.A(_07336_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_2 _22880_ (.A0(\fetch.bht.bhtTable_tag[11][20] ),
    .A1(_10760_),
    .S(_07335_),
    .X(_07337_));
 sky130_fd_sc_hd__buf_1 _22881_ (.A(_07337_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_2 _22882_ (.A0(\fetch.bht.bhtTable_tag[11][21] ),
    .A1(_10759_),
    .S(_07335_),
    .X(_07338_));
 sky130_fd_sc_hd__buf_1 _22883_ (.A(_07338_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_2 _22884_ (.A0(\fetch.bht.bhtTable_tag[11][22] ),
    .A1(_10771_),
    .S(_07335_),
    .X(_07339_));
 sky130_fd_sc_hd__buf_1 _22885_ (.A(_07339_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_2 _22886_ (.A0(\fetch.bht.bhtTable_tag[11][23] ),
    .A1(\csr.io_mem_pc[29] ),
    .S(_07335_),
    .X(_07340_));
 sky130_fd_sc_hd__buf_1 _22887_ (.A(_07340_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_2 _22888_ (.A0(\fetch.bht.bhtTable_tag[11][24] ),
    .A1(_10777_),
    .S(_07335_),
    .X(_07341_));
 sky130_fd_sc_hd__buf_1 _22889_ (.A(_07341_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_2 _22890_ (.A0(\fetch.bht.bhtTable_tag[11][25] ),
    .A1(\csr.io_mem_pc[31] ),
    .S(_07335_),
    .X(_07342_));
 sky130_fd_sc_hd__buf_1 _22891_ (.A(_07342_),
    .X(_01395_));
 sky130_fd_sc_hd__buf_1 _22892_ (.A(_06248_),
    .X(_07343_));
 sky130_fd_sc_hd__buf_1 _22893_ (.A(_03500_),
    .X(_07344_));
 sky130_fd_sc_hd__buf_1 _22894_ (.A(_03592_),
    .X(_07345_));
 sky130_fd_sc_hd__nor2_2 _22895_ (.A(_06032_),
    .B(_07345_),
    .Y(_07346_));
 sky130_fd_sc_hd__and3_2 _22896_ (.A(_03592_),
    .B(_10672_),
    .C(_03590_),
    .X(_07347_));
 sky130_fd_sc_hd__buf_1 _22897_ (.A(_07347_),
    .X(_07348_));
 sky130_fd_sc_hd__nand2_2 _22898_ (.A(_06820_),
    .B(_07037_),
    .Y(_07349_));
 sky130_fd_sc_hd__o2bb2a_2 _22899_ (.A1_N(io_fetch_address[9]),
    .A2_N(_06717_),
    .B1(_06698_),
    .B2(io_fetch_address[13]),
    .X(_07350_));
 sky130_fd_sc_hd__o2111ai_2 _22900_ (.A1(_06718_),
    .A2(_06717_),
    .B1(_07048_),
    .C1(_07058_),
    .D1(_07350_),
    .Y(_07351_));
 sky130_fd_sc_hd__or4bb_2 _22901_ (.A(_06976_),
    .B(_07351_),
    .C_N(_06956_),
    .D_N(_06964_),
    .X(_07352_));
 sky130_fd_sc_hd__or4b_2 _22902_ (.A(_06785_),
    .B(_07349_),
    .C(_07352_),
    .D_N(_07035_),
    .X(_07353_));
 sky130_fd_sc_hd__nor4_2 _22903_ (.A(_06944_),
    .B(_06928_),
    .C(_07018_),
    .D(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__a22oi_2 _22904_ (.A1(io_fetch_address[11]),
    .A2(_06794_),
    .B1(_06806_),
    .B2(io_fetch_address[30]),
    .Y(_07355_));
 sky130_fd_sc_hd__o221a_2 _22905_ (.A1(io_fetch_address[30]),
    .A2(_06806_),
    .B1(_06670_),
    .B2(io_fetch_address[24]),
    .C1(_07355_),
    .X(_07356_));
 sky130_fd_sc_hd__nand2_2 _22906_ (.A(_06656_),
    .B(_06795_),
    .Y(_07357_));
 sky130_fd_sc_hd__or2_2 _22907_ (.A(io_fetch_address[10]),
    .B(_06739_),
    .X(_07358_));
 sky130_fd_sc_hd__and4b_2 _22908_ (.A_N(_06671_),
    .B(_07356_),
    .C(_07357_),
    .D(_07358_),
    .X(_07359_));
 sky130_fd_sc_hd__a2bb2o_2 _22909_ (.A1_N(io_fetch_address[17]),
    .A2_N(_06886_),
    .B1(_06862_),
    .B2(io_fetch_address[23]),
    .X(_07360_));
 sky130_fd_sc_hd__a221oi_2 _22910_ (.A1(io_fetch_address[21]),
    .A2(_06833_),
    .B1(_06767_),
    .B2(io_fetch_address[19]),
    .C1(_06893_),
    .Y(_07361_));
 sky130_fd_sc_hd__or4b_2 _22911_ (.A(_06834_),
    .B(_07360_),
    .C(_06849_),
    .D_N(_07361_),
    .X(_07362_));
 sky130_fd_sc_hd__a2111oi_2 _22912_ (.A1(io_fetch_address[13]),
    .A2(_06698_),
    .B1(_06916_),
    .C1(_06894_),
    .D1(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__o22a_2 _22913_ (.A1(io_fetch_address[11]),
    .A2(_06794_),
    .B1(_06862_),
    .B2(io_fetch_address[23]),
    .X(_07364_));
 sky130_fd_sc_hd__and4bb_2 _22914_ (.A_N(_06888_),
    .B_N(_07007_),
    .C(_07363_),
    .D(_07364_),
    .X(_07365_));
 sky130_fd_sc_hd__and4_2 _22915_ (.A(_06768_),
    .B(_07359_),
    .C(_07365_),
    .D(_06896_),
    .X(_07366_));
 sky130_fd_sc_hd__and2_2 _22916_ (.A(_07354_),
    .B(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__buf_1 _22917_ (.A(_07367_),
    .X(_07368_));
 sky130_fd_sc_hd__mux4_2 _22918_ (.A0(\fetch.bht.bhtTable_target_pc[4][2] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][2] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][2] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][2] ),
    .S0(_07107_),
    .S1(_07071_),
    .X(_07369_));
 sky130_fd_sc_hd__mux4_2 _22919_ (.A0(\fetch.bht.bhtTable_target_pc[0][2] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][2] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][2] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][2] ),
    .S0(_07119_),
    .S1(_07071_),
    .X(_07370_));
 sky130_fd_sc_hd__buf_1 _22920_ (.A(_07080_),
    .X(_07371_));
 sky130_fd_sc_hd__mux2_2 _22921_ (.A0(_07369_),
    .A1(_07370_),
    .S(_07371_),
    .X(_07372_));
 sky130_fd_sc_hd__mux2_2 _22922_ (.A0(\fetch.bht.bhtTable_target_pc[12][2] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][2] ),
    .S(_07068_),
    .X(_07373_));
 sky130_fd_sc_hd__and2b_2 _22923_ (.A_N(_07103_),
    .B(_07373_),
    .X(_07374_));
 sky130_fd_sc_hd__mux2_2 _22924_ (.A0(\fetch.bht.bhtTable_target_pc[14][2] ),
    .A1(\fetch.bht.bhtTable_target_pc[15][2] ),
    .S(_07119_),
    .X(_07375_));
 sky130_fd_sc_hd__a21o_2 _22925_ (.A1(_07375_),
    .A2(_07101_),
    .B1(_07081_),
    .X(_07376_));
 sky130_fd_sc_hd__mux4_2 _22926_ (.A0(\fetch.bht.bhtTable_target_pc[8][2] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][2] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][2] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][2] ),
    .S0(_07107_),
    .S1(_07114_),
    .X(_07377_));
 sky130_fd_sc_hd__o221a_2 _22927_ (.A1(_07374_),
    .A2(_07376_),
    .B1(_07377_),
    .B2(_07122_),
    .C1(_06740_),
    .X(_07378_));
 sky130_fd_sc_hd__a21oi_2 _22928_ (.A1(_07372_),
    .A2(_07085_),
    .B1(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__and2_2 _22929_ (.A(_07130_),
    .B(io_fetch_address[2]),
    .X(_07380_));
 sky130_fd_sc_hd__a211oi_2 _22930_ (.A1(_07368_),
    .A2(_07379_),
    .B1(_05246_),
    .C1(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__a221o_2 _22931_ (.A1(\csr._csr_read_data_T_8[2] ),
    .A2(_06039_),
    .B1(\csr.io_mret_vector[2] ),
    .B2(_06463_),
    .C1(_07381_),
    .X(_07382_));
 sky130_fd_sc_hd__a211o_2 _22932_ (.A1(\execute.io_target_pc[2] ),
    .A2(_07346_),
    .B1(_07348_),
    .C1(_07382_),
    .X(_07383_));
 sky130_fd_sc_hd__o311a_2 _22933_ (.A1(io_fetch_address[2]),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07383_),
    .C1(_06566_),
    .X(_01396_));
 sky130_fd_sc_hd__buf_1 _22934_ (.A(_07066_),
    .X(_07384_));
 sky130_fd_sc_hd__mux4_2 _22935_ (.A0(\fetch.bht.bhtTable_target_pc[12][3] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][3] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][3] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][3] ),
    .S0(_07384_),
    .S1(_07113_),
    .X(_07385_));
 sky130_fd_sc_hd__buf_1 _22936_ (.A(_06661_),
    .X(_07386_));
 sky130_fd_sc_hd__mux4_2 _22937_ (.A0(\fetch.bht.bhtTable_target_pc[8][3] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][3] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][3] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][3] ),
    .S0(_07106_),
    .S1(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__mux4_2 _22938_ (.A0(\fetch.bht.bhtTable_target_pc[4][3] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][3] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][3] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][3] ),
    .S0(_07106_),
    .S1(_07386_),
    .X(_07388_));
 sky130_fd_sc_hd__mux4_2 _22939_ (.A0(\fetch.bht.bhtTable_target_pc[0][3] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][3] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][3] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][3] ),
    .S0(_07384_),
    .S1(_07113_),
    .X(_07389_));
 sky130_fd_sc_hd__mux4_2 _22940_ (.A0(_07385_),
    .A1(_07387_),
    .A2(_07388_),
    .A3(_07389_),
    .S0(_07080_),
    .S1(_06637_),
    .X(_07390_));
 sky130_fd_sc_hd__buf_1 _22941_ (.A(_07354_),
    .X(_07391_));
 sky130_fd_sc_hd__buf_1 _22942_ (.A(_07366_),
    .X(_07392_));
 sky130_fd_sc_hd__and2_2 _22943_ (.A(io_fetch_address[3]),
    .B(io_fetch_address[2]),
    .X(_07393_));
 sky130_fd_sc_hd__nor2_2 _22944_ (.A(io_fetch_address[3]),
    .B(io_fetch_address[2]),
    .Y(_07394_));
 sky130_fd_sc_hd__a211oi_2 _22945_ (.A1(_07391_),
    .A2(_07392_),
    .B1(_07393_),
    .C1(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__a211o_2 _22946_ (.A1(_07390_),
    .A2(_07367_),
    .B1(_07090_),
    .C1(_07395_),
    .X(_07396_));
 sky130_fd_sc_hd__o211a_2 _22947_ (.A1(\execute.io_target_pc[3] ),
    .A2(_03592_),
    .B1(_03590_),
    .C1(_07396_),
    .X(_07397_));
 sky130_fd_sc_hd__a221o_2 _22948_ (.A1(\csr._csr_read_data_T_8[3] ),
    .A2(_06481_),
    .B1(\csr.io_mret_vector[3] ),
    .B2(_06463_),
    .C1(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__o31a_2 _22949_ (.A1(_06032_),
    .A2(_07091_),
    .A3(_10915_),
    .B1(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__a211o_2 _22950_ (.A1(io_fetch_address[3]),
    .A2(_07348_),
    .B1(_07399_),
    .C1(_03580_),
    .X(_01397_));
 sky130_fd_sc_hd__a22o_2 _22951_ (.A1(\csr._csr_read_data_T_8[4] ),
    .A2(_06039_),
    .B1(\csr.io_mret_vector[4] ),
    .B2(_06463_),
    .X(_07400_));
 sky130_fd_sc_hd__mux4_2 _22952_ (.A0(\fetch.bht.bhtTable_target_pc[12][4] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][4] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][4] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][4] ),
    .S0(_07123_),
    .S1(_07101_),
    .X(_07401_));
 sky130_fd_sc_hd__mux4_2 _22953_ (.A0(\fetch.bht.bhtTable_target_pc[8][4] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][4] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][4] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][4] ),
    .S0(_07123_),
    .S1(_07101_),
    .X(_07402_));
 sky130_fd_sc_hd__mux2_2 _22954_ (.A0(_07401_),
    .A1(_07402_),
    .S(_07082_),
    .X(_07403_));
 sky130_fd_sc_hd__mux4_2 _22955_ (.A0(\fetch.bht.bhtTable_target_pc[0][4] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][4] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][4] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][4] ),
    .S0(_07108_),
    .S1(_07115_),
    .X(_07404_));
 sky130_fd_sc_hd__nor2_2 _22956_ (.A(_07076_),
    .B(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__buf_1 _22957_ (.A(_07371_),
    .X(_07406_));
 sky130_fd_sc_hd__buf_1 _22958_ (.A(_07119_),
    .X(_07407_));
 sky130_fd_sc_hd__mux4_2 _22959_ (.A0(\fetch.bht.bhtTable_target_pc[4][4] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][4] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][4] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][4] ),
    .S0(_07407_),
    .S1(_07115_),
    .X(_07408_));
 sky130_fd_sc_hd__o21ai_2 _22960_ (.A1(_07406_),
    .A2(_07408_),
    .B1(_07085_),
    .Y(_07409_));
 sky130_fd_sc_hd__o2bb2a_2 _22961_ (.A1_N(_07097_),
    .A2_N(_07403_),
    .B1(_07405_),
    .B2(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__and3_2 _22962_ (.A(io_fetch_address[4]),
    .B(io_fetch_address[3]),
    .C(io_fetch_address[2]),
    .X(_07411_));
 sky130_fd_sc_hd__a21oi_2 _22963_ (.A1(io_fetch_address[3]),
    .A2(io_fetch_address[2]),
    .B1(io_fetch_address[4]),
    .Y(_07412_));
 sky130_fd_sc_hd__o2bb2a_2 _22964_ (.A1_N(_07391_),
    .A2_N(_07392_),
    .B1(_07411_),
    .B2(_07412_),
    .X(_07413_));
 sky130_fd_sc_hd__a211oi_2 _22965_ (.A1(_07368_),
    .A2(_07410_),
    .B1(_05246_),
    .C1(_07413_),
    .Y(_07414_));
 sky130_fd_sc_hd__a2111o_2 _22966_ (.A1(\execute.io_target_pc[4] ),
    .A2(_07346_),
    .B1(_07400_),
    .C1(_07414_),
    .D1(_07348_),
    .X(_07415_));
 sky130_fd_sc_hd__o311a_2 _22967_ (.A1(io_fetch_address[4]),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07415_),
    .C1(_06566_),
    .X(_01398_));
 sky130_fd_sc_hd__buf_1 _22968_ (.A(_06461_),
    .X(_07416_));
 sky130_fd_sc_hd__nand2_2 _22969_ (.A(_06461_),
    .B(_06041_),
    .Y(_07417_));
 sky130_fd_sc_hd__o22a_2 _22970_ (.A1(\csr._csr_read_data_T_8[5] ),
    .A2(_07416_),
    .B1(\csr.io_mret_vector[5] ),
    .B2(_07417_),
    .X(_07418_));
 sky130_fd_sc_hd__mux4_2 _22971_ (.A0(\fetch.bht.bhtTable_target_pc[0][5] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][5] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][5] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][5] ),
    .S0(_07098_),
    .S1(_07100_),
    .X(_07419_));
 sky130_fd_sc_hd__mux4_2 _22972_ (.A0(\fetch.bht.bhtTable_target_pc[4][5] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][5] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][5] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][5] ),
    .S0(_07098_),
    .S1(_07100_),
    .X(_07420_));
 sky130_fd_sc_hd__mux2_2 _22973_ (.A0(_07419_),
    .A1(_07420_),
    .S(_06633_),
    .X(_07421_));
 sky130_fd_sc_hd__mux4_2 _22974_ (.A0(\fetch.bht.bhtTable_target_pc[8][5] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][5] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][5] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][5] ),
    .S0(_07068_),
    .S1(_07110_),
    .X(_07422_));
 sky130_fd_sc_hd__and2_2 _22975_ (.A(_07422_),
    .B(_07371_),
    .X(_07423_));
 sky130_fd_sc_hd__mux4_2 _22976_ (.A0(\fetch.bht.bhtTable_target_pc[12][5] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][5] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][5] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][5] ),
    .S0(_07068_),
    .S1(_07110_),
    .X(_07424_));
 sky130_fd_sc_hd__a21o_2 _22977_ (.A1(_07075_),
    .A2(_07424_),
    .B1(_07084_),
    .X(_07425_));
 sky130_fd_sc_hd__o221a_2 _22978_ (.A1(_07127_),
    .A2(_07421_),
    .B1(_07423_),
    .B2(_07425_),
    .C1(_07367_),
    .X(_07426_));
 sky130_fd_sc_hd__and3_2 _22979_ (.A(io_fetch_address[5]),
    .B(io_fetch_address[4]),
    .C(_07393_),
    .X(_07427_));
 sky130_fd_sc_hd__a31o_2 _22980_ (.A1(io_fetch_address[4]),
    .A2(io_fetch_address[3]),
    .A3(io_fetch_address[2]),
    .B1(io_fetch_address[5]),
    .X(_07428_));
 sky130_fd_sc_hd__or3b_2 _22981_ (.A(_07367_),
    .B(_07427_),
    .C_N(_07428_),
    .X(_07429_));
 sky130_fd_sc_hd__or3b_2 _22982_ (.A(_07426_),
    .B(_10758_),
    .C_N(_07429_),
    .X(_07430_));
 sky130_fd_sc_hd__o311a_2 _22983_ (.A1(\execute.io_target_pc[5] ),
    .A2(_06032_),
    .A3(_07345_),
    .B1(_07418_),
    .C1(_07430_),
    .X(_07431_));
 sky130_fd_sc_hd__o21a_2 _22984_ (.A1(_07348_),
    .A2(_07431_),
    .B1(_10019_),
    .X(_07432_));
 sky130_fd_sc_hd__o31a_2 _22985_ (.A1(io_fetch_address[5]),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07432_),
    .X(_01399_));
 sky130_fd_sc_hd__mux4_2 _22986_ (.A0(\fetch.bht.bhtTable_target_pc[0][6] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][6] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][6] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][6] ),
    .S0(_07407_),
    .S1(_07115_),
    .X(_07433_));
 sky130_fd_sc_hd__mux2_2 _22987_ (.A0(\fetch.bht.bhtTable_target_pc[4][6] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][6] ),
    .S(_07123_),
    .X(_07434_));
 sky130_fd_sc_hd__and2b_2 _22988_ (.A_N(_07125_),
    .B(_07434_),
    .X(_07435_));
 sky130_fd_sc_hd__mux2_2 _22989_ (.A0(\fetch.bht.bhtTable_target_pc[6][6] ),
    .A1(\fetch.bht.bhtTable_target_pc[7][6] ),
    .S(_07069_),
    .X(_07436_));
 sky130_fd_sc_hd__a21o_2 _22990_ (.A1(_07112_),
    .A2(_07436_),
    .B1(_07082_),
    .X(_07437_));
 sky130_fd_sc_hd__o22a_2 _22991_ (.A1(_07076_),
    .A2(_07433_),
    .B1(_07435_),
    .B2(_07437_),
    .X(_07438_));
 sky130_fd_sc_hd__buf_1 _22992_ (.A(_07069_),
    .X(_07439_));
 sky130_fd_sc_hd__a21bo_2 _22993_ (.A1(_07439_),
    .A2(\fetch.bht.bhtTable_target_pc[15][6] ),
    .B1_N(_07125_),
    .X(_07440_));
 sky130_fd_sc_hd__and2b_2 _22994_ (.A_N(_07439_),
    .B(\fetch.bht.bhtTable_target_pc[14][6] ),
    .X(_07441_));
 sky130_fd_sc_hd__mux2_2 _22995_ (.A0(\fetch.bht.bhtTable_target_pc[12][6] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][6] ),
    .S(_07439_),
    .X(_07442_));
 sky130_fd_sc_hd__o221ai_2 _22996_ (.A1(_07440_),
    .A2(_07441_),
    .B1(_07112_),
    .B2(_07442_),
    .C1(_07076_),
    .Y(_07443_));
 sky130_fd_sc_hd__mux4_2 _22997_ (.A0(\fetch.bht.bhtTable_target_pc[8][6] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][6] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][6] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][6] ),
    .S0(_07108_),
    .S1(_07125_),
    .X(_07444_));
 sky130_fd_sc_hd__a21oi_2 _22998_ (.A1(_07444_),
    .A2(_07406_),
    .B1(_07085_),
    .Y(_07445_));
 sky130_fd_sc_hd__a2bb2o_2 _22999_ (.A1_N(_07097_),
    .A2_N(_07438_),
    .B1(_07443_),
    .B2(_07445_),
    .X(_07446_));
 sky130_fd_sc_hd__a31o_2 _23000_ (.A1(io_fetch_address[5]),
    .A2(io_fetch_address[4]),
    .A3(_07393_),
    .B1(io_fetch_address[6]),
    .X(_07447_));
 sky130_fd_sc_hd__nand2_2 _23001_ (.A(io_fetch_address[6]),
    .B(_07427_),
    .Y(_07448_));
 sky130_fd_sc_hd__a21oi_2 _23002_ (.A1(_07447_),
    .A2(_07448_),
    .B1(_07368_),
    .Y(_07449_));
 sky130_fd_sc_hd__a31o_2 _23003_ (.A1(_07391_),
    .A2(_07392_),
    .A3(_07446_),
    .B1(_07449_),
    .X(_07450_));
 sky130_fd_sc_hd__a22o_2 _23004_ (.A1(\csr._csr_read_data_T_8[6] ),
    .A2(_06038_),
    .B1(\csr.io_mret_vector[6] ),
    .B2(_06462_),
    .X(_07451_));
 sky130_fd_sc_hd__a311oi_2 _23005_ (.A1(\execute.io_target_pc[6] ),
    .A2(_05857_),
    .A3(_07091_),
    .B1(_07451_),
    .C1(_07348_),
    .Y(_07452_));
 sky130_fd_sc_hd__o21ai_2 _23006_ (.A1(_06248_),
    .A2(_07450_),
    .B1(_07452_),
    .Y(_07453_));
 sky130_fd_sc_hd__o311a_2 _23007_ (.A1(io_fetch_address[6]),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07453_),
    .C1(_06566_),
    .X(_01400_));
 sky130_fd_sc_hd__mux4_2 _23008_ (.A0(\fetch.bht.bhtTable_target_pc[0][7] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][7] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][7] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][7] ),
    .S0(_07407_),
    .S1(_07072_),
    .X(_07454_));
 sky130_fd_sc_hd__mux4_2 _23009_ (.A0(\fetch.bht.bhtTable_target_pc[4][7] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][7] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][7] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][7] ),
    .S0(_07407_),
    .S1(_07072_),
    .X(_07455_));
 sky130_fd_sc_hd__mux2_2 _23010_ (.A0(_07454_),
    .A1(_07455_),
    .S(_07076_),
    .X(_07456_));
 sky130_fd_sc_hd__a21bo_2 _23011_ (.A1(_07439_),
    .A2(\fetch.bht.bhtTable_target_pc[15][7] ),
    .B1_N(_07125_),
    .X(_07457_));
 sky130_fd_sc_hd__and2b_2 _23012_ (.A_N(_07439_),
    .B(\fetch.bht.bhtTable_target_pc[14][7] ),
    .X(_07458_));
 sky130_fd_sc_hd__mux2_2 _23013_ (.A0(\fetch.bht.bhtTable_target_pc[12][7] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][7] ),
    .S(_07439_),
    .X(_07459_));
 sky130_fd_sc_hd__o221ai_2 _23014_ (.A1(_07457_),
    .A2(_07458_),
    .B1(_07112_),
    .B2(_07459_),
    .C1(_07076_),
    .Y(_07460_));
 sky130_fd_sc_hd__mux4_2 _23015_ (.A0(\fetch.bht.bhtTable_target_pc[8][7] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][7] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][7] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][7] ),
    .S0(_07108_),
    .S1(_07125_),
    .X(_07461_));
 sky130_fd_sc_hd__a21oi_2 _23016_ (.A1(_07461_),
    .A2(_07406_),
    .B1(_07085_),
    .Y(_07462_));
 sky130_fd_sc_hd__a2bb2o_2 _23017_ (.A1_N(_07097_),
    .A2_N(_07456_),
    .B1(_07460_),
    .B2(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__and3_2 _23018_ (.A(io_fetch_address[7]),
    .B(io_fetch_address[6]),
    .C(_07427_),
    .X(_07464_));
 sky130_fd_sc_hd__a21oi_2 _23019_ (.A1(io_fetch_address[6]),
    .A2(_07427_),
    .B1(io_fetch_address[7]),
    .Y(_07465_));
 sky130_fd_sc_hd__o2bb2a_2 _23020_ (.A1_N(_07391_),
    .A2_N(_07392_),
    .B1(_07464_),
    .B2(_07465_),
    .X(_07466_));
 sky130_fd_sc_hd__a31o_2 _23021_ (.A1(_07391_),
    .A2(_07392_),
    .A3(_07463_),
    .B1(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__a22o_2 _23022_ (.A1(\csr._csr_read_data_T_8[7] ),
    .A2(_06038_),
    .B1(\csr.io_mret_vector[7] ),
    .B2(_06462_),
    .X(_07468_));
 sky130_fd_sc_hd__a311oi_2 _23023_ (.A1(\execute.io_target_pc[7] ),
    .A2(_05857_),
    .A3(_07091_),
    .B1(_07468_),
    .C1(_07347_),
    .Y(_07469_));
 sky130_fd_sc_hd__o21ai_2 _23024_ (.A1(_06248_),
    .A2(_07467_),
    .B1(_07469_),
    .Y(_07470_));
 sky130_fd_sc_hd__o311a_2 _23025_ (.A1(io_fetch_address[7]),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07470_),
    .C1(_06566_),
    .X(_01401_));
 sky130_fd_sc_hd__nor2_2 _23026_ (.A(io_fetch_address[8]),
    .B(_07464_),
    .Y(_07471_));
 sky130_fd_sc_hd__and4_2 _23027_ (.A(io_fetch_address[8]),
    .B(io_fetch_address[7]),
    .C(io_fetch_address[6]),
    .D(_07427_),
    .X(_07472_));
 sky130_fd_sc_hd__nor2_2 _23028_ (.A(_07471_),
    .B(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__mux4_2 _23029_ (.A0(\fetch.bht.bhtTable_target_pc[12][8] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][8] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][8] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][8] ),
    .S0(_07069_),
    .S1(_07111_),
    .X(_07474_));
 sky130_fd_sc_hd__a21o_2 _23030_ (.A1(_07076_),
    .A2(_07474_),
    .B1(_07084_),
    .X(_07475_));
 sky130_fd_sc_hd__a21bo_2 _23031_ (.A1(_07108_),
    .A2(\fetch.bht.bhtTable_target_pc[11][8] ),
    .B1_N(_07111_),
    .X(_07476_));
 sky130_fd_sc_hd__and2b_2 _23032_ (.A_N(_07108_),
    .B(\fetch.bht.bhtTable_target_pc[10][8] ),
    .X(_07477_));
 sky130_fd_sc_hd__mux2_2 _23033_ (.A0(\fetch.bht.bhtTable_target_pc[8][8] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][8] ),
    .S(_07407_),
    .X(_07478_));
 sky130_fd_sc_hd__o221a_2 _23034_ (.A1(_07476_),
    .A2(_07477_),
    .B1(_07112_),
    .B2(_07478_),
    .C1(_07082_),
    .X(_07479_));
 sky130_fd_sc_hd__mux4_2 _23035_ (.A0(\fetch.bht.bhtTable_target_pc[4][8] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][8] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][8] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][8] ),
    .S0(_07123_),
    .S1(_07101_),
    .X(_07480_));
 sky130_fd_sc_hd__mux4_2 _23036_ (.A0(\fetch.bht.bhtTable_target_pc[0][8] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][8] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][8] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][8] ),
    .S0(_07123_),
    .S1(_07101_),
    .X(_07481_));
 sky130_fd_sc_hd__mux2_2 _23037_ (.A0(_07480_),
    .A1(_07481_),
    .S(_07082_),
    .X(_07482_));
 sky130_fd_sc_hd__o22a_2 _23038_ (.A1(_07475_),
    .A2(_07479_),
    .B1(_07097_),
    .B2(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__mux2_2 _23039_ (.A0(_07473_),
    .A1(_07483_),
    .S(_07368_),
    .X(_07484_));
 sky130_fd_sc_hd__a22o_2 _23040_ (.A1(\csr._csr_read_data_T_8[8] ),
    .A2(_06038_),
    .B1(\csr.io_mret_vector[8] ),
    .B2(_06462_),
    .X(_07485_));
 sky130_fd_sc_hd__a311o_2 _23041_ (.A1(\execute.io_target_pc[8] ),
    .A2(_05864_),
    .A3(_07091_),
    .B1(_07485_),
    .C1(_07347_),
    .X(_07486_));
 sky130_fd_sc_hd__a31o_2 _23042_ (.A1(_06025_),
    .A2(_07484_),
    .A3(_07345_),
    .B1(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__o311a_2 _23043_ (.A1(io_fetch_address[8]),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07487_),
    .C1(_06566_),
    .X(_01402_));
 sky130_fd_sc_hd__a22o_2 _23044_ (.A1(\csr._csr_read_data_T_8[9] ),
    .A2(_06039_),
    .B1(\csr.io_mret_vector[9] ),
    .B2(_06463_),
    .X(_07488_));
 sky130_fd_sc_hd__mux4_2 _23045_ (.A0(\fetch.bht.bhtTable_target_pc[12][9] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][9] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][9] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][9] ),
    .S0(_07407_),
    .S1(_07115_),
    .X(_07489_));
 sky130_fd_sc_hd__mux4_2 _23046_ (.A0(\fetch.bht.bhtTable_target_pc[8][9] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][9] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][9] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][9] ),
    .S0(_07407_),
    .S1(_07115_),
    .X(_07490_));
 sky130_fd_sc_hd__mux2_2 _23047_ (.A0(_07489_),
    .A1(_07490_),
    .S(_07406_),
    .X(_07491_));
 sky130_fd_sc_hd__mux4_2 _23048_ (.A0(\fetch.bht.bhtTable_target_pc[0][9] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][9] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][9] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][9] ),
    .S0(_07108_),
    .S1(_07125_),
    .X(_07492_));
 sky130_fd_sc_hd__mux4_2 _23049_ (.A0(\fetch.bht.bhtTable_target_pc[4][9] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][9] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][9] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][9] ),
    .S0(_07123_),
    .S1(_07111_),
    .X(_07493_));
 sky130_fd_sc_hd__a21o_2 _23050_ (.A1(_07122_),
    .A2(_07493_),
    .B1(_07127_),
    .X(_07494_));
 sky130_fd_sc_hd__a21o_2 _23051_ (.A1(_07406_),
    .A2(_07492_),
    .B1(_07494_),
    .X(_07495_));
 sky130_fd_sc_hd__o21ai_2 _23052_ (.A1(_07085_),
    .A2(_07491_),
    .B1(_07495_),
    .Y(_07496_));
 sky130_fd_sc_hd__nand2_2 _23053_ (.A(_06718_),
    .B(_07472_),
    .Y(_07497_));
 sky130_fd_sc_hd__a41o_2 _23054_ (.A1(io_fetch_address[8]),
    .A2(io_fetch_address[7]),
    .A3(io_fetch_address[6]),
    .A4(_07427_),
    .B1(_06718_),
    .X(_07498_));
 sky130_fd_sc_hd__a21oi_2 _23055_ (.A1(_07497_),
    .A2(_07498_),
    .B1(_07368_),
    .Y(_07499_));
 sky130_fd_sc_hd__a211oi_2 _23056_ (.A1(_07368_),
    .A2(_07496_),
    .B1(_05246_),
    .C1(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__a2111o_2 _23057_ (.A1(\execute.io_target_pc[9] ),
    .A2(_07346_),
    .B1(_07488_),
    .C1(_07500_),
    .D1(_07348_),
    .X(_07501_));
 sky130_fd_sc_hd__o311a_2 _23058_ (.A1(_06718_),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07501_),
    .C1(_06566_),
    .X(_01403_));
 sky130_fd_sc_hd__a22o_2 _23059_ (.A1(\csr._csr_read_data_T_8[10] ),
    .A2(_06039_),
    .B1(\csr.io_mret_vector[10] ),
    .B2(_06463_),
    .X(_07502_));
 sky130_fd_sc_hd__a21oi_2 _23060_ (.A1(_06718_),
    .A2(_07472_),
    .B1(io_fetch_address[10]),
    .Y(_07503_));
 sky130_fd_sc_hd__and3_2 _23061_ (.A(io_fetch_address[10]),
    .B(_06718_),
    .C(_07472_),
    .X(_07504_));
 sky130_fd_sc_hd__o2bb2a_2 _23062_ (.A1_N(_07391_),
    .A2_N(_07392_),
    .B1(_07503_),
    .B2(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__mux4_2 _23063_ (.A0(\fetch.bht.bhtTable_target_pc[4][10] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][10] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][10] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][10] ),
    .S0(_07108_),
    .S1(_07115_),
    .X(_07506_));
 sky130_fd_sc_hd__mux4_2 _23064_ (.A0(\fetch.bht.bhtTable_target_pc[0][10] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][10] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][10] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][10] ),
    .S0(_07407_),
    .S1(_07115_),
    .X(_07507_));
 sky130_fd_sc_hd__mux2_2 _23065_ (.A0(_07506_),
    .A1(_07507_),
    .S(_07406_),
    .X(_07508_));
 sky130_fd_sc_hd__mux2_2 _23066_ (.A0(\fetch.bht.bhtTable_target_pc[12][10] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][10] ),
    .S(_07123_),
    .X(_07509_));
 sky130_fd_sc_hd__and2b_2 _23067_ (.A_N(_07125_),
    .B(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__or2b_2 _23068_ (.A(\fetch.bht.bhtTable_target_pc[15][10] ),
    .B_N(_07407_),
    .X(_07511_));
 sky130_fd_sc_hd__o211a_2 _23069_ (.A1(_07439_),
    .A2(\fetch.bht.bhtTable_target_pc[14][10] ),
    .B1(_07125_),
    .C1(_07511_),
    .X(_07512_));
 sky130_fd_sc_hd__mux2_2 _23070_ (.A0(\fetch.bht.bhtTable_target_pc[10][10] ),
    .A1(\fetch.bht.bhtTable_target_pc[11][10] ),
    .S(_07069_),
    .X(_07513_));
 sky130_fd_sc_hd__mux2_2 _23071_ (.A0(\fetch.bht.bhtTable_target_pc[8][10] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][10] ),
    .S(_07119_),
    .X(_07514_));
 sky130_fd_sc_hd__and2b_2 _23072_ (.A_N(_07072_),
    .B(_07514_),
    .X(_07515_));
 sky130_fd_sc_hd__a211o_2 _23073_ (.A1(_07513_),
    .A2(_07112_),
    .B1(_07122_),
    .C1(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__o311a_2 _23074_ (.A1(_07406_),
    .A2(_07510_),
    .A3(_07512_),
    .B1(_07097_),
    .C1(_07516_),
    .X(_07517_));
 sky130_fd_sc_hd__a211oi_2 _23075_ (.A1(_07085_),
    .A2(_07508_),
    .B1(_07517_),
    .C1(_07130_),
    .Y(_07518_));
 sky130_fd_sc_hd__nor3_2 _23076_ (.A(_05246_),
    .B(_07505_),
    .C(_07518_),
    .Y(_07519_));
 sky130_fd_sc_hd__a2111o_2 _23077_ (.A1(\execute.io_target_pc[10] ),
    .A2(_07346_),
    .B1(_07502_),
    .C1(_07519_),
    .D1(_07348_),
    .X(_07520_));
 sky130_fd_sc_hd__o311a_2 _23078_ (.A1(io_fetch_address[10]),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07520_),
    .C1(_06566_),
    .X(_01404_));
 sky130_fd_sc_hd__a22o_2 _23079_ (.A1(\csr._csr_read_data_T_8[11] ),
    .A2(_06039_),
    .B1(\csr.io_mret_vector[11] ),
    .B2(_06463_),
    .X(_07521_));
 sky130_fd_sc_hd__mux4_2 _23080_ (.A0(\fetch.bht.bhtTable_target_pc[12][11] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][11] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][11] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][11] ),
    .S0(_07069_),
    .S1(_07111_),
    .X(_07522_));
 sky130_fd_sc_hd__mux4_2 _23081_ (.A0(\fetch.bht.bhtTable_target_pc[8][11] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][11] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][11] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][11] ),
    .S0(_07123_),
    .S1(_07111_),
    .X(_07523_));
 sky130_fd_sc_hd__mux2_2 _23082_ (.A0(_07522_),
    .A1(_07523_),
    .S(_07082_),
    .X(_07524_));
 sky130_fd_sc_hd__mux4_2 _23083_ (.A0(\fetch.bht.bhtTable_target_pc[0][11] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][11] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][11] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][11] ),
    .S0(_07407_),
    .S1(_07115_),
    .X(_07525_));
 sky130_fd_sc_hd__a21oi_2 _23084_ (.A1(_07525_),
    .A2(_07406_),
    .B1(_07097_),
    .Y(_07526_));
 sky130_fd_sc_hd__mux4_2 _23085_ (.A0(\fetch.bht.bhtTable_target_pc[4][11] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][11] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][11] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][11] ),
    .S0(_07108_),
    .S1(_07125_),
    .X(_07527_));
 sky130_fd_sc_hd__nand2_2 _23086_ (.A(_07076_),
    .B(_07527_),
    .Y(_07528_));
 sky130_fd_sc_hd__a2bb2o_2 _23087_ (.A1_N(_07085_),
    .A2_N(_07524_),
    .B1(_07526_),
    .B2(_07528_),
    .X(_07529_));
 sky130_fd_sc_hd__and4_2 _23088_ (.A(io_fetch_address[11]),
    .B(io_fetch_address[10]),
    .C(io_fetch_address[9]),
    .D(_07472_),
    .X(_07530_));
 sky130_fd_sc_hd__nor2_2 _23089_ (.A(io_fetch_address[11]),
    .B(_07504_),
    .Y(_07531_));
 sky130_fd_sc_hd__o2bb2a_2 _23090_ (.A1_N(_07391_),
    .A2_N(_07392_),
    .B1(_07530_),
    .B2(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__a211oi_2 _23091_ (.A1(_07368_),
    .A2(_07529_),
    .B1(_05246_),
    .C1(_07532_),
    .Y(_07533_));
 sky130_fd_sc_hd__a2111o_2 _23092_ (.A1(\execute.io_target_pc[11] ),
    .A2(_07346_),
    .B1(_07521_),
    .C1(_07533_),
    .D1(_07348_),
    .X(_07534_));
 sky130_fd_sc_hd__buf_1 _23093_ (.A(_09956_),
    .X(_07535_));
 sky130_fd_sc_hd__o311a_2 _23094_ (.A1(io_fetch_address[11]),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07534_),
    .C1(_07535_),
    .X(_01405_));
 sky130_fd_sc_hd__buf_1 _23095_ (.A(_06248_),
    .X(_07536_));
 sky130_fd_sc_hd__buf_1 _23096_ (.A(_03500_),
    .X(_07537_));
 sky130_fd_sc_hd__a22o_2 _23097_ (.A1(\csr._csr_read_data_T_8[12] ),
    .A2(_06039_),
    .B1(\csr.io_mret_vector[12] ),
    .B2(_06463_),
    .X(_07538_));
 sky130_fd_sc_hd__mux4_2 _23098_ (.A0(\fetch.bht.bhtTable_target_pc[4][12] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][12] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][12] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][12] ),
    .S0(_07107_),
    .S1(_07114_),
    .X(_07539_));
 sky130_fd_sc_hd__mux4_2 _23099_ (.A0(\fetch.bht.bhtTable_target_pc[0][12] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][12] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][12] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][12] ),
    .S0(_07107_),
    .S1(_07071_),
    .X(_07540_));
 sky130_fd_sc_hd__mux2_2 _23100_ (.A0(_07539_),
    .A1(_07540_),
    .S(_07371_),
    .X(_07541_));
 sky130_fd_sc_hd__mux4_2 _23101_ (.A0(\fetch.bht.bhtTable_target_pc[8][12] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][12] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][12] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][12] ),
    .S0(_07107_),
    .S1(_07114_),
    .X(_07542_));
 sky130_fd_sc_hd__mux2_2 _23102_ (.A0(\fetch.bht.bhtTable_target_pc[12][12] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][12] ),
    .S(_07068_),
    .X(_07543_));
 sky130_fd_sc_hd__and2b_2 _23103_ (.A_N(_07101_),
    .B(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__mux2_2 _23104_ (.A0(\fetch.bht.bhtTable_target_pc[14][12] ),
    .A1(\fetch.bht.bhtTable_target_pc[15][12] ),
    .S(_07119_),
    .X(_07545_));
 sky130_fd_sc_hd__a21o_2 _23105_ (.A1(_07545_),
    .A2(_07111_),
    .B1(_07081_),
    .X(_07546_));
 sky130_fd_sc_hd__o221a_2 _23106_ (.A1(_07122_),
    .A2(_07542_),
    .B1(_07544_),
    .B2(_07546_),
    .C1(_07127_),
    .X(_07547_));
 sky130_fd_sc_hd__a21oi_2 _23107_ (.A1(_07541_),
    .A2(_07085_),
    .B1(_07547_),
    .Y(_07548_));
 sky130_fd_sc_hd__a41o_2 _23108_ (.A1(io_fetch_address[11]),
    .A2(io_fetch_address[10]),
    .A3(_06718_),
    .A4(_07472_),
    .B1(io_fetch_address[12]),
    .X(_07549_));
 sky130_fd_sc_hd__nand2_2 _23109_ (.A(io_fetch_address[12]),
    .B(_07530_),
    .Y(_07550_));
 sky130_fd_sc_hd__nand3_2 _23110_ (.A(_07130_),
    .B(_07549_),
    .C(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__o211ai_2 _23111_ (.A1(_07130_),
    .A2(_07548_),
    .B1(_07551_),
    .C1(_03592_),
    .Y(_07552_));
 sky130_fd_sc_hd__o211a_2 _23112_ (.A1(\execute.io_target_pc[12] ),
    .A2(_07345_),
    .B1(_05864_),
    .C1(_07552_),
    .X(_07553_));
 sky130_fd_sc_hd__or3_2 _23113_ (.A(_07347_),
    .B(_07538_),
    .C(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__o311a_2 _23114_ (.A1(io_fetch_address[12]),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07554_),
    .C1(_07535_),
    .X(_01406_));
 sky130_fd_sc_hd__buf_1 _23115_ (.A(_07098_),
    .X(_07555_));
 sky130_fd_sc_hd__mux4_2 _23116_ (.A0(\fetch.bht.bhtTable_target_pc[8][13] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][13] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][13] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][13] ),
    .S0(_07555_),
    .S1(_07114_),
    .X(_07556_));
 sky130_fd_sc_hd__o21ai_2 _23117_ (.A1(_07122_),
    .A2(_07556_),
    .B1(_07127_),
    .Y(_07557_));
 sky130_fd_sc_hd__mux4_2 _23118_ (.A0(\fetch.bht.bhtTable_target_pc[12][13] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][13] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][13] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][13] ),
    .S0(_07099_),
    .S1(_07101_),
    .X(_07558_));
 sky130_fd_sc_hd__nor2_2 _23119_ (.A(_07082_),
    .B(_07558_),
    .Y(_07559_));
 sky130_fd_sc_hd__mux4_2 _23120_ (.A0(\fetch.bht.bhtTable_target_pc[4][13] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][13] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][13] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][13] ),
    .S0(_07099_),
    .S1(_07101_),
    .X(_07560_));
 sky130_fd_sc_hd__mux2_2 _23121_ (.A0(\fetch.bht.bhtTable_target_pc[2][13] ),
    .A1(\fetch.bht.bhtTable_target_pc[3][13] ),
    .S(_07119_),
    .X(_07561_));
 sky130_fd_sc_hd__mux2_2 _23122_ (.A0(\fetch.bht.bhtTable_target_pc[0][13] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][13] ),
    .S(_07067_),
    .X(_07562_));
 sky130_fd_sc_hd__and2b_2 _23123_ (.A_N(_07071_),
    .B(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__a211o_2 _23124_ (.A1(_07561_),
    .A2(_07072_),
    .B1(_07075_),
    .C1(_07563_),
    .X(_07564_));
 sky130_fd_sc_hd__o21ai_2 _23125_ (.A1(_07082_),
    .A2(_07560_),
    .B1(_07564_),
    .Y(_07565_));
 sky130_fd_sc_hd__o22a_2 _23126_ (.A1(_07557_),
    .A2(_07559_),
    .B1(_07097_),
    .B2(_07565_),
    .X(_07566_));
 sky130_fd_sc_hd__and3_2 _23127_ (.A(io_fetch_address[13]),
    .B(io_fetch_address[12]),
    .C(_07530_),
    .X(_07567_));
 sky130_fd_sc_hd__a21oi_2 _23128_ (.A1(io_fetch_address[12]),
    .A2(_07530_),
    .B1(io_fetch_address[13]),
    .Y(_07568_));
 sky130_fd_sc_hd__o2bb2a_2 _23129_ (.A1_N(_07391_),
    .A2_N(_07392_),
    .B1(_07567_),
    .B2(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__a211oi_2 _23130_ (.A1(_07368_),
    .A2(_07566_),
    .B1(_05246_),
    .C1(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__a221o_2 _23131_ (.A1(\csr._csr_read_data_T_8[13] ),
    .A2(_06039_),
    .B1(\csr.io_mret_vector[13] ),
    .B2(_06463_),
    .C1(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__a211o_2 _23132_ (.A1(\execute.io_target_pc[13] ),
    .A2(_07346_),
    .B1(_07348_),
    .C1(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__o311a_2 _23133_ (.A1(io_fetch_address[13]),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07572_),
    .C1(_07535_),
    .X(_01407_));
 sky130_fd_sc_hd__buf_1 _23134_ (.A(_07345_),
    .X(_07573_));
 sky130_fd_sc_hd__mux4_2 _23135_ (.A0(\fetch.bht.bhtTable_target_pc[0][14] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][14] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][14] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][14] ),
    .S0(_07099_),
    .S1(_07103_),
    .X(_07574_));
 sky130_fd_sc_hd__mux4_2 _23136_ (.A0(\fetch.bht.bhtTable_target_pc[4][14] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][14] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][14] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][14] ),
    .S0(_07099_),
    .S1(_07103_),
    .X(_07575_));
 sky130_fd_sc_hd__mux2_2 _23137_ (.A0(_07574_),
    .A1(_07575_),
    .S(_07122_),
    .X(_07576_));
 sky130_fd_sc_hd__mux4_2 _23138_ (.A0(\fetch.bht.bhtTable_target_pc[8][14] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][14] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][14] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][14] ),
    .S0(_07123_),
    .S1(_07111_),
    .X(_07577_));
 sky130_fd_sc_hd__and2_2 _23139_ (.A(_07577_),
    .B(_07082_),
    .X(_07578_));
 sky130_fd_sc_hd__mux4_2 _23140_ (.A0(\fetch.bht.bhtTable_target_pc[12][14] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][14] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][14] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][14] ),
    .S0(_07069_),
    .S1(_07111_),
    .X(_07579_));
 sky130_fd_sc_hd__a21o_2 _23141_ (.A1(_07122_),
    .A2(_07579_),
    .B1(_07084_),
    .X(_07580_));
 sky130_fd_sc_hd__o221a_2 _23142_ (.A1(_07097_),
    .A2(_07576_),
    .B1(_07578_),
    .B2(_07580_),
    .C1(_07368_),
    .X(_07581_));
 sky130_fd_sc_hd__and4_2 _23143_ (.A(io_fetch_address[14]),
    .B(io_fetch_address[13]),
    .C(io_fetch_address[12]),
    .D(_07530_),
    .X(_07582_));
 sky130_fd_sc_hd__nor2_2 _23144_ (.A(io_fetch_address[14]),
    .B(_07567_),
    .Y(_07583_));
 sky130_fd_sc_hd__a211oi_2 _23145_ (.A1(_07391_),
    .A2(_07392_),
    .B1(_07582_),
    .C1(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__or4_2 _23146_ (.A(\execute.io_target_pc[14] ),
    .B(_06037_),
    .C(_10970_),
    .D(_03592_),
    .X(_07585_));
 sky130_fd_sc_hd__o221a_2 _23147_ (.A1(\csr._csr_read_data_T_8[14] ),
    .A2(_06461_),
    .B1(\csr.io_mret_vector[14] ),
    .B2(_07417_),
    .C1(_07585_),
    .X(_07586_));
 sky130_fd_sc_hd__o31a_2 _23148_ (.A1(_07581_),
    .A2(_05246_),
    .A3(_07584_),
    .B1(_07586_),
    .X(_07587_));
 sky130_fd_sc_hd__a31o_2 _23149_ (.A1(_06025_),
    .A2(_07573_),
    .A3(_03546_),
    .B1(_07587_),
    .X(_07588_));
 sky130_fd_sc_hd__o311a_2 _23150_ (.A1(io_fetch_address[14]),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07588_),
    .C1(_07535_),
    .X(_01408_));
 sky130_fd_sc_hd__nand2_2 _23151_ (.A(io_fetch_address[15]),
    .B(_07582_),
    .Y(_07589_));
 sky130_fd_sc_hd__a41o_2 _23152_ (.A1(io_fetch_address[14]),
    .A2(io_fetch_address[13]),
    .A3(io_fetch_address[12]),
    .A4(_07530_),
    .B1(io_fetch_address[15]),
    .X(_07590_));
 sky130_fd_sc_hd__and3_2 _23153_ (.A(_07130_),
    .B(_07589_),
    .C(_07590_),
    .X(_07591_));
 sky130_fd_sc_hd__mux4_2 _23154_ (.A0(\fetch.bht.bhtTable_target_pc[4][15] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][15] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][15] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][15] ),
    .S0(_07555_),
    .S1(_07114_),
    .X(_07592_));
 sky130_fd_sc_hd__mux4_2 _23155_ (.A0(\fetch.bht.bhtTable_target_pc[0][15] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][15] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][15] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][15] ),
    .S0(_07107_),
    .S1(_07114_),
    .X(_07593_));
 sky130_fd_sc_hd__mux4_2 _23156_ (.A0(\fetch.bht.bhtTable_target_pc[12][15] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][15] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][15] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][15] ),
    .S0(_07107_),
    .S1(_07114_),
    .X(_07594_));
 sky130_fd_sc_hd__mux4_2 _23157_ (.A0(\fetch.bht.bhtTable_target_pc[8][15] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][15] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][15] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][15] ),
    .S0(_07555_),
    .S1(_07114_),
    .X(_07595_));
 sky130_fd_sc_hd__mux4_2 _23158_ (.A0(_07592_),
    .A1(_07593_),
    .A2(_07594_),
    .A3(_07595_),
    .S0(_07371_),
    .S1(_07127_),
    .X(_07596_));
 sky130_fd_sc_hd__and2b_2 _23159_ (.A_N(_07130_),
    .B(_07596_),
    .X(_07597_));
 sky130_fd_sc_hd__or4_2 _23160_ (.A(\execute.io_target_pc[15] ),
    .B(_06037_),
    .C(_10970_),
    .D(_03592_),
    .X(_07598_));
 sky130_fd_sc_hd__o221a_2 _23161_ (.A1(\csr._csr_read_data_T_8[15] ),
    .A2(_06461_),
    .B1(\csr.io_mret_vector[15] ),
    .B2(_07417_),
    .C1(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__o31a_2 _23162_ (.A1(_05246_),
    .A2(_07591_),
    .A3(_07597_),
    .B1(_07599_),
    .X(_07600_));
 sky130_fd_sc_hd__a31o_2 _23163_ (.A1(_06025_),
    .A2(_07573_),
    .A3(_03546_),
    .B1(_07600_),
    .X(_07601_));
 sky130_fd_sc_hd__o311a_2 _23164_ (.A1(io_fetch_address[15]),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07601_),
    .C1(_07535_),
    .X(_01409_));
 sky130_fd_sc_hd__mux4_2 _23165_ (.A0(\fetch.bht.bhtTable_target_pc[4][16] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][16] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][16] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][16] ),
    .S0(_07439_),
    .S1(_07112_),
    .X(_07602_));
 sky130_fd_sc_hd__mux4_2 _23166_ (.A0(\fetch.bht.bhtTable_target_pc[0][16] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][16] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][16] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][16] ),
    .S0(_07439_),
    .S1(_07112_),
    .X(_07603_));
 sky130_fd_sc_hd__mux2_2 _23167_ (.A0(_07602_),
    .A1(_07603_),
    .S(_07406_),
    .X(_07604_));
 sky130_fd_sc_hd__mux4_2 _23168_ (.A0(\fetch.bht.bhtTable_target_pc[12][16] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][16] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][16] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][16] ),
    .S0(_07439_),
    .S1(_07112_),
    .X(_07605_));
 sky130_fd_sc_hd__mux2_2 _23169_ (.A0(\fetch.bht.bhtTable_target_pc[10][16] ),
    .A1(\fetch.bht.bhtTable_target_pc[11][16] ),
    .S(_07108_),
    .X(_07606_));
 sky130_fd_sc_hd__mux2_2 _23170_ (.A0(\fetch.bht.bhtTable_target_pc[8][16] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][16] ),
    .S(_07099_),
    .X(_07607_));
 sky130_fd_sc_hd__and2b_2 _23171_ (.A_N(_07115_),
    .B(_07607_),
    .X(_07608_));
 sky130_fd_sc_hd__a211o_2 _23172_ (.A1(_07606_),
    .A2(_07112_),
    .B1(_07076_),
    .C1(_07608_),
    .X(_07609_));
 sky130_fd_sc_hd__o211a_2 _23173_ (.A1(_07406_),
    .A2(_07605_),
    .B1(_07097_),
    .C1(_07609_),
    .X(_07610_));
 sky130_fd_sc_hd__a211o_2 _23174_ (.A1(_07085_),
    .A2(_07604_),
    .B1(_07610_),
    .C1(_07130_),
    .X(_07611_));
 sky130_fd_sc_hd__a21oi_2 _23175_ (.A1(io_fetch_address[15]),
    .A2(_07582_),
    .B1(io_fetch_address[16]),
    .Y(_07612_));
 sky130_fd_sc_hd__and3_2 _23176_ (.A(io_fetch_address[16]),
    .B(io_fetch_address[15]),
    .C(_07582_),
    .X(_07613_));
 sky130_fd_sc_hd__nor2_2 _23177_ (.A(_07612_),
    .B(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__o211a_2 _23178_ (.A1(_07368_),
    .A2(_07614_),
    .B1(_05864_),
    .C1(_07345_),
    .X(_07615_));
 sky130_fd_sc_hd__a22o_2 _23179_ (.A1(\csr._csr_read_data_T_8[16] ),
    .A2(_06038_),
    .B1(\csr.io_mret_vector[16] ),
    .B2(_06462_),
    .X(_07616_));
 sky130_fd_sc_hd__a311o_2 _23180_ (.A1(\execute.io_target_pc[16] ),
    .A2(_05864_),
    .A3(_07091_),
    .B1(_07616_),
    .C1(_07347_),
    .X(_07617_));
 sky130_fd_sc_hd__a21o_2 _23181_ (.A1(_07611_),
    .A2(_07615_),
    .B1(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__o311a_2 _23182_ (.A1(io_fetch_address[16]),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07618_),
    .C1(_07535_),
    .X(_01410_));
 sky130_fd_sc_hd__buf_1 _23183_ (.A(_05864_),
    .X(_07619_));
 sky130_fd_sc_hd__buf_1 _23184_ (.A(_10672_),
    .X(_07620_));
 sky130_fd_sc_hd__buf_1 _23185_ (.A(_07417_),
    .X(_07621_));
 sky130_fd_sc_hd__mux4_2 _23186_ (.A0(\fetch.bht.bhtTable_target_pc[12][17] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][17] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][17] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][17] ),
    .S0(_07384_),
    .S1(_07113_),
    .X(_07622_));
 sky130_fd_sc_hd__mux4_2 _23187_ (.A0(\fetch.bht.bhtTable_target_pc[8][17] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][17] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][17] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][17] ),
    .S0(_07106_),
    .S1(_07386_),
    .X(_07623_));
 sky130_fd_sc_hd__mux4_2 _23188_ (.A0(\fetch.bht.bhtTable_target_pc[4][17] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][17] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][17] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][17] ),
    .S0(_07384_),
    .S1(_07386_),
    .X(_07624_));
 sky130_fd_sc_hd__mux4_2 _23189_ (.A0(\fetch.bht.bhtTable_target_pc[0][17] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][17] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][17] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][17] ),
    .S0(_07384_),
    .S1(_07113_),
    .X(_07625_));
 sky130_fd_sc_hd__mux4_2 _23190_ (.A0(_07622_),
    .A1(_07623_),
    .A2(_07624_),
    .A3(_07625_),
    .S0(_07080_),
    .S1(_06637_),
    .X(_07626_));
 sky130_fd_sc_hd__a31o_2 _23191_ (.A1(io_fetch_address[16]),
    .A2(io_fetch_address[15]),
    .A3(_07582_),
    .B1(_06887_),
    .X(_07627_));
 sky130_fd_sc_hd__nand2_2 _23192_ (.A(_06887_),
    .B(_07613_),
    .Y(_07628_));
 sky130_fd_sc_hd__a22o_2 _23193_ (.A1(_07627_),
    .A2(_07628_),
    .B1(_07391_),
    .B2(_07392_),
    .X(_07629_));
 sky130_fd_sc_hd__o211a_2 _23194_ (.A1(_07626_),
    .A2(_07130_),
    .B1(_03592_),
    .C1(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__a211o_2 _23195_ (.A1(\execute.io_target_pc[17] ),
    .A2(_07091_),
    .B1(_06032_),
    .C1(_07630_),
    .X(_07631_));
 sky130_fd_sc_hd__o221a_2 _23196_ (.A1(\csr._csr_read_data_T_8[17] ),
    .A2(_06480_),
    .B1(\csr.io_mret_vector[17] ),
    .B2(_07621_),
    .C1(_07631_),
    .X(_07632_));
 sky130_fd_sc_hd__a31o_2 _23197_ (.A1(_07619_),
    .A2(_07573_),
    .A3(_07620_),
    .B1(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__o311a_2 _23198_ (.A1(_06887_),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07633_),
    .C1(_07535_),
    .X(_01411_));
 sky130_fd_sc_hd__a22o_2 _23199_ (.A1(\csr._csr_read_data_T_8[18] ),
    .A2(_06038_),
    .B1(\csr.io_mret_vector[18] ),
    .B2(_06463_),
    .X(_07634_));
 sky130_fd_sc_hd__a21oi_2 _23200_ (.A1(_06887_),
    .A2(_07613_),
    .B1(io_fetch_address[18]),
    .Y(_07635_));
 sky130_fd_sc_hd__and3_2 _23201_ (.A(io_fetch_address[18]),
    .B(_06887_),
    .C(_07613_),
    .X(_07636_));
 sky130_fd_sc_hd__nor2_2 _23202_ (.A(_07635_),
    .B(_07636_),
    .Y(_07637_));
 sky130_fd_sc_hd__mux4_2 _23203_ (.A0(\fetch.bht.bhtTable_target_pc[0][18] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][18] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][18] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][18] ),
    .S0(_07098_),
    .S1(_07113_),
    .X(_07638_));
 sky130_fd_sc_hd__mux4_2 _23204_ (.A0(\fetch.bht.bhtTable_target_pc[4][18] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][18] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][18] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][18] ),
    .S0(_07384_),
    .S1(_07113_),
    .X(_07639_));
 sky130_fd_sc_hd__mux2_2 _23205_ (.A0(_07638_),
    .A1(_07639_),
    .S(_06633_),
    .X(_07640_));
 sky130_fd_sc_hd__mux2_2 _23206_ (.A0(\fetch.bht.bhtTable_target_pc[8][18] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][18] ),
    .S(_07067_),
    .X(_07641_));
 sky130_fd_sc_hd__o21a_2 _23207_ (.A1(_07110_),
    .A2(_07641_),
    .B1(_07080_),
    .X(_07642_));
 sky130_fd_sc_hd__mux2_2 _23208_ (.A0(\fetch.bht.bhtTable_target_pc[10][18] ),
    .A1(\fetch.bht.bhtTable_target_pc[11][18] ),
    .S(_07067_),
    .X(_07643_));
 sky130_fd_sc_hd__or2b_2 _23209_ (.A(_07643_),
    .B_N(_07110_),
    .X(_07644_));
 sky130_fd_sc_hd__mux4_2 _23210_ (.A0(\fetch.bht.bhtTable_target_pc[12][18] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][18] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][18] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][18] ),
    .S0(_07098_),
    .S1(_07100_),
    .X(_07645_));
 sky130_fd_sc_hd__a221o_2 _23211_ (.A1(_07642_),
    .A2(_07644_),
    .B1(_07645_),
    .B2(_07075_),
    .C1(_06637_),
    .X(_07646_));
 sky130_fd_sc_hd__o211a_2 _23212_ (.A1(_07127_),
    .A2(_07640_),
    .B1(_07646_),
    .C1(_07367_),
    .X(_07647_));
 sky130_fd_sc_hd__a211o_2 _23213_ (.A1(_07130_),
    .A2(_07637_),
    .B1(_07647_),
    .C1(_07090_),
    .X(_07648_));
 sky130_fd_sc_hd__o211a_2 _23214_ (.A1(\execute.io_target_pc[18] ),
    .A2(_03592_),
    .B1(_03590_),
    .C1(_07648_),
    .X(_07649_));
 sky130_fd_sc_hd__or3_2 _23215_ (.A(_07347_),
    .B(_07634_),
    .C(_07649_),
    .X(_07650_));
 sky130_fd_sc_hd__o311a_2 _23216_ (.A1(io_fetch_address[18]),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07650_),
    .C1(_07535_),
    .X(_01412_));
 sky130_fd_sc_hd__and4_2 _23217_ (.A(io_fetch_address[19]),
    .B(io_fetch_address[18]),
    .C(io_fetch_address[17]),
    .D(_07613_),
    .X(_07651_));
 sky130_fd_sc_hd__a31o_2 _23218_ (.A1(io_fetch_address[18]),
    .A2(_06887_),
    .A3(_07613_),
    .B1(io_fetch_address[19]),
    .X(_07652_));
 sky130_fd_sc_hd__and3b_2 _23219_ (.A_N(_07651_),
    .B(_07652_),
    .C(_07063_),
    .X(_07653_));
 sky130_fd_sc_hd__a211o_2 _23220_ (.A1(\execute.io_target_pc[19] ),
    .A2(_10757_),
    .B1(_10970_),
    .C1(_06037_),
    .X(_07654_));
 sky130_fd_sc_hd__and2b_2 _23221_ (.A_N(_07107_),
    .B(\fetch.bht.bhtTable_target_pc[14][19] ),
    .X(_07655_));
 sky130_fd_sc_hd__buf_1 _23222_ (.A(_07070_),
    .X(_07656_));
 sky130_fd_sc_hd__a21bo_2 _23223_ (.A1(_07555_),
    .A2(\fetch.bht.bhtTable_target_pc[15][19] ),
    .B1_N(_07656_),
    .X(_07657_));
 sky130_fd_sc_hd__mux2_2 _23224_ (.A0(\fetch.bht.bhtTable_target_pc[12][19] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][19] ),
    .S(_07119_),
    .X(_07658_));
 sky130_fd_sc_hd__o221a_2 _23225_ (.A1(_07655_),
    .A2(_07657_),
    .B1(_07111_),
    .B2(_07658_),
    .C1(_07075_),
    .X(_07659_));
 sky130_fd_sc_hd__mux2_2 _23226_ (.A0(\fetch.bht.bhtTable_target_pc[10][19] ),
    .A1(\fetch.bht.bhtTable_target_pc[11][19] ),
    .S(_07067_),
    .X(_07660_));
 sky130_fd_sc_hd__or2b_2 _23227_ (.A(_07660_),
    .B_N(_07071_),
    .X(_07661_));
 sky130_fd_sc_hd__mux2_2 _23228_ (.A0(\fetch.bht.bhtTable_target_pc[8][19] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][19] ),
    .S(_07067_),
    .X(_07662_));
 sky130_fd_sc_hd__or2_2 _23229_ (.A(_07110_),
    .B(_07662_),
    .X(_07663_));
 sky130_fd_sc_hd__a31o_2 _23230_ (.A1(_07371_),
    .A2(_07661_),
    .A3(_07663_),
    .B1(_06637_),
    .X(_07664_));
 sky130_fd_sc_hd__mux2_2 _23231_ (.A0(\fetch.bht.bhtTable_target_pc[2][19] ),
    .A1(\fetch.bht.bhtTable_target_pc[3][19] ),
    .S(_07067_),
    .X(_07665_));
 sky130_fd_sc_hd__or2b_2 _23232_ (.A(_07665_),
    .B_N(_07110_),
    .X(_07666_));
 sky130_fd_sc_hd__mux2_2 _23233_ (.A0(\fetch.bht.bhtTable_target_pc[0][19] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][19] ),
    .S(_07067_),
    .X(_07667_));
 sky130_fd_sc_hd__o21a_2 _23234_ (.A1(_07110_),
    .A2(_07667_),
    .B1(_07080_),
    .X(_07668_));
 sky130_fd_sc_hd__buf_1 _23235_ (.A(_07066_),
    .X(_07669_));
 sky130_fd_sc_hd__mux4_2 _23236_ (.A0(\fetch.bht.bhtTable_target_pc[4][19] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][19] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][19] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][19] ),
    .S0(_07669_),
    .S1(_07100_),
    .X(_07670_));
 sky130_fd_sc_hd__a221o_2 _23237_ (.A1(_07666_),
    .A2(_07668_),
    .B1(_07670_),
    .B2(_07075_),
    .C1(_06740_),
    .X(_07671_));
 sky130_fd_sc_hd__o211a_2 _23238_ (.A1(_07659_),
    .A2(_07664_),
    .B1(_07671_),
    .C1(_07088_),
    .X(_07672_));
 sky130_fd_sc_hd__or3_2 _23239_ (.A(_07653_),
    .B(_07654_),
    .C(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__o221a_2 _23240_ (.A1(\csr._csr_read_data_T_8[19] ),
    .A2(_06480_),
    .B1(\csr.io_mret_vector[19] ),
    .B2(_07621_),
    .C1(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__a31o_2 _23241_ (.A1(_07619_),
    .A2(_07573_),
    .A3(_07620_),
    .B1(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__o311a_2 _23242_ (.A1(io_fetch_address[19]),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07675_),
    .C1(_07535_),
    .X(_01413_));
 sky130_fd_sc_hd__a41o_2 _23243_ (.A1(io_fetch_address[19]),
    .A2(io_fetch_address[18]),
    .A3(_06887_),
    .A4(_07613_),
    .B1(io_fetch_address[20]),
    .X(_07676_));
 sky130_fd_sc_hd__nand2_2 _23244_ (.A(io_fetch_address[20]),
    .B(_07651_),
    .Y(_07677_));
 sky130_fd_sc_hd__mux4_2 _23245_ (.A0(\fetch.bht.bhtTable_target_pc[4][20] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][20] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][20] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][20] ),
    .S0(_07068_),
    .S1(_07656_),
    .X(_07678_));
 sky130_fd_sc_hd__mux4_2 _23246_ (.A0(\fetch.bht.bhtTable_target_pc[0][20] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][20] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][20] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][20] ),
    .S0(_07669_),
    .S1(_07100_),
    .X(_07679_));
 sky130_fd_sc_hd__mux4_2 _23247_ (.A0(\fetch.bht.bhtTable_target_pc[12][20] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][20] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][20] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][20] ),
    .S0(_07669_),
    .S1(_07100_),
    .X(_07680_));
 sky130_fd_sc_hd__mux4_2 _23248_ (.A0(\fetch.bht.bhtTable_target_pc[8][20] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][20] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][20] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][20] ),
    .S0(_07669_),
    .S1(_07656_),
    .X(_07681_));
 sky130_fd_sc_hd__mux4_2 _23249_ (.A0(_07678_),
    .A1(_07679_),
    .A2(_07680_),
    .A3(_07681_),
    .S0(_07081_),
    .S1(_06740_),
    .X(_07682_));
 sky130_fd_sc_hd__a211o_2 _23250_ (.A1(\execute.io_target_pc[20] ),
    .A2(_10757_),
    .B1(_10970_),
    .C1(_06037_),
    .X(_07683_));
 sky130_fd_sc_hd__a21o_2 _23251_ (.A1(_07088_),
    .A2(_07682_),
    .B1(_07683_),
    .X(_07684_));
 sky130_fd_sc_hd__a31o_2 _23252_ (.A1(_07064_),
    .A2(_07676_),
    .A3(_07677_),
    .B1(_07684_),
    .X(_07685_));
 sky130_fd_sc_hd__o221a_2 _23253_ (.A1(\csr._csr_read_data_T_8[20] ),
    .A2(_06480_),
    .B1(\csr.io_mret_vector[20] ),
    .B2(_07621_),
    .C1(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__a31o_2 _23254_ (.A1(_07619_),
    .A2(_07573_),
    .A3(_07620_),
    .B1(_07686_),
    .X(_07687_));
 sky130_fd_sc_hd__o311a_2 _23255_ (.A1(io_fetch_address[20]),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07687_),
    .C1(_07535_),
    .X(_01414_));
 sky130_fd_sc_hd__o22a_2 _23256_ (.A1(\csr._csr_read_data_T_8[21] ),
    .A2(_06480_),
    .B1(\csr.io_mret_vector[21] ),
    .B2(_07621_),
    .X(_07688_));
 sky130_fd_sc_hd__a31o_2 _23257_ (.A1(io_fetch_address[20]),
    .A2(io_fetch_address[19]),
    .A3(_07636_),
    .B1(io_fetch_address[21]),
    .X(_07689_));
 sky130_fd_sc_hd__nand4_2 _23258_ (.A(io_fetch_address[21]),
    .B(io_fetch_address[20]),
    .C(io_fetch_address[19]),
    .D(_07636_),
    .Y(_07690_));
 sky130_fd_sc_hd__mux4_2 _23259_ (.A0(\fetch.bht.bhtTable_target_pc[0][21] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][21] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][21] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][21] ),
    .S0(_07119_),
    .S1(_07071_),
    .X(_07691_));
 sky130_fd_sc_hd__nor2_2 _23260_ (.A(_07122_),
    .B(_07691_),
    .Y(_07692_));
 sky130_fd_sc_hd__mux2_2 _23261_ (.A0(\fetch.bht.bhtTable_target_pc[4][21] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][21] ),
    .S(_07106_),
    .X(_07693_));
 sky130_fd_sc_hd__or2b_2 _23262_ (.A(_07110_),
    .B_N(_07693_),
    .X(_07694_));
 sky130_fd_sc_hd__mux2_2 _23263_ (.A0(\fetch.bht.bhtTable_target_pc[6][21] ),
    .A1(\fetch.bht.bhtTable_target_pc[7][21] ),
    .S(_07068_),
    .X(_07695_));
 sky130_fd_sc_hd__nand2_2 _23264_ (.A(_07695_),
    .B(_07114_),
    .Y(_07696_));
 sky130_fd_sc_hd__a31o_2 _23265_ (.A1(_07694_),
    .A2(_07075_),
    .A3(_07696_),
    .B1(_06740_),
    .X(_07697_));
 sky130_fd_sc_hd__mux4_2 _23266_ (.A0(\fetch.bht.bhtTable_target_pc[12][21] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][21] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][21] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][21] ),
    .S0(_07098_),
    .S1(_07113_),
    .X(_07698_));
 sky130_fd_sc_hd__mux4_2 _23267_ (.A0(\fetch.bht.bhtTable_target_pc[8][21] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][21] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][21] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][21] ),
    .S0(_07098_),
    .S1(_07113_),
    .X(_07699_));
 sky130_fd_sc_hd__mux2_2 _23268_ (.A0(_07698_),
    .A1(_07699_),
    .S(_07081_),
    .X(_07700_));
 sky130_fd_sc_hd__a2bb2o_2 _23269_ (.A1_N(_07692_),
    .A2_N(_07697_),
    .B1(_07127_),
    .B2(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__a221o_2 _23270_ (.A1(\execute.io_target_pc[21] ),
    .A2(_07090_),
    .B1(_07089_),
    .B2(_07701_),
    .C1(_06032_),
    .X(_07702_));
 sky130_fd_sc_hd__a31o_2 _23271_ (.A1(_07064_),
    .A2(_07689_),
    .A3(_07690_),
    .B1(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__a2bb2o_2 _23272_ (.A1_N(_06248_),
    .A2_N(_10915_),
    .B1(_07688_),
    .B2(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__buf_1 _23273_ (.A(_09956_),
    .X(_07705_));
 sky130_fd_sc_hd__o311a_2 _23274_ (.A1(io_fetch_address[21]),
    .A2(_07536_),
    .A3(_07537_),
    .B1(_07704_),
    .C1(_07705_),
    .X(_01415_));
 sky130_fd_sc_hd__buf_1 _23275_ (.A(_06248_),
    .X(_07706_));
 sky130_fd_sc_hd__buf_1 _23276_ (.A(_03500_),
    .X(_07707_));
 sky130_fd_sc_hd__buf_1 _23277_ (.A(_07098_),
    .X(_07708_));
 sky130_fd_sc_hd__mux4_2 _23278_ (.A0(\fetch.bht.bhtTable_target_pc[8][22] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][22] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][22] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][22] ),
    .S0(_07708_),
    .S1(_07103_),
    .X(_07709_));
 sky130_fd_sc_hd__buf_1 _23279_ (.A(_07100_),
    .X(_07710_));
 sky130_fd_sc_hd__mux4_2 _23280_ (.A0(\fetch.bht.bhtTable_target_pc[12][22] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][22] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][22] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][22] ),
    .S0(_07555_),
    .S1(_07710_),
    .X(_07711_));
 sky130_fd_sc_hd__mux4_2 _23281_ (.A0(\fetch.bht.bhtTable_target_pc[0][22] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][22] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][22] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][22] ),
    .S0(_07708_),
    .S1(_07710_),
    .X(_07712_));
 sky130_fd_sc_hd__mux4_2 _23282_ (.A0(\fetch.bht.bhtTable_target_pc[4][22] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][22] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][22] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][22] ),
    .S0(_07708_),
    .S1(_07103_),
    .X(_07713_));
 sky130_fd_sc_hd__mux4_2 _23283_ (.A0(_07709_),
    .A1(_07711_),
    .A2(_07712_),
    .A3(_07713_),
    .S0(_07122_),
    .S1(_07084_),
    .X(_07714_));
 sky130_fd_sc_hd__a211o_2 _23284_ (.A1(\execute.io_target_pc[22] ),
    .A2(_07090_),
    .B1(_06041_),
    .C1(_06038_),
    .X(_07715_));
 sky130_fd_sc_hd__and3_2 _23285_ (.A(io_fetch_address[21]),
    .B(io_fetch_address[20]),
    .C(_07651_),
    .X(_07716_));
 sky130_fd_sc_hd__nand2_2 _23286_ (.A(io_fetch_address[22]),
    .B(_07716_),
    .Y(_07717_));
 sky130_fd_sc_hd__o211a_2 _23287_ (.A1(io_fetch_address[22]),
    .A2(_07716_),
    .B1(_07717_),
    .C1(_07064_),
    .X(_07718_));
 sky130_fd_sc_hd__a211o_2 _23288_ (.A1(_07089_),
    .A2(_07714_),
    .B1(_07715_),
    .C1(_07718_),
    .X(_07719_));
 sky130_fd_sc_hd__o221a_2 _23289_ (.A1(\csr._csr_read_data_T_8[22] ),
    .A2(_07416_),
    .B1(\csr.io_mret_vector[22] ),
    .B2(_07621_),
    .C1(_07719_),
    .X(_07720_));
 sky130_fd_sc_hd__a31o_2 _23290_ (.A1(_07619_),
    .A2(_07573_),
    .A3(_07620_),
    .B1(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__o311a_2 _23291_ (.A1(io_fetch_address[22]),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07721_),
    .C1(_07705_),
    .X(_01416_));
 sky130_fd_sc_hd__mux4_2 _23292_ (.A0(\fetch.bht.bhtTable_target_pc[4][23] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][23] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][23] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][23] ),
    .S0(_07708_),
    .S1(_07103_),
    .X(_07722_));
 sky130_fd_sc_hd__mux4_2 _23293_ (.A0(\fetch.bht.bhtTable_target_pc[0][23] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][23] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][23] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][23] ),
    .S0(_07555_),
    .S1(_07710_),
    .X(_07723_));
 sky130_fd_sc_hd__mux4_2 _23294_ (.A0(\fetch.bht.bhtTable_target_pc[12][23] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][23] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][23] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][23] ),
    .S0(_07708_),
    .S1(_07710_),
    .X(_07724_));
 sky130_fd_sc_hd__mux4_2 _23295_ (.A0(\fetch.bht.bhtTable_target_pc[8][23] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][23] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][23] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][23] ),
    .S0(_07708_),
    .S1(_07103_),
    .X(_07725_));
 sky130_fd_sc_hd__mux4_2 _23296_ (.A0(_07722_),
    .A1(_07723_),
    .A2(_07724_),
    .A3(_07725_),
    .S0(_07371_),
    .S1(_07127_),
    .X(_07726_));
 sky130_fd_sc_hd__a211o_2 _23297_ (.A1(\execute.io_target_pc[23] ),
    .A2(_07090_),
    .B1(_06041_),
    .C1(_06038_),
    .X(_07727_));
 sky130_fd_sc_hd__and3_2 _23298_ (.A(io_fetch_address[23]),
    .B(io_fetch_address[22]),
    .C(_07716_),
    .X(_07728_));
 sky130_fd_sc_hd__a41o_2 _23299_ (.A1(io_fetch_address[22]),
    .A2(io_fetch_address[21]),
    .A3(io_fetch_address[20]),
    .A4(_07651_),
    .B1(io_fetch_address[23]),
    .X(_07729_));
 sky130_fd_sc_hd__and3b_2 _23300_ (.A_N(_07728_),
    .B(_07729_),
    .C(_07063_),
    .X(_07730_));
 sky130_fd_sc_hd__a211o_2 _23301_ (.A1(_07089_),
    .A2(_07726_),
    .B1(_07727_),
    .C1(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__o221a_2 _23302_ (.A1(\csr._csr_read_data_T_8[23] ),
    .A2(_07416_),
    .B1(\csr.io_mret_vector[23] ),
    .B2(_07621_),
    .C1(_07731_),
    .X(_07732_));
 sky130_fd_sc_hd__a31o_2 _23303_ (.A1(_07619_),
    .A2(_07573_),
    .A3(_07620_),
    .B1(_07732_),
    .X(_07733_));
 sky130_fd_sc_hd__o311a_2 _23304_ (.A1(io_fetch_address[23]),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07733_),
    .C1(_07705_),
    .X(_01417_));
 sky130_fd_sc_hd__mux4_2 _23305_ (.A0(\fetch.bht.bhtTable_target_pc[4][24] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][24] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][24] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][24] ),
    .S0(_07708_),
    .S1(_07103_),
    .X(_07734_));
 sky130_fd_sc_hd__mux4_2 _23306_ (.A0(\fetch.bht.bhtTable_target_pc[0][24] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][24] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][24] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][24] ),
    .S0(_07555_),
    .S1(_07710_),
    .X(_07735_));
 sky130_fd_sc_hd__mux4_2 _23307_ (.A0(\fetch.bht.bhtTable_target_pc[12][24] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][24] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][24] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][24] ),
    .S0(_07555_),
    .S1(_07710_),
    .X(_07736_));
 sky130_fd_sc_hd__mux4_2 _23308_ (.A0(\fetch.bht.bhtTable_target_pc[8][24] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][24] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][24] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][24] ),
    .S0(_07708_),
    .S1(_07710_),
    .X(_07737_));
 sky130_fd_sc_hd__mux4_2 _23309_ (.A0(_07734_),
    .A1(_07735_),
    .A2(_07736_),
    .A3(_07737_),
    .S0(_07371_),
    .S1(_07127_),
    .X(_07738_));
 sky130_fd_sc_hd__a211o_2 _23310_ (.A1(\execute.io_target_pc[24] ),
    .A2(_07090_),
    .B1(_06041_),
    .C1(_06037_),
    .X(_07739_));
 sky130_fd_sc_hd__and4_2 _23311_ (.A(io_fetch_address[24]),
    .B(io_fetch_address[23]),
    .C(io_fetch_address[22]),
    .D(_07716_),
    .X(_07740_));
 sky130_fd_sc_hd__a31o_2 _23312_ (.A1(io_fetch_address[23]),
    .A2(io_fetch_address[22]),
    .A3(_07716_),
    .B1(io_fetch_address[24]),
    .X(_07741_));
 sky130_fd_sc_hd__and3b_2 _23313_ (.A_N(_07740_),
    .B(_07063_),
    .C(_07741_),
    .X(_07742_));
 sky130_fd_sc_hd__a211o_2 _23314_ (.A1(_07089_),
    .A2(_07738_),
    .B1(_07739_),
    .C1(_07742_),
    .X(_07743_));
 sky130_fd_sc_hd__o221a_2 _23315_ (.A1(\csr._csr_read_data_T_8[24] ),
    .A2(_07416_),
    .B1(\csr.io_mret_vector[24] ),
    .B2(_07621_),
    .C1(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__a31o_2 _23316_ (.A1(_07619_),
    .A2(_07573_),
    .A3(_07620_),
    .B1(_07744_),
    .X(_07745_));
 sky130_fd_sc_hd__o311a_2 _23317_ (.A1(io_fetch_address[24]),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07745_),
    .C1(_07705_),
    .X(_01418_));
 sky130_fd_sc_hd__o22a_2 _23318_ (.A1(\csr._csr_read_data_T_8[25] ),
    .A2(_06480_),
    .B1(\csr.io_mret_vector[25] ),
    .B2(_07621_),
    .X(_07746_));
 sky130_fd_sc_hd__nand2_2 _23319_ (.A(io_fetch_address[25]),
    .B(_07740_),
    .Y(_07747_));
 sky130_fd_sc_hd__a41o_2 _23320_ (.A1(io_fetch_address[24]),
    .A2(io_fetch_address[23]),
    .A3(io_fetch_address[22]),
    .A4(_07716_),
    .B1(io_fetch_address[25]),
    .X(_07748_));
 sky130_fd_sc_hd__mux4_2 _23321_ (.A0(\fetch.bht.bhtTable_target_pc[12][25] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][25] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][25] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][25] ),
    .S0(_07384_),
    .S1(_07386_),
    .X(_07749_));
 sky130_fd_sc_hd__mux4_2 _23322_ (.A0(\fetch.bht.bhtTable_target_pc[8][25] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][25] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][25] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][25] ),
    .S0(_07384_),
    .S1(_07386_),
    .X(_07750_));
 sky130_fd_sc_hd__mux2_2 _23323_ (.A0(_07749_),
    .A1(_07750_),
    .S(_07081_),
    .X(_07751_));
 sky130_fd_sc_hd__mux4_2 _23324_ (.A0(\fetch.bht.bhtTable_target_pc[0][25] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][25] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][25] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][25] ),
    .S0(_07098_),
    .S1(_07113_),
    .X(_07752_));
 sky130_fd_sc_hd__mux2_2 _23325_ (.A0(\fetch.bht.bhtTable_target_pc[4][25] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][25] ),
    .S(_07067_),
    .X(_07753_));
 sky130_fd_sc_hd__and2b_2 _23326_ (.A_N(_07110_),
    .B(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__mux2_2 _23327_ (.A0(\fetch.bht.bhtTable_target_pc[6][25] ),
    .A1(\fetch.bht.bhtTable_target_pc[7][25] ),
    .S(_07106_),
    .X(_07755_));
 sky130_fd_sc_hd__a21o_2 _23328_ (.A1(_07755_),
    .A2(_07071_),
    .B1(_07080_),
    .X(_07756_));
 sky130_fd_sc_hd__o22a_2 _23329_ (.A1(_07075_),
    .A2(_07752_),
    .B1(_07754_),
    .B2(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__mux2_2 _23330_ (.A0(_07751_),
    .A1(_07757_),
    .S(_07084_),
    .X(_07758_));
 sky130_fd_sc_hd__a221o_2 _23331_ (.A1(\execute.io_target_pc[25] ),
    .A2(_07090_),
    .B1(_07089_),
    .B2(_07758_),
    .C1(_06032_),
    .X(_07759_));
 sky130_fd_sc_hd__a31o_2 _23332_ (.A1(_07064_),
    .A2(_07747_),
    .A3(_07748_),
    .B1(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__a2bb2o_2 _23333_ (.A1_N(_06248_),
    .A2_N(_10915_),
    .B1(_07746_),
    .B2(_07760_),
    .X(_07761_));
 sky130_fd_sc_hd__o311a_2 _23334_ (.A1(io_fetch_address[25]),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07761_),
    .C1(_07705_),
    .X(_01419_));
 sky130_fd_sc_hd__mux4_2 _23335_ (.A0(\fetch.bht.bhtTable_target_pc[8][26] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][26] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][26] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][26] ),
    .S0(_07068_),
    .S1(_07656_),
    .X(_07762_));
 sky130_fd_sc_hd__mux4_2 _23336_ (.A0(\fetch.bht.bhtTable_target_pc[12][26] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][26] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][26] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][26] ),
    .S0(_07669_),
    .S1(_07656_),
    .X(_07763_));
 sky130_fd_sc_hd__mux2_2 _23337_ (.A0(_07762_),
    .A1(_07763_),
    .S(_07075_),
    .X(_07764_));
 sky130_fd_sc_hd__mux4_2 _23338_ (.A0(\fetch.bht.bhtTable_target_pc[4][26] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][26] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][26] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][26] ),
    .S0(_07669_),
    .S1(_07656_),
    .X(_07765_));
 sky130_fd_sc_hd__mux4_2 _23339_ (.A0(\fetch.bht.bhtTable_target_pc[0][26] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][26] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][26] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][26] ),
    .S0(_07669_),
    .S1(_07656_),
    .X(_07766_));
 sky130_fd_sc_hd__mux2_2 _23340_ (.A0(_07765_),
    .A1(_07766_),
    .S(_07081_),
    .X(_07767_));
 sky130_fd_sc_hd__mux2_2 _23341_ (.A0(_07764_),
    .A1(_07767_),
    .S(_07084_),
    .X(_07768_));
 sky130_fd_sc_hd__a211o_2 _23342_ (.A1(\execute.io_target_pc[26] ),
    .A2(_07090_),
    .B1(_10970_),
    .C1(_06037_),
    .X(_07769_));
 sky130_fd_sc_hd__nand4_2 _23343_ (.A(io_fetch_address[26]),
    .B(io_fetch_address[25]),
    .C(io_fetch_address[24]),
    .D(_07728_),
    .Y(_07770_));
 sky130_fd_sc_hd__a31o_2 _23344_ (.A1(io_fetch_address[25]),
    .A2(io_fetch_address[24]),
    .A3(_07728_),
    .B1(io_fetch_address[26]),
    .X(_07771_));
 sky130_fd_sc_hd__and3_2 _23345_ (.A(_07064_),
    .B(_07770_),
    .C(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__a211o_2 _23346_ (.A1(_07089_),
    .A2(_07768_),
    .B1(_07769_),
    .C1(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__o221a_2 _23347_ (.A1(\csr._csr_read_data_T_8[26] ),
    .A2(_07416_),
    .B1(\csr.io_mret_vector[26] ),
    .B2(_07621_),
    .C1(_07773_),
    .X(_07774_));
 sky130_fd_sc_hd__a31o_2 _23348_ (.A1(_07619_),
    .A2(_07573_),
    .A3(_07620_),
    .B1(_07774_),
    .X(_07775_));
 sky130_fd_sc_hd__o311a_2 _23349_ (.A1(io_fetch_address[26]),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07775_),
    .C1(_07705_),
    .X(_01420_));
 sky130_fd_sc_hd__mux4_2 _23350_ (.A0(\fetch.bht.bhtTable_target_pc[12][27] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][27] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][27] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][27] ),
    .S0(_07708_),
    .S1(_07103_),
    .X(_07776_));
 sky130_fd_sc_hd__mux4_2 _23351_ (.A0(\fetch.bht.bhtTable_target_pc[8][27] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][27] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][27] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][27] ),
    .S0(_07555_),
    .S1(_07710_),
    .X(_07777_));
 sky130_fd_sc_hd__mux4_2 _23352_ (.A0(\fetch.bht.bhtTable_target_pc[4][27] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][27] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][27] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][27] ),
    .S0(_07555_),
    .S1(_07710_),
    .X(_07778_));
 sky130_fd_sc_hd__mux4_2 _23353_ (.A0(\fetch.bht.bhtTable_target_pc[0][27] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][27] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][27] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][27] ),
    .S0(_07708_),
    .S1(_07710_),
    .X(_07779_));
 sky130_fd_sc_hd__mux4_2 _23354_ (.A0(_07776_),
    .A1(_07777_),
    .A2(_07778_),
    .A3(_07779_),
    .S0(_07371_),
    .S1(_07084_),
    .X(_07780_));
 sky130_fd_sc_hd__a211o_2 _23355_ (.A1(\execute.io_target_pc[27] ),
    .A2(_10757_),
    .B1(_10970_),
    .C1(_06037_),
    .X(_07781_));
 sky130_fd_sc_hd__and4_2 _23356_ (.A(io_fetch_address[27]),
    .B(io_fetch_address[26]),
    .C(io_fetch_address[25]),
    .D(_07740_),
    .X(_07782_));
 sky130_fd_sc_hd__buf_1 _23357_ (.A(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__a31o_2 _23358_ (.A1(io_fetch_address[26]),
    .A2(io_fetch_address[25]),
    .A3(_07740_),
    .B1(io_fetch_address[27]),
    .X(_07784_));
 sky130_fd_sc_hd__and3b_2 _23359_ (.A_N(_07783_),
    .B(_07784_),
    .C(_07063_),
    .X(_07785_));
 sky130_fd_sc_hd__a211o_2 _23360_ (.A1(_07089_),
    .A2(_07780_),
    .B1(_07781_),
    .C1(_07785_),
    .X(_07786_));
 sky130_fd_sc_hd__o221a_2 _23361_ (.A1(\csr._csr_read_data_T_8[27] ),
    .A2(_07416_),
    .B1(\csr.io_mret_vector[27] ),
    .B2(_07621_),
    .C1(_07786_),
    .X(_07787_));
 sky130_fd_sc_hd__a31o_2 _23362_ (.A1(_07619_),
    .A2(_07573_),
    .A3(_07620_),
    .B1(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__o311a_2 _23363_ (.A1(io_fetch_address[27]),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07788_),
    .C1(_07705_),
    .X(_01421_));
 sky130_fd_sc_hd__nand2_2 _23364_ (.A(_06795_),
    .B(_07783_),
    .Y(_07789_));
 sky130_fd_sc_hd__o211a_2 _23365_ (.A1(_06795_),
    .A2(_07783_),
    .B1(_07789_),
    .C1(_07064_),
    .X(_07790_));
 sky130_fd_sc_hd__mux4_2 _23366_ (.A0(\fetch.bht.bhtTable_target_pc[8][28] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][28] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][28] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][28] ),
    .S0(_07119_),
    .S1(_07071_),
    .X(_07791_));
 sky130_fd_sc_hd__o21ai_2 _23367_ (.A1(_07075_),
    .A2(_07791_),
    .B1(_06740_),
    .Y(_07792_));
 sky130_fd_sc_hd__or2b_2 _23368_ (.A(\fetch.bht.bhtTable_target_pc[13][28] ),
    .B_N(_07099_),
    .X(_07793_));
 sky130_fd_sc_hd__o21ba_2 _23369_ (.A1(_07099_),
    .A2(\fetch.bht.bhtTable_target_pc[12][28] ),
    .B1_N(_07071_),
    .X(_07794_));
 sky130_fd_sc_hd__mux2_2 _23370_ (.A0(\fetch.bht.bhtTable_target_pc[14][28] ),
    .A1(\fetch.bht.bhtTable_target_pc[15][28] ),
    .S(_07107_),
    .X(_07795_));
 sky130_fd_sc_hd__a221oi_2 _23371_ (.A1(_07793_),
    .A2(_07794_),
    .B1(_07795_),
    .B2(_07072_),
    .C1(_07371_),
    .Y(_07796_));
 sky130_fd_sc_hd__mux4_2 _23372_ (.A0(\fetch.bht.bhtTable_target_pc[4][28] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][28] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][28] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][28] ),
    .S0(_07384_),
    .S1(_07386_),
    .X(_07797_));
 sky130_fd_sc_hd__mux4_2 _23373_ (.A0(\fetch.bht.bhtTable_target_pc[0][28] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][28] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][28] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][28] ),
    .S0(_07384_),
    .S1(_07386_),
    .X(_07798_));
 sky130_fd_sc_hd__mux2_2 _23374_ (.A0(_07797_),
    .A1(_07798_),
    .S(_07081_),
    .X(_07799_));
 sky130_fd_sc_hd__a2bb2o_2 _23375_ (.A1_N(_07792_),
    .A2_N(_07796_),
    .B1(_07084_),
    .B2(_07799_),
    .X(_07800_));
 sky130_fd_sc_hd__a221o_2 _23376_ (.A1(\execute.io_target_pc[28] ),
    .A2(_07090_),
    .B1(_07089_),
    .B2(_07800_),
    .C1(_06032_),
    .X(_07801_));
 sky130_fd_sc_hd__or3b_2 _23377_ (.A(_06038_),
    .B(\csr.io_mret_vector[28] ),
    .C_N(_06041_),
    .X(_07802_));
 sky130_fd_sc_hd__o221a_2 _23378_ (.A1(\csr._csr_read_data_T_8[28] ),
    .A2(_07416_),
    .B1(_07790_),
    .B2(_07801_),
    .C1(_07802_),
    .X(_07803_));
 sky130_fd_sc_hd__a31o_2 _23379_ (.A1(_07619_),
    .A2(_07345_),
    .A3(_07620_),
    .B1(_07803_),
    .X(_07804_));
 sky130_fd_sc_hd__o311a_2 _23380_ (.A1(_06795_),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07804_),
    .C1(_07705_),
    .X(_01422_));
 sky130_fd_sc_hd__mux4_2 _23381_ (.A0(\fetch.bht.bhtTable_target_pc[12][29] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][29] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][29] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][29] ),
    .S0(_07068_),
    .S1(_07656_),
    .X(_07805_));
 sky130_fd_sc_hd__mux4_2 _23382_ (.A0(\fetch.bht.bhtTable_target_pc[8][29] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][29] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][29] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][29] ),
    .S0(_07669_),
    .S1(_07656_),
    .X(_07806_));
 sky130_fd_sc_hd__mux2_2 _23383_ (.A0(_07805_),
    .A1(_07806_),
    .S(_07081_),
    .X(_07807_));
 sky130_fd_sc_hd__mux4_2 _23384_ (.A0(\fetch.bht.bhtTable_target_pc[4][29] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][29] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][29] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][29] ),
    .S0(_07669_),
    .S1(_07656_),
    .X(_07808_));
 sky130_fd_sc_hd__mux4_2 _23385_ (.A0(\fetch.bht.bhtTable_target_pc[0][29] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][29] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][29] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][29] ),
    .S0(_07669_),
    .S1(_07100_),
    .X(_07809_));
 sky130_fd_sc_hd__mux2_2 _23386_ (.A0(_07808_),
    .A1(_07809_),
    .S(_07081_),
    .X(_07810_));
 sky130_fd_sc_hd__mux2_2 _23387_ (.A0(_07807_),
    .A1(_07810_),
    .S(_07084_),
    .X(_07811_));
 sky130_fd_sc_hd__a211o_2 _23388_ (.A1(\execute.io_target_pc[29] ),
    .A2(_10757_),
    .B1(_10970_),
    .C1(_06037_),
    .X(_07812_));
 sky130_fd_sc_hd__nand3_2 _23389_ (.A(io_fetch_address[29]),
    .B(_06795_),
    .C(_07783_),
    .Y(_07813_));
 sky130_fd_sc_hd__a21o_2 _23390_ (.A1(_06795_),
    .A2(_07783_),
    .B1(io_fetch_address[29]),
    .X(_07814_));
 sky130_fd_sc_hd__and3_2 _23391_ (.A(_07064_),
    .B(_07813_),
    .C(_07814_),
    .X(_07815_));
 sky130_fd_sc_hd__a211o_2 _23392_ (.A1(_07089_),
    .A2(_07811_),
    .B1(_07812_),
    .C1(_07815_),
    .X(_07816_));
 sky130_fd_sc_hd__o221a_2 _23393_ (.A1(\csr._csr_read_data_T_8[29] ),
    .A2(_07416_),
    .B1(\csr.io_mret_vector[29] ),
    .B2(_07417_),
    .C1(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__a31o_2 _23394_ (.A1(_07619_),
    .A2(_07345_),
    .A3(_07620_),
    .B1(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__o311a_2 _23395_ (.A1(io_fetch_address[29]),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07818_),
    .C1(_07705_),
    .X(_01423_));
 sky130_fd_sc_hd__nand4_2 _23396_ (.A(io_fetch_address[30]),
    .B(io_fetch_address[29]),
    .C(_06795_),
    .D(_07783_),
    .Y(_07819_));
 sky130_fd_sc_hd__a31o_2 _23397_ (.A1(io_fetch_address[29]),
    .A2(_06795_),
    .A3(_07783_),
    .B1(io_fetch_address[30]),
    .X(_07820_));
 sky130_fd_sc_hd__mux4_2 _23398_ (.A0(\fetch.bht.bhtTable_target_pc[12][30] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][30] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][30] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][30] ),
    .S0(_07106_),
    .S1(_07386_),
    .X(_07821_));
 sky130_fd_sc_hd__mux4_2 _23399_ (.A0(\fetch.bht.bhtTable_target_pc[8][30] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][30] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][30] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][30] ),
    .S0(_07106_),
    .S1(_07070_),
    .X(_07822_));
 sky130_fd_sc_hd__mux4_2 _23400_ (.A0(\fetch.bht.bhtTable_target_pc[4][30] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][30] ),
    .A2(\fetch.bht.bhtTable_target_pc[6][30] ),
    .A3(\fetch.bht.bhtTable_target_pc[7][30] ),
    .S0(_07106_),
    .S1(_07070_),
    .X(_07823_));
 sky130_fd_sc_hd__mux4_2 _23401_ (.A0(\fetch.bht.bhtTable_target_pc[0][30] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][30] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][30] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][30] ),
    .S0(_07106_),
    .S1(_07386_),
    .X(_07824_));
 sky130_fd_sc_hd__mux4_2 _23402_ (.A0(_07821_),
    .A1(_07822_),
    .A2(_07823_),
    .A3(_07824_),
    .S0(_07080_),
    .S1(_06637_),
    .X(_07825_));
 sky130_fd_sc_hd__a221o_2 _23403_ (.A1(\execute.io_target_pc[30] ),
    .A2(_10757_),
    .B1(_07088_),
    .B2(_07825_),
    .C1(_10971_),
    .X(_07826_));
 sky130_fd_sc_hd__a31o_2 _23404_ (.A1(_07064_),
    .A2(_07819_),
    .A3(_07820_),
    .B1(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__o221a_2 _23405_ (.A1(\csr._csr_read_data_T_8[30] ),
    .A2(_07416_),
    .B1(\csr.io_mret_vector[30] ),
    .B2(_07417_),
    .C1(_07827_),
    .X(_07828_));
 sky130_fd_sc_hd__a31o_2 _23406_ (.A1(_05857_),
    .A2(_07345_),
    .A3(_10672_),
    .B1(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__o311a_2 _23407_ (.A1(io_fetch_address[30]),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07829_),
    .C1(_07705_),
    .X(_01424_));
 sky130_fd_sc_hd__o21ai_2 _23408_ (.A1(io_fetch_address[31]),
    .A2(_07819_),
    .B1(_07087_),
    .Y(_07830_));
 sky130_fd_sc_hd__a21o_2 _23409_ (.A1(io_fetch_address[31]),
    .A2(_07819_),
    .B1(_07830_),
    .X(_07831_));
 sky130_fd_sc_hd__mux4_2 _23410_ (.A0(\fetch.bht.bhtTable_target_pc[12][31] ),
    .A1(\fetch.bht.bhtTable_target_pc[13][31] ),
    .A2(\fetch.bht.bhtTable_target_pc[14][31] ),
    .A3(\fetch.bht.bhtTable_target_pc[15][31] ),
    .S0(_07066_),
    .S1(_07070_),
    .X(_07832_));
 sky130_fd_sc_hd__mux4_2 _23411_ (.A0(\fetch.bht.bhtTable_target_pc[8][31] ),
    .A1(\fetch.bht.bhtTable_target_pc[9][31] ),
    .A2(\fetch.bht.bhtTable_target_pc[10][31] ),
    .A3(\fetch.bht.bhtTable_target_pc[11][31] ),
    .S0(_07066_),
    .S1(_06661_),
    .X(_07833_));
 sky130_fd_sc_hd__mux2_2 _23412_ (.A0(_07832_),
    .A1(_07833_),
    .S(_07080_),
    .X(_07834_));
 sky130_fd_sc_hd__mux4_2 _23413_ (.A0(\fetch.bht.bhtTable_target_pc[0][31] ),
    .A1(\fetch.bht.bhtTable_target_pc[1][31] ),
    .A2(\fetch.bht.bhtTable_target_pc[2][31] ),
    .A3(\fetch.bht.bhtTable_target_pc[3][31] ),
    .S0(_07066_),
    .S1(_07070_),
    .X(_07835_));
 sky130_fd_sc_hd__mux2_2 _23414_ (.A0(\fetch.bht.bhtTable_target_pc[4][31] ),
    .A1(\fetch.bht.bhtTable_target_pc[5][31] ),
    .S(_07066_),
    .X(_07836_));
 sky130_fd_sc_hd__and2b_2 _23415_ (.A_N(_07070_),
    .B(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__mux2_2 _23416_ (.A0(\fetch.bht.bhtTable_target_pc[6][31] ),
    .A1(\fetch.bht.bhtTable_target_pc[7][31] ),
    .S(_07066_),
    .X(_07838_));
 sky130_fd_sc_hd__a21o_2 _23417_ (.A1(_07838_),
    .A2(_07070_),
    .B1(_07080_),
    .X(_07839_));
 sky130_fd_sc_hd__o22a_2 _23418_ (.A1(_06633_),
    .A2(_07835_),
    .B1(_07837_),
    .B2(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__mux2_2 _23419_ (.A0(_07834_),
    .A1(_07840_),
    .S(_06637_),
    .X(_07841_));
 sky130_fd_sc_hd__a21o_2 _23420_ (.A1(_03592_),
    .A2(_07841_),
    .B1(_07064_),
    .X(_07842_));
 sky130_fd_sc_hd__a221o_2 _23421_ (.A1(\execute.io_target_pc[31] ),
    .A2(_07091_),
    .B1(_07831_),
    .B2(_07842_),
    .C1(_06032_),
    .X(_07843_));
 sky130_fd_sc_hd__o221a_2 _23422_ (.A1(\csr._csr_read_data_T_8[31] ),
    .A2(_07416_),
    .B1(\csr.io_mret_vector[31] ),
    .B2(_07417_),
    .C1(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__a31o_2 _23423_ (.A1(_05857_),
    .A2(_07345_),
    .A3(_10672_),
    .B1(_07844_),
    .X(_07845_));
 sky130_fd_sc_hd__o311a_2 _23424_ (.A1(io_fetch_address[31]),
    .A2(_07706_),
    .A3(_07707_),
    .B1(_07845_),
    .C1(_05856_),
    .X(_01425_));
 sky130_fd_sc_hd__buf_1 _23425_ (.A(_03546_),
    .X(_07846_));
 sky130_fd_sc_hd__buf_1 _23426_ (.A(_10670_),
    .X(_07847_));
 sky130_fd_sc_hd__or3b_2 _23427_ (.A(\decode.control.io_opcode[2] ),
    .B(_07847_),
    .C_N(_05206_),
    .X(_07848_));
 sky130_fd_sc_hd__o211a_2 _23428_ (.A1(io_fetch_data[2]),
    .A2(_07846_),
    .B1(_07848_),
    .C1(_05454_),
    .X(_01426_));
 sky130_fd_sc_hd__and4bb_2 _23429_ (.A_N(_06422_),
    .B_N(_10910_),
    .C(_03500_),
    .D(io_fetch_data[3]),
    .X(_07849_));
 sky130_fd_sc_hd__buf_1 _23430_ (.A(_07849_),
    .X(_01427_));
 sky130_fd_sc_hd__or3b_2 _23431_ (.A(_10965_),
    .B(_07847_),
    .C_N(_05206_),
    .X(_07850_));
 sky130_fd_sc_hd__buf_1 _23432_ (.A(_04459_),
    .X(_07851_));
 sky130_fd_sc_hd__o211a_2 _23433_ (.A1(io_fetch_data[5]),
    .A2(_07846_),
    .B1(_07850_),
    .C1(_07851_),
    .X(_01428_));
 sky130_fd_sc_hd__or3b_2 _23434_ (.A(_10579_),
    .B(_07847_),
    .C_N(_05206_),
    .X(_07852_));
 sky130_fd_sc_hd__o211a_2 _23435_ (.A1(io_fetch_data[6]),
    .A2(_07846_),
    .B1(_07852_),
    .C1(_07851_),
    .X(_01429_));
 sky130_fd_sc_hd__or3b_2 _23436_ (.A(\decode.immGen._imm_T_10[0] ),
    .B(_07847_),
    .C_N(_05206_),
    .X(_07853_));
 sky130_fd_sc_hd__o211a_2 _23437_ (.A1(io_fetch_data[7]),
    .A2(_07846_),
    .B1(_07853_),
    .C1(_07851_),
    .X(_01430_));
 sky130_fd_sc_hd__or3b_2 _23438_ (.A(\decode.immGen._imm_T_10[1] ),
    .B(_07847_),
    .C_N(_05206_),
    .X(_07854_));
 sky130_fd_sc_hd__o211a_2 _23439_ (.A1(io_fetch_data[8]),
    .A2(_07846_),
    .B1(_07854_),
    .C1(_07851_),
    .X(_01431_));
 sky130_fd_sc_hd__or3b_2 _23440_ (.A(\decode.immGen._imm_T_10[2] ),
    .B(_07847_),
    .C_N(_05206_),
    .X(_07855_));
 sky130_fd_sc_hd__o211a_2 _23441_ (.A1(io_fetch_data[9]),
    .A2(_07846_),
    .B1(_07855_),
    .C1(_07851_),
    .X(_01432_));
 sky130_fd_sc_hd__or3b_2 _23442_ (.A(\decode.immGen._imm_T_10[3] ),
    .B(_07847_),
    .C_N(_05206_),
    .X(_07856_));
 sky130_fd_sc_hd__o211a_2 _23443_ (.A1(io_fetch_data[10]),
    .A2(_07846_),
    .B1(_07856_),
    .C1(_07851_),
    .X(_01433_));
 sky130_fd_sc_hd__or3b_2 _23444_ (.A(\decode.immGen._imm_T_10[4] ),
    .B(_07847_),
    .C_N(_05206_),
    .X(_07857_));
 sky130_fd_sc_hd__o211a_2 _23445_ (.A1(io_fetch_data[11]),
    .A2(_07846_),
    .B1(_07857_),
    .C1(_07851_),
    .X(_01434_));
 sky130_fd_sc_hd__or3b_2 _23446_ (.A(_10941_),
    .B(_07847_),
    .C_N(_05206_),
    .X(_07858_));
 sky130_fd_sc_hd__o211a_2 _23447_ (.A1(io_fetch_data[12]),
    .A2(_07846_),
    .B1(_07858_),
    .C1(_07851_),
    .X(_01435_));
 sky130_fd_sc_hd__buf_1 _23448_ (.A(\decode.id_ex_memread_reg ),
    .X(_07859_));
 sky130_fd_sc_hd__or3b_2 _23449_ (.A(_10944_),
    .B(_07847_),
    .C_N(_07859_),
    .X(_07860_));
 sky130_fd_sc_hd__o211a_2 _23450_ (.A1(io_fetch_data[13]),
    .A2(_07846_),
    .B1(_07860_),
    .C1(_07851_),
    .X(_01436_));
 sky130_fd_sc_hd__buf_1 _23451_ (.A(_03546_),
    .X(_07861_));
 sky130_fd_sc_hd__buf_1 _23452_ (.A(_10670_),
    .X(_07862_));
 sky130_fd_sc_hd__or3b_2 _23453_ (.A(_10946_),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07863_));
 sky130_fd_sc_hd__o211a_2 _23454_ (.A1(io_fetch_data[14]),
    .A2(_07861_),
    .B1(_07863_),
    .C1(_07851_),
    .X(_01437_));
 sky130_fd_sc_hd__or3b_2 _23455_ (.A(_12765_),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07864_));
 sky130_fd_sc_hd__buf_1 _23456_ (.A(_04459_),
    .X(_07865_));
 sky130_fd_sc_hd__o211a_2 _23457_ (.A1(io_fetch_data[15]),
    .A2(_07861_),
    .B1(_07864_),
    .C1(_07865_),
    .X(_01438_));
 sky130_fd_sc_hd__or3b_2 _23458_ (.A(_11011_),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07866_));
 sky130_fd_sc_hd__o211a_2 _23459_ (.A1(io_fetch_data[16]),
    .A2(_07861_),
    .B1(_07866_),
    .C1(_07865_),
    .X(_01439_));
 sky130_fd_sc_hd__or3b_2 _23460_ (.A(_11012_),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07867_));
 sky130_fd_sc_hd__o211a_2 _23461_ (.A1(io_fetch_data[17]),
    .A2(_07861_),
    .B1(_07867_),
    .C1(_07865_),
    .X(_01440_));
 sky130_fd_sc_hd__or3b_2 _23462_ (.A(_11015_),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07868_));
 sky130_fd_sc_hd__o211a_2 _23463_ (.A1(io_fetch_data[18]),
    .A2(_07861_),
    .B1(_07868_),
    .C1(_07865_),
    .X(_01441_));
 sky130_fd_sc_hd__or3b_2 _23464_ (.A(_11027_),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07869_));
 sky130_fd_sc_hd__o211a_2 _23465_ (.A1(io_fetch_data[19]),
    .A2(_07861_),
    .B1(_07869_),
    .C1(_07865_),
    .X(_01442_));
 sky130_fd_sc_hd__or3b_2 _23466_ (.A(_10962_),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07870_));
 sky130_fd_sc_hd__o211a_2 _23467_ (.A1(io_fetch_data[20]),
    .A2(_07861_),
    .B1(_07870_),
    .C1(_07865_),
    .X(_01443_));
 sky130_fd_sc_hd__or3b_2 _23468_ (.A(_10981_),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07871_));
 sky130_fd_sc_hd__o211a_2 _23469_ (.A1(io_fetch_data[21]),
    .A2(_07861_),
    .B1(_07871_),
    .C1(_07865_),
    .X(_01444_));
 sky130_fd_sc_hd__or3b_2 _23470_ (.A(_10657_),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07872_));
 sky130_fd_sc_hd__o211a_2 _23471_ (.A1(io_fetch_data[22]),
    .A2(_07861_),
    .B1(_07872_),
    .C1(_07865_),
    .X(_01445_));
 sky130_fd_sc_hd__buf_1 _23472_ (.A(\decode.id_ex_memread_reg ),
    .X(_07873_));
 sky130_fd_sc_hd__or3b_2 _23473_ (.A(_10662_),
    .B(_07862_),
    .C_N(_07873_),
    .X(_07874_));
 sky130_fd_sc_hd__o211a_2 _23474_ (.A1(io_fetch_data[23]),
    .A2(_07861_),
    .B1(_07874_),
    .C1(_07865_),
    .X(_01446_));
 sky130_fd_sc_hd__buf_1 _23475_ (.A(_03546_),
    .X(_07875_));
 sky130_fd_sc_hd__buf_1 _23476_ (.A(_10670_),
    .X(_07876_));
 sky130_fd_sc_hd__or3b_2 _23477_ (.A(_10994_),
    .B(_07876_),
    .C_N(_07873_),
    .X(_07877_));
 sky130_fd_sc_hd__o211a_2 _23478_ (.A1(io_fetch_data[24]),
    .A2(_07875_),
    .B1(_07877_),
    .C1(_07865_),
    .X(_01447_));
 sky130_fd_sc_hd__or3b_2 _23479_ (.A(\decode.control.io_funct7[0] ),
    .B(_07876_),
    .C_N(_07873_),
    .X(_07878_));
 sky130_fd_sc_hd__buf_1 _23480_ (.A(_04459_),
    .X(_07879_));
 sky130_fd_sc_hd__o211a_2 _23481_ (.A1(io_fetch_data[25]),
    .A2(_07875_),
    .B1(_07878_),
    .C1(_07879_),
    .X(_01448_));
 sky130_fd_sc_hd__or3b_2 _23482_ (.A(\decode.control.io_funct7[1] ),
    .B(_07876_),
    .C_N(_07873_),
    .X(_07880_));
 sky130_fd_sc_hd__o211a_2 _23483_ (.A1(io_fetch_data[26]),
    .A2(_07875_),
    .B1(_07880_),
    .C1(_07879_),
    .X(_01449_));
 sky130_fd_sc_hd__or3b_2 _23484_ (.A(\decode.control.io_funct7[2] ),
    .B(_07876_),
    .C_N(_07873_),
    .X(_07881_));
 sky130_fd_sc_hd__o211a_2 _23485_ (.A1(io_fetch_data[27]),
    .A2(_07875_),
    .B1(_07881_),
    .C1(_07879_),
    .X(_01450_));
 sky130_fd_sc_hd__or3b_2 _23486_ (.A(\decode.control.io_funct7[3] ),
    .B(_07876_),
    .C_N(_07873_),
    .X(_07882_));
 sky130_fd_sc_hd__o211a_2 _23487_ (.A1(io_fetch_data[28]),
    .A2(_07875_),
    .B1(_07882_),
    .C1(_07879_),
    .X(_01451_));
 sky130_fd_sc_hd__or3b_2 _23488_ (.A(\decode.control.io_funct7[4] ),
    .B(_07876_),
    .C_N(_07873_),
    .X(_07883_));
 sky130_fd_sc_hd__o211a_2 _23489_ (.A1(io_fetch_data[29]),
    .A2(_07875_),
    .B1(_07883_),
    .C1(_07879_),
    .X(_01452_));
 sky130_fd_sc_hd__or3b_2 _23490_ (.A(\decode.control.io_funct7[5] ),
    .B(_07876_),
    .C_N(_07873_),
    .X(_07884_));
 sky130_fd_sc_hd__o211a_2 _23491_ (.A1(io_fetch_data[30]),
    .A2(_07875_),
    .B1(_07884_),
    .C1(_07879_),
    .X(_01453_));
 sky130_fd_sc_hd__or3b_2 _23492_ (.A(\decode.control.io_funct7[6] ),
    .B(_07876_),
    .C_N(_07873_),
    .X(_07885_));
 sky130_fd_sc_hd__o211a_2 _23493_ (.A1(io_fetch_data[31]),
    .A2(_07875_),
    .B1(_07885_),
    .C1(_07879_),
    .X(_01454_));
 sky130_fd_sc_hd__or3b_2 _23494_ (.A(\decode.io_id_pc[0] ),
    .B(_07876_),
    .C_N(_07873_),
    .X(_07886_));
 sky130_fd_sc_hd__o211a_2 _23495_ (.A1(io_fetch_address[0]),
    .A2(_07875_),
    .B1(_07886_),
    .C1(_07879_),
    .X(_01455_));
 sky130_fd_sc_hd__buf_1 _23496_ (.A(\decode.id_ex_memread_reg ),
    .X(_07887_));
 sky130_fd_sc_hd__or3b_2 _23497_ (.A(\decode.io_id_pc[1] ),
    .B(_07876_),
    .C_N(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__o211a_2 _23498_ (.A1(io_fetch_address[1]),
    .A2(_07875_),
    .B1(_07888_),
    .C1(_07879_),
    .X(_01456_));
 sky130_fd_sc_hd__buf_1 _23499_ (.A(_03546_),
    .X(_07889_));
 sky130_fd_sc_hd__buf_1 _23500_ (.A(_10670_),
    .X(_07890_));
 sky130_fd_sc_hd__or3b_2 _23501_ (.A(\decode.io_id_pc[2] ),
    .B(_07890_),
    .C_N(_07887_),
    .X(_07891_));
 sky130_fd_sc_hd__o211a_2 _23502_ (.A1(io_fetch_address[2]),
    .A2(_07889_),
    .B1(_07891_),
    .C1(_07879_),
    .X(_01457_));
 sky130_fd_sc_hd__or3b_2 _23503_ (.A(\decode.io_id_pc[3] ),
    .B(_07890_),
    .C_N(_07887_),
    .X(_07892_));
 sky130_fd_sc_hd__buf_1 _23504_ (.A(_04459_),
    .X(_07893_));
 sky130_fd_sc_hd__o211a_2 _23505_ (.A1(io_fetch_address[3]),
    .A2(_07889_),
    .B1(_07892_),
    .C1(_07893_),
    .X(_01458_));
 sky130_fd_sc_hd__or3b_2 _23506_ (.A(\decode.io_id_pc[4] ),
    .B(_07890_),
    .C_N(_07887_),
    .X(_07894_));
 sky130_fd_sc_hd__o211a_2 _23507_ (.A1(io_fetch_address[4]),
    .A2(_07889_),
    .B1(_07894_),
    .C1(_07893_),
    .X(_01459_));
 sky130_fd_sc_hd__or3b_2 _23508_ (.A(\decode.io_id_pc[5] ),
    .B(_07890_),
    .C_N(_07887_),
    .X(_07895_));
 sky130_fd_sc_hd__o211a_2 _23509_ (.A1(io_fetch_address[5]),
    .A2(_07889_),
    .B1(_07895_),
    .C1(_07893_),
    .X(_01460_));
 sky130_fd_sc_hd__or3b_2 _23510_ (.A(\decode.io_id_pc[6] ),
    .B(_07890_),
    .C_N(_07887_),
    .X(_07896_));
 sky130_fd_sc_hd__o211a_2 _23511_ (.A1(io_fetch_address[6]),
    .A2(_07889_),
    .B1(_07896_),
    .C1(_07893_),
    .X(_01461_));
 sky130_fd_sc_hd__or3b_2 _23512_ (.A(\decode.io_id_pc[7] ),
    .B(_07890_),
    .C_N(_07887_),
    .X(_07897_));
 sky130_fd_sc_hd__o211a_2 _23513_ (.A1(io_fetch_address[7]),
    .A2(_07889_),
    .B1(_07897_),
    .C1(_07893_),
    .X(_01462_));
 sky130_fd_sc_hd__or3b_2 _23514_ (.A(\decode.io_id_pc[8] ),
    .B(_07890_),
    .C_N(_07887_),
    .X(_07898_));
 sky130_fd_sc_hd__o211a_2 _23515_ (.A1(io_fetch_address[8]),
    .A2(_07889_),
    .B1(_07898_),
    .C1(_07893_),
    .X(_01463_));
 sky130_fd_sc_hd__or3b_2 _23516_ (.A(\decode.io_id_pc[9] ),
    .B(_07890_),
    .C_N(_07887_),
    .X(_07899_));
 sky130_fd_sc_hd__o211a_2 _23517_ (.A1(_06718_),
    .A2(_07889_),
    .B1(_07899_),
    .C1(_07893_),
    .X(_01464_));
 sky130_fd_sc_hd__or3b_2 _23518_ (.A(\decode.io_id_pc[10] ),
    .B(_07890_),
    .C_N(_07887_),
    .X(_07900_));
 sky130_fd_sc_hd__o211a_2 _23519_ (.A1(io_fetch_address[10]),
    .A2(_07889_),
    .B1(_07900_),
    .C1(_07893_),
    .X(_01465_));
 sky130_fd_sc_hd__buf_1 _23520_ (.A(\decode.id_ex_memread_reg ),
    .X(_07901_));
 sky130_fd_sc_hd__or3b_2 _23521_ (.A(\decode.io_id_pc[11] ),
    .B(_07890_),
    .C_N(_07901_),
    .X(_07902_));
 sky130_fd_sc_hd__o211a_2 _23522_ (.A1(io_fetch_address[11]),
    .A2(_07889_),
    .B1(_07902_),
    .C1(_07893_),
    .X(_01466_));
 sky130_fd_sc_hd__buf_1 _23523_ (.A(_03546_),
    .X(_07903_));
 sky130_fd_sc_hd__buf_1 _23524_ (.A(_10670_),
    .X(_07904_));
 sky130_fd_sc_hd__or3b_2 _23525_ (.A(\decode.io_id_pc[12] ),
    .B(_07904_),
    .C_N(_07901_),
    .X(_07905_));
 sky130_fd_sc_hd__o211a_2 _23526_ (.A1(io_fetch_address[12]),
    .A2(_07903_),
    .B1(_07905_),
    .C1(_07893_),
    .X(_01467_));
 sky130_fd_sc_hd__or3b_2 _23527_ (.A(\decode.io_id_pc[13] ),
    .B(_07904_),
    .C_N(_07901_),
    .X(_07906_));
 sky130_fd_sc_hd__buf_1 _23528_ (.A(_04459_),
    .X(_07907_));
 sky130_fd_sc_hd__o211a_2 _23529_ (.A1(io_fetch_address[13]),
    .A2(_07903_),
    .B1(_07906_),
    .C1(_07907_),
    .X(_01468_));
 sky130_fd_sc_hd__or3b_2 _23530_ (.A(\decode.io_id_pc[14] ),
    .B(_07904_),
    .C_N(_07901_),
    .X(_07908_));
 sky130_fd_sc_hd__o211a_2 _23531_ (.A1(io_fetch_address[14]),
    .A2(_07903_),
    .B1(_07908_),
    .C1(_07907_),
    .X(_01469_));
 sky130_fd_sc_hd__or3b_2 _23532_ (.A(\decode.io_id_pc[15] ),
    .B(_07904_),
    .C_N(_07901_),
    .X(_07909_));
 sky130_fd_sc_hd__o211a_2 _23533_ (.A1(io_fetch_address[15]),
    .A2(_07903_),
    .B1(_07909_),
    .C1(_07907_),
    .X(_01470_));
 sky130_fd_sc_hd__or3b_2 _23534_ (.A(\decode.io_id_pc[16] ),
    .B(_07904_),
    .C_N(_07901_),
    .X(_07910_));
 sky130_fd_sc_hd__o211a_2 _23535_ (.A1(io_fetch_address[16]),
    .A2(_07903_),
    .B1(_07910_),
    .C1(_07907_),
    .X(_01471_));
 sky130_fd_sc_hd__or3b_2 _23536_ (.A(\decode.io_id_pc[17] ),
    .B(_07904_),
    .C_N(_07901_),
    .X(_07911_));
 sky130_fd_sc_hd__o211a_2 _23537_ (.A1(_06887_),
    .A2(_07903_),
    .B1(_07911_),
    .C1(_07907_),
    .X(_01472_));
 sky130_fd_sc_hd__or3b_2 _23538_ (.A(\decode.io_id_pc[18] ),
    .B(_07904_),
    .C_N(_07901_),
    .X(_07912_));
 sky130_fd_sc_hd__o211a_2 _23539_ (.A1(io_fetch_address[18]),
    .A2(_07903_),
    .B1(_07912_),
    .C1(_07907_),
    .X(_01473_));
 sky130_fd_sc_hd__or3b_2 _23540_ (.A(\decode.io_id_pc[19] ),
    .B(_07904_),
    .C_N(_07901_),
    .X(_07913_));
 sky130_fd_sc_hd__o211a_2 _23541_ (.A1(io_fetch_address[19]),
    .A2(_07903_),
    .B1(_07913_),
    .C1(_07907_),
    .X(_01474_));
 sky130_fd_sc_hd__or3b_2 _23542_ (.A(\decode.io_id_pc[20] ),
    .B(_07904_),
    .C_N(_07901_),
    .X(_07914_));
 sky130_fd_sc_hd__o211a_2 _23543_ (.A1(io_fetch_address[20]),
    .A2(_07903_),
    .B1(_07914_),
    .C1(_07907_),
    .X(_01475_));
 sky130_fd_sc_hd__buf_1 _23544_ (.A(\decode.id_ex_memread_reg ),
    .X(_07915_));
 sky130_fd_sc_hd__or3b_2 _23545_ (.A(\decode.io_id_pc[21] ),
    .B(_07904_),
    .C_N(_07915_),
    .X(_07916_));
 sky130_fd_sc_hd__o211a_2 _23546_ (.A1(io_fetch_address[21]),
    .A2(_07903_),
    .B1(_07916_),
    .C1(_07907_),
    .X(_01476_));
 sky130_fd_sc_hd__buf_1 _23547_ (.A(_03546_),
    .X(_07917_));
 sky130_fd_sc_hd__buf_1 _23548_ (.A(_10670_),
    .X(_07918_));
 sky130_fd_sc_hd__or3b_2 _23549_ (.A(\decode.io_id_pc[22] ),
    .B(_07918_),
    .C_N(_07915_),
    .X(_07919_));
 sky130_fd_sc_hd__o211a_2 _23550_ (.A1(io_fetch_address[22]),
    .A2(_07917_),
    .B1(_07919_),
    .C1(_07907_),
    .X(_01477_));
 sky130_fd_sc_hd__or3b_2 _23551_ (.A(\decode.io_id_pc[23] ),
    .B(_07918_),
    .C_N(_07915_),
    .X(_07920_));
 sky130_fd_sc_hd__o211a_2 _23552_ (.A1(io_fetch_address[23]),
    .A2(_07917_),
    .B1(_07920_),
    .C1(_05805_),
    .X(_01478_));
 sky130_fd_sc_hd__or3b_2 _23553_ (.A(\decode.io_id_pc[24] ),
    .B(_07918_),
    .C_N(_07915_),
    .X(_07921_));
 sky130_fd_sc_hd__o211a_2 _23554_ (.A1(io_fetch_address[24]),
    .A2(_07917_),
    .B1(_07921_),
    .C1(_05805_),
    .X(_01479_));
 sky130_fd_sc_hd__or3b_2 _23555_ (.A(\decode.io_id_pc[25] ),
    .B(_07918_),
    .C_N(_07915_),
    .X(_07922_));
 sky130_fd_sc_hd__o211a_2 _23556_ (.A1(io_fetch_address[25]),
    .A2(_07917_),
    .B1(_07922_),
    .C1(_05805_),
    .X(_01480_));
 sky130_fd_sc_hd__or3b_2 _23557_ (.A(\decode.io_id_pc[26] ),
    .B(_07918_),
    .C_N(_07915_),
    .X(_07923_));
 sky130_fd_sc_hd__o211a_2 _23558_ (.A1(io_fetch_address[26]),
    .A2(_07917_),
    .B1(_07923_),
    .C1(_05805_),
    .X(_01481_));
 sky130_fd_sc_hd__or3b_2 _23559_ (.A(\decode.io_id_pc[27] ),
    .B(_07918_),
    .C_N(_07915_),
    .X(_07924_));
 sky130_fd_sc_hd__o211a_2 _23560_ (.A1(io_fetch_address[27]),
    .A2(_07917_),
    .B1(_07924_),
    .C1(_05805_),
    .X(_01482_));
 sky130_fd_sc_hd__or3b_2 _23561_ (.A(\decode.io_id_pc[28] ),
    .B(_07918_),
    .C_N(_07915_),
    .X(_07925_));
 sky130_fd_sc_hd__o211a_2 _23562_ (.A1(_06795_),
    .A2(_07917_),
    .B1(_07925_),
    .C1(_05805_),
    .X(_01483_));
 sky130_fd_sc_hd__or3b_2 _23563_ (.A(\decode.io_id_pc[29] ),
    .B(_07918_),
    .C_N(_07915_),
    .X(_07926_));
 sky130_fd_sc_hd__o211a_2 _23564_ (.A1(io_fetch_address[29]),
    .A2(_07917_),
    .B1(_07926_),
    .C1(_05805_),
    .X(_01484_));
 sky130_fd_sc_hd__or3b_2 _23565_ (.A(\decode.io_id_pc[30] ),
    .B(_07918_),
    .C_N(_07915_),
    .X(_07927_));
 sky130_fd_sc_hd__o211a_2 _23566_ (.A1(io_fetch_address[30]),
    .A2(_07917_),
    .B1(_07927_),
    .C1(_05805_),
    .X(_01485_));
 sky130_fd_sc_hd__or3b_2 _23567_ (.A(\decode.io_id_pc[31] ),
    .B(_07918_),
    .C_N(\decode.id_ex_memread_reg ),
    .X(_07928_));
 sky130_fd_sc_hd__o211a_2 _23568_ (.A1(io_fetch_address[31]),
    .A2(_07917_),
    .B1(_07928_),
    .C1(_05805_),
    .X(_01486_));
 sky130_fd_sc_hd__or3b_2 _23569_ (.A(_09900_),
    .B(_06281_),
    .C_N(_09894_),
    .X(_07929_));
 sky130_fd_sc_hd__buf_1 _23570_ (.A(_07929_),
    .X(_07930_));
 sky130_fd_sc_hd__a22o_2 _23571_ (.A1(_09914_),
    .A2(_10761_),
    .B1(_07930_),
    .B2(\fetch.bht.bhtTable_tag[15][0] ),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_2 _23572_ (.A0(_06103_),
    .A1(\fetch.bht.bhtTable_tag[15][1] ),
    .S(_07930_),
    .X(_07931_));
 sky130_fd_sc_hd__buf_1 _23573_ (.A(_07931_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_2 _23574_ (.A0(_06105_),
    .A1(\fetch.bht.bhtTable_tag[15][2] ),
    .S(_07930_),
    .X(_07932_));
 sky130_fd_sc_hd__buf_1 _23575_ (.A(_07932_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_2 _23576_ (.A0(_06107_),
    .A1(\fetch.bht.bhtTable_tag[15][3] ),
    .S(_07930_),
    .X(_07933_));
 sky130_fd_sc_hd__buf_1 _23577_ (.A(_07933_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_2 _23578_ (.A0(_06109_),
    .A1(\fetch.bht.bhtTable_tag[15][4] ),
    .S(_07930_),
    .X(_07934_));
 sky130_fd_sc_hd__buf_1 _23579_ (.A(_07934_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_2 _23580_ (.A0(_06111_),
    .A1(\fetch.bht.bhtTable_tag[15][5] ),
    .S(_07930_),
    .X(_07935_));
 sky130_fd_sc_hd__buf_1 _23581_ (.A(_07935_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_2 _23582_ (.A0(_06113_),
    .A1(\fetch.bht.bhtTable_tag[15][6] ),
    .S(_07930_),
    .X(_07936_));
 sky130_fd_sc_hd__buf_1 _23583_ (.A(_07936_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_2 _23584_ (.A0(_06115_),
    .A1(\fetch.bht.bhtTable_tag[15][7] ),
    .S(_07930_),
    .X(_07937_));
 sky130_fd_sc_hd__buf_1 _23585_ (.A(_07937_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_2 _23586_ (.A0(_06117_),
    .A1(\fetch.bht.bhtTable_tag[15][8] ),
    .S(_07930_),
    .X(_07938_));
 sky130_fd_sc_hd__buf_1 _23587_ (.A(_07938_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_2 _23588_ (.A0(_06119_),
    .A1(\fetch.bht.bhtTable_tag[15][9] ),
    .S(_07930_),
    .X(_07939_));
 sky130_fd_sc_hd__buf_1 _23589_ (.A(_07939_),
    .X(_01496_));
 sky130_fd_sc_hd__buf_1 _23590_ (.A(_07929_),
    .X(_07940_));
 sky130_fd_sc_hd__buf_1 _23591_ (.A(_07940_),
    .X(_07941_));
 sky130_fd_sc_hd__mux2_2 _23592_ (.A0(_06122_),
    .A1(\fetch.bht.bhtTable_tag[15][10] ),
    .S(_07941_),
    .X(_07942_));
 sky130_fd_sc_hd__buf_1 _23593_ (.A(_07942_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_2 _23594_ (.A0(_06124_),
    .A1(\fetch.bht.bhtTable_tag[15][11] ),
    .S(_07941_),
    .X(_07943_));
 sky130_fd_sc_hd__buf_1 _23595_ (.A(_07943_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_2 _23596_ (.A0(_06126_),
    .A1(\fetch.bht.bhtTable_tag[15][12] ),
    .S(_07941_),
    .X(_07944_));
 sky130_fd_sc_hd__buf_1 _23597_ (.A(_07944_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_2 _23598_ (.A0(_06128_),
    .A1(\fetch.bht.bhtTable_tag[15][13] ),
    .S(_07941_),
    .X(_07945_));
 sky130_fd_sc_hd__buf_1 _23599_ (.A(_07945_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_2 _23600_ (.A0(_06130_),
    .A1(\fetch.bht.bhtTable_tag[15][14] ),
    .S(_07941_),
    .X(_07946_));
 sky130_fd_sc_hd__buf_1 _23601_ (.A(_07946_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_2 _23602_ (.A0(_06132_),
    .A1(\fetch.bht.bhtTable_tag[15][15] ),
    .S(_07941_),
    .X(_07947_));
 sky130_fd_sc_hd__buf_1 _23603_ (.A(_07947_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_2 _23604_ (.A0(_06134_),
    .A1(\fetch.bht.bhtTable_tag[15][16] ),
    .S(_07941_),
    .X(_07948_));
 sky130_fd_sc_hd__buf_1 _23605_ (.A(_07948_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_2 _23606_ (.A0(_06136_),
    .A1(\fetch.bht.bhtTable_tag[15][17] ),
    .S(_07941_),
    .X(_07949_));
 sky130_fd_sc_hd__buf_1 _23607_ (.A(_07949_),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_2 _23608_ (.A0(_06138_),
    .A1(\fetch.bht.bhtTable_tag[15][18] ),
    .S(_07941_),
    .X(_07950_));
 sky130_fd_sc_hd__buf_1 _23609_ (.A(_07950_),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_2 _23610_ (.A0(_06140_),
    .A1(\fetch.bht.bhtTable_tag[15][19] ),
    .S(_07941_),
    .X(_07951_));
 sky130_fd_sc_hd__buf_1 _23611_ (.A(_07951_),
    .X(_01506_));
 sky130_fd_sc_hd__buf_1 _23612_ (.A(_07940_),
    .X(_07952_));
 sky130_fd_sc_hd__mux2_2 _23613_ (.A0(_06143_),
    .A1(\fetch.bht.bhtTable_tag[15][20] ),
    .S(_07952_),
    .X(_07953_));
 sky130_fd_sc_hd__buf_1 _23614_ (.A(_07953_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_2 _23615_ (.A0(_06145_),
    .A1(\fetch.bht.bhtTable_tag[15][21] ),
    .S(_07952_),
    .X(_07954_));
 sky130_fd_sc_hd__buf_1 _23616_ (.A(_07954_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_2 _23617_ (.A0(_06147_),
    .A1(\fetch.bht.bhtTable_tag[15][22] ),
    .S(_07952_),
    .X(_07955_));
 sky130_fd_sc_hd__buf_1 _23618_ (.A(_07955_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_2 _23619_ (.A0(_06149_),
    .A1(\fetch.bht.bhtTable_tag[15][23] ),
    .S(_07952_),
    .X(_07956_));
 sky130_fd_sc_hd__buf_1 _23620_ (.A(_07956_),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_2 _23621_ (.A0(_06151_),
    .A1(\fetch.bht.bhtTable_tag[15][24] ),
    .S(_07952_),
    .X(_07957_));
 sky130_fd_sc_hd__buf_1 _23622_ (.A(_07957_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_2 _23623_ (.A0(_06153_),
    .A1(\fetch.bht.bhtTable_tag[15][25] ),
    .S(_07952_),
    .X(_07958_));
 sky130_fd_sc_hd__buf_1 _23624_ (.A(_07958_),
    .X(_01512_));
 sky130_fd_sc_hd__and3_2 _23625_ (.A(_09885_),
    .B(_09887_),
    .C(_09917_),
    .X(_07959_));
 sky130_fd_sc_hd__buf_1 _23626_ (.A(_07959_),
    .X(_07960_));
 sky130_fd_sc_hd__buf_1 _23627_ (.A(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__mux2_2 _23628_ (.A0(\fetch.bht.bhtTable_tag[2][0] ),
    .A1(_10820_),
    .S(_07961_),
    .X(_07962_));
 sky130_fd_sc_hd__buf_1 _23629_ (.A(_07962_),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_2 _23630_ (.A0(\fetch.bht.bhtTable_tag[2][1] ),
    .A1(_10821_),
    .S(_07961_),
    .X(_07963_));
 sky130_fd_sc_hd__buf_1 _23631_ (.A(_07963_),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_2 _23632_ (.A0(\fetch.bht.bhtTable_tag[2][2] ),
    .A1(_10881_),
    .S(_07961_),
    .X(_07964_));
 sky130_fd_sc_hd__buf_1 _23633_ (.A(_07964_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_2 _23634_ (.A0(\fetch.bht.bhtTable_tag[2][3] ),
    .A1(_10817_),
    .S(_07961_),
    .X(_07965_));
 sky130_fd_sc_hd__buf_1 _23635_ (.A(_07965_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_2 _23636_ (.A0(\fetch.bht.bhtTable_tag[2][4] ),
    .A1(_10878_),
    .S(_07961_),
    .X(_07966_));
 sky130_fd_sc_hd__buf_1 _23637_ (.A(_07966_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_2 _23638_ (.A0(\fetch.bht.bhtTable_tag[2][5] ),
    .A1(_10812_),
    .S(_07961_),
    .X(_07967_));
 sky130_fd_sc_hd__buf_1 _23639_ (.A(_07967_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_2 _23640_ (.A0(\fetch.bht.bhtTable_tag[2][6] ),
    .A1(\csr.io_mem_pc[12] ),
    .S(_07961_),
    .X(_07968_));
 sky130_fd_sc_hd__buf_1 _23641_ (.A(_07968_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_2 _23642_ (.A0(\fetch.bht.bhtTable_tag[2][7] ),
    .A1(_10871_),
    .S(_07961_),
    .X(_07969_));
 sky130_fd_sc_hd__buf_1 _23643_ (.A(_07969_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_2 _23644_ (.A0(\fetch.bht.bhtTable_tag[2][8] ),
    .A1(_10872_),
    .S(_07961_),
    .X(_07970_));
 sky130_fd_sc_hd__buf_1 _23645_ (.A(_07970_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_2 _23646_ (.A0(\fetch.bht.bhtTable_tag[2][9] ),
    .A1(_10807_),
    .S(_07961_),
    .X(_07971_));
 sky130_fd_sc_hd__buf_1 _23647_ (.A(_07971_),
    .X(_01522_));
 sky130_fd_sc_hd__buf_1 _23648_ (.A(_07960_),
    .X(_07972_));
 sky130_fd_sc_hd__mux2_2 _23649_ (.A0(\fetch.bht.bhtTable_tag[2][10] ),
    .A1(_10868_),
    .S(_07972_),
    .X(_07973_));
 sky130_fd_sc_hd__buf_1 _23650_ (.A(_07973_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_2 _23651_ (.A0(\fetch.bht.bhtTable_tag[2][11] ),
    .A1(_10803_),
    .S(_07972_),
    .X(_07974_));
 sky130_fd_sc_hd__buf_1 _23652_ (.A(_07974_),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_2 _23653_ (.A0(\fetch.bht.bhtTable_tag[2][12] ),
    .A1(\csr.io_mem_pc[18] ),
    .S(_07972_),
    .X(_07975_));
 sky130_fd_sc_hd__buf_1 _23654_ (.A(_07975_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_2 _23655_ (.A0(\fetch.bht.bhtTable_tag[2][13] ),
    .A1(_10800_),
    .S(_07972_),
    .X(_07976_));
 sky130_fd_sc_hd__buf_1 _23656_ (.A(_07976_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_2 _23657_ (.A0(\fetch.bht.bhtTable_tag[2][14] ),
    .A1(_10795_),
    .S(_07972_),
    .X(_07977_));
 sky130_fd_sc_hd__buf_1 _23658_ (.A(_07977_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_2 _23659_ (.A0(\fetch.bht.bhtTable_tag[2][15] ),
    .A1(\csr.io_mem_pc[21] ),
    .S(_07972_),
    .X(_07978_));
 sky130_fd_sc_hd__buf_1 _23660_ (.A(_07978_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_2 _23661_ (.A0(\fetch.bht.bhtTable_tag[2][16] ),
    .A1(_10787_),
    .S(_07972_),
    .X(_07979_));
 sky130_fd_sc_hd__buf_1 _23662_ (.A(_07979_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_2 _23663_ (.A0(\fetch.bht.bhtTable_tag[2][17] ),
    .A1(\csr.io_mem_pc[23] ),
    .S(_07972_),
    .X(_07980_));
 sky130_fd_sc_hd__buf_1 _23664_ (.A(_07980_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_2 _23665_ (.A0(\fetch.bht.bhtTable_tag[2][18] ),
    .A1(_10772_),
    .S(_07972_),
    .X(_07981_));
 sky130_fd_sc_hd__buf_1 _23666_ (.A(_07981_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_2 _23667_ (.A0(\fetch.bht.bhtTable_tag[2][19] ),
    .A1(_10773_),
    .S(_07972_),
    .X(_07982_));
 sky130_fd_sc_hd__buf_1 _23668_ (.A(_07982_),
    .X(_01532_));
 sky130_fd_sc_hd__buf_1 _23669_ (.A(_07959_),
    .X(_07983_));
 sky130_fd_sc_hd__mux2_2 _23670_ (.A0(\fetch.bht.bhtTable_tag[2][20] ),
    .A1(_10760_),
    .S(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__buf_1 _23671_ (.A(_07984_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_2 _23672_ (.A0(\fetch.bht.bhtTable_tag[2][21] ),
    .A1(_10759_),
    .S(_07983_),
    .X(_07985_));
 sky130_fd_sc_hd__buf_1 _23673_ (.A(_07985_),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_2 _23674_ (.A0(\fetch.bht.bhtTable_tag[2][22] ),
    .A1(_10771_),
    .S(_07983_),
    .X(_07986_));
 sky130_fd_sc_hd__buf_1 _23675_ (.A(_07986_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_2 _23676_ (.A0(\fetch.bht.bhtTable_tag[2][23] ),
    .A1(\csr.io_mem_pc[29] ),
    .S(_07983_),
    .X(_07987_));
 sky130_fd_sc_hd__buf_1 _23677_ (.A(_07987_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_2 _23678_ (.A0(\fetch.bht.bhtTable_tag[2][24] ),
    .A1(_10777_),
    .S(_07983_),
    .X(_07988_));
 sky130_fd_sc_hd__buf_1 _23679_ (.A(_07988_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_2 _23680_ (.A0(\fetch.bht.bhtTable_tag[2][25] ),
    .A1(\csr.io_mem_pc[31] ),
    .S(_07983_),
    .X(_07989_));
 sky130_fd_sc_hd__buf_1 _23681_ (.A(_07989_),
    .X(_01538_));
 sky130_fd_sc_hd__and3_2 _23682_ (.A(_09885_),
    .B(_09894_),
    .C(_09917_),
    .X(_07990_));
 sky130_fd_sc_hd__buf_1 _23683_ (.A(_07990_),
    .X(_07991_));
 sky130_fd_sc_hd__buf_1 _23684_ (.A(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__mux2_2 _23685_ (.A0(\fetch.bht.bhtTable_tag[3][0] ),
    .A1(_10820_),
    .S(_07992_),
    .X(_07993_));
 sky130_fd_sc_hd__buf_1 _23686_ (.A(_07993_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_2 _23687_ (.A0(\fetch.bht.bhtTable_tag[3][1] ),
    .A1(_10821_),
    .S(_07992_),
    .X(_07994_));
 sky130_fd_sc_hd__buf_1 _23688_ (.A(_07994_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_2 _23689_ (.A0(\fetch.bht.bhtTable_tag[3][2] ),
    .A1(_10881_),
    .S(_07992_),
    .X(_07995_));
 sky130_fd_sc_hd__buf_1 _23690_ (.A(_07995_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_2 _23691_ (.A0(\fetch.bht.bhtTable_tag[3][3] ),
    .A1(_10817_),
    .S(_07992_),
    .X(_07996_));
 sky130_fd_sc_hd__buf_1 _23692_ (.A(_07996_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_2 _23693_ (.A0(\fetch.bht.bhtTable_tag[3][4] ),
    .A1(_10878_),
    .S(_07992_),
    .X(_07997_));
 sky130_fd_sc_hd__buf_1 _23694_ (.A(_07997_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_2 _23695_ (.A0(\fetch.bht.bhtTable_tag[3][5] ),
    .A1(_10812_),
    .S(_07992_),
    .X(_07998_));
 sky130_fd_sc_hd__buf_1 _23696_ (.A(_07998_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_2 _23697_ (.A0(\fetch.bht.bhtTable_tag[3][6] ),
    .A1(\csr.io_mem_pc[12] ),
    .S(_07992_),
    .X(_07999_));
 sky130_fd_sc_hd__buf_1 _23698_ (.A(_07999_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_2 _23699_ (.A0(\fetch.bht.bhtTable_tag[3][7] ),
    .A1(_10871_),
    .S(_07992_),
    .X(_08000_));
 sky130_fd_sc_hd__buf_1 _23700_ (.A(_08000_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_2 _23701_ (.A0(\fetch.bht.bhtTable_tag[3][8] ),
    .A1(_10872_),
    .S(_07992_),
    .X(_08001_));
 sky130_fd_sc_hd__buf_1 _23702_ (.A(_08001_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_2 _23703_ (.A0(\fetch.bht.bhtTable_tag[3][9] ),
    .A1(_10807_),
    .S(_07992_),
    .X(_08002_));
 sky130_fd_sc_hd__buf_1 _23704_ (.A(_08002_),
    .X(_01548_));
 sky130_fd_sc_hd__buf_1 _23705_ (.A(_07991_),
    .X(_08003_));
 sky130_fd_sc_hd__mux2_2 _23706_ (.A0(\fetch.bht.bhtTable_tag[3][10] ),
    .A1(_10868_),
    .S(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__buf_1 _23707_ (.A(_08004_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_2 _23708_ (.A0(\fetch.bht.bhtTable_tag[3][11] ),
    .A1(_10803_),
    .S(_08003_),
    .X(_08005_));
 sky130_fd_sc_hd__buf_1 _23709_ (.A(_08005_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_2 _23710_ (.A0(\fetch.bht.bhtTable_tag[3][12] ),
    .A1(\csr.io_mem_pc[18] ),
    .S(_08003_),
    .X(_08006_));
 sky130_fd_sc_hd__buf_1 _23711_ (.A(_08006_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_2 _23712_ (.A0(\fetch.bht.bhtTable_tag[3][13] ),
    .A1(_10800_),
    .S(_08003_),
    .X(_08007_));
 sky130_fd_sc_hd__buf_1 _23713_ (.A(_08007_),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_2 _23714_ (.A0(\fetch.bht.bhtTable_tag[3][14] ),
    .A1(_10795_),
    .S(_08003_),
    .X(_08008_));
 sky130_fd_sc_hd__buf_1 _23715_ (.A(_08008_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_2 _23716_ (.A0(\fetch.bht.bhtTable_tag[3][15] ),
    .A1(\csr.io_mem_pc[21] ),
    .S(_08003_),
    .X(_08009_));
 sky130_fd_sc_hd__buf_1 _23717_ (.A(_08009_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_2 _23718_ (.A0(\fetch.bht.bhtTable_tag[3][16] ),
    .A1(_10787_),
    .S(_08003_),
    .X(_08010_));
 sky130_fd_sc_hd__buf_1 _23719_ (.A(_08010_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_2 _23720_ (.A0(\fetch.bht.bhtTable_tag[3][17] ),
    .A1(\csr.io_mem_pc[23] ),
    .S(_08003_),
    .X(_08011_));
 sky130_fd_sc_hd__buf_1 _23721_ (.A(_08011_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_2 _23722_ (.A0(\fetch.bht.bhtTable_tag[3][18] ),
    .A1(_10772_),
    .S(_08003_),
    .X(_08012_));
 sky130_fd_sc_hd__buf_1 _23723_ (.A(_08012_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_2 _23724_ (.A0(\fetch.bht.bhtTable_tag[3][19] ),
    .A1(_10773_),
    .S(_08003_),
    .X(_08013_));
 sky130_fd_sc_hd__buf_1 _23725_ (.A(_08013_),
    .X(_01558_));
 sky130_fd_sc_hd__buf_1 _23726_ (.A(_07990_),
    .X(_08014_));
 sky130_fd_sc_hd__mux2_2 _23727_ (.A0(\fetch.bht.bhtTable_tag[3][20] ),
    .A1(_10760_),
    .S(_08014_),
    .X(_08015_));
 sky130_fd_sc_hd__buf_1 _23728_ (.A(_08015_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_2 _23729_ (.A0(\fetch.bht.bhtTable_tag[3][21] ),
    .A1(_10759_),
    .S(_08014_),
    .X(_08016_));
 sky130_fd_sc_hd__buf_1 _23730_ (.A(_08016_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_2 _23731_ (.A0(\fetch.bht.bhtTable_tag[3][22] ),
    .A1(_10771_),
    .S(_08014_),
    .X(_08017_));
 sky130_fd_sc_hd__buf_1 _23732_ (.A(_08017_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_2 _23733_ (.A0(\fetch.bht.bhtTable_tag[3][23] ),
    .A1(\csr.io_mem_pc[29] ),
    .S(_08014_),
    .X(_08018_));
 sky130_fd_sc_hd__buf_1 _23734_ (.A(_08018_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_2 _23735_ (.A0(\fetch.bht.bhtTable_tag[3][24] ),
    .A1(_10777_),
    .S(_08014_),
    .X(_08019_));
 sky130_fd_sc_hd__buf_1 _23736_ (.A(_08019_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_2 _23737_ (.A0(\fetch.bht.bhtTable_tag[3][25] ),
    .A1(\csr.io_mem_pc[31] ),
    .S(_08014_),
    .X(_08020_));
 sky130_fd_sc_hd__buf_1 _23738_ (.A(_08020_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_2 _23739_ (.A0(_06101_),
    .A1(\fetch.bht.bhtTable_tag[9][0] ),
    .S(_09907_),
    .X(_08021_));
 sky130_fd_sc_hd__buf_1 _23740_ (.A(_08021_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_2 _23741_ (.A0(_06103_),
    .A1(\fetch.bht.bhtTable_tag[9][1] ),
    .S(_09907_),
    .X(_08022_));
 sky130_fd_sc_hd__buf_1 _23742_ (.A(_08022_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_2 _23743_ (.A0(_06105_),
    .A1(\fetch.bht.bhtTable_tag[9][2] ),
    .S(_09907_),
    .X(_08023_));
 sky130_fd_sc_hd__buf_1 _23744_ (.A(_08023_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_2 _23745_ (.A0(_06107_),
    .A1(\fetch.bht.bhtTable_tag[9][3] ),
    .S(_09907_),
    .X(_08024_));
 sky130_fd_sc_hd__buf_1 _23746_ (.A(_08024_),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_2 _23747_ (.A0(_06109_),
    .A1(\fetch.bht.bhtTable_tag[9][4] ),
    .S(_09907_),
    .X(_08025_));
 sky130_fd_sc_hd__buf_1 _23748_ (.A(_08025_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_2 _23749_ (.A0(_06111_),
    .A1(\fetch.bht.bhtTable_tag[9][5] ),
    .S(_09907_),
    .X(_08026_));
 sky130_fd_sc_hd__buf_1 _23750_ (.A(_08026_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_2 _23751_ (.A0(_06113_),
    .A1(\fetch.bht.bhtTable_tag[9][6] ),
    .S(_09907_),
    .X(_08027_));
 sky130_fd_sc_hd__buf_1 _23752_ (.A(_08027_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_2 _23753_ (.A0(_06115_),
    .A1(\fetch.bht.bhtTable_tag[9][7] ),
    .S(_09907_),
    .X(_08028_));
 sky130_fd_sc_hd__buf_1 _23754_ (.A(_08028_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_2 _23755_ (.A0(_06117_),
    .A1(\fetch.bht.bhtTable_tag[9][8] ),
    .S(_09907_),
    .X(_08029_));
 sky130_fd_sc_hd__buf_1 _23756_ (.A(_08029_),
    .X(_01573_));
 sky130_fd_sc_hd__buf_1 _23757_ (.A(_09905_),
    .X(_08030_));
 sky130_fd_sc_hd__mux2_2 _23758_ (.A0(_06119_),
    .A1(\fetch.bht.bhtTable_tag[9][9] ),
    .S(_08030_),
    .X(_08031_));
 sky130_fd_sc_hd__buf_1 _23759_ (.A(_08031_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_2 _23760_ (.A0(_06122_),
    .A1(\fetch.bht.bhtTable_tag[9][10] ),
    .S(_08030_),
    .X(_08032_));
 sky130_fd_sc_hd__buf_1 _23761_ (.A(_08032_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_2 _23762_ (.A0(_06124_),
    .A1(\fetch.bht.bhtTable_tag[9][11] ),
    .S(_08030_),
    .X(_08033_));
 sky130_fd_sc_hd__buf_1 _23763_ (.A(_08033_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_2 _23764_ (.A0(_06126_),
    .A1(\fetch.bht.bhtTable_tag[9][12] ),
    .S(_08030_),
    .X(_08034_));
 sky130_fd_sc_hd__buf_1 _23765_ (.A(_08034_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_2 _23766_ (.A0(_06128_),
    .A1(\fetch.bht.bhtTable_tag[9][13] ),
    .S(_08030_),
    .X(_08035_));
 sky130_fd_sc_hd__buf_1 _23767_ (.A(_08035_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_2 _23768_ (.A0(_06130_),
    .A1(\fetch.bht.bhtTable_tag[9][14] ),
    .S(_08030_),
    .X(_08036_));
 sky130_fd_sc_hd__buf_1 _23769_ (.A(_08036_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_2 _23770_ (.A0(_06132_),
    .A1(\fetch.bht.bhtTable_tag[9][15] ),
    .S(_08030_),
    .X(_08037_));
 sky130_fd_sc_hd__buf_1 _23771_ (.A(_08037_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_2 _23772_ (.A0(_06134_),
    .A1(\fetch.bht.bhtTable_tag[9][16] ),
    .S(_08030_),
    .X(_08038_));
 sky130_fd_sc_hd__buf_1 _23773_ (.A(_08038_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_2 _23774_ (.A0(_06136_),
    .A1(\fetch.bht.bhtTable_tag[9][17] ),
    .S(_08030_),
    .X(_08039_));
 sky130_fd_sc_hd__buf_1 _23775_ (.A(_08039_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_2 _23776_ (.A0(_06138_),
    .A1(\fetch.bht.bhtTable_tag[9][18] ),
    .S(_08030_),
    .X(_08040_));
 sky130_fd_sc_hd__buf_1 _23777_ (.A(_08040_),
    .X(_01583_));
 sky130_fd_sc_hd__buf_1 _23778_ (.A(_09905_),
    .X(_08041_));
 sky130_fd_sc_hd__mux2_2 _23779_ (.A0(_06140_),
    .A1(\fetch.bht.bhtTable_tag[9][19] ),
    .S(_08041_),
    .X(_08042_));
 sky130_fd_sc_hd__buf_1 _23780_ (.A(_08042_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_2 _23781_ (.A0(_06143_),
    .A1(\fetch.bht.bhtTable_tag[9][20] ),
    .S(_08041_),
    .X(_08043_));
 sky130_fd_sc_hd__buf_1 _23782_ (.A(_08043_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_2 _23783_ (.A0(_06145_),
    .A1(\fetch.bht.bhtTable_tag[9][21] ),
    .S(_08041_),
    .X(_08044_));
 sky130_fd_sc_hd__buf_1 _23784_ (.A(_08044_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_2 _23785_ (.A0(_06147_),
    .A1(\fetch.bht.bhtTable_tag[9][22] ),
    .S(_08041_),
    .X(_08045_));
 sky130_fd_sc_hd__buf_1 _23786_ (.A(_08045_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_2 _23787_ (.A0(_06149_),
    .A1(\fetch.bht.bhtTable_tag[9][23] ),
    .S(_08041_),
    .X(_08046_));
 sky130_fd_sc_hd__buf_1 _23788_ (.A(_08046_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_2 _23789_ (.A0(_06151_),
    .A1(\fetch.bht.bhtTable_tag[9][24] ),
    .S(_08041_),
    .X(_08047_));
 sky130_fd_sc_hd__buf_1 _23790_ (.A(_08047_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_2 _23791_ (.A0(_06153_),
    .A1(\fetch.bht.bhtTable_tag[9][25] ),
    .S(_08041_),
    .X(_08048_));
 sky130_fd_sc_hd__buf_1 _23792_ (.A(_08048_),
    .X(_01590_));
 sky130_fd_sc_hd__buf_1 _23793_ (.A(\execute.io_target_pc[0] ),
    .X(_08049_));
 sky130_fd_sc_hd__mux2_2 _23794_ (.A0(_08049_),
    .A1(\fetch.bht.bhtTable_target_pc[15][0] ),
    .S(_07952_),
    .X(_08050_));
 sky130_fd_sc_hd__buf_1 _23795_ (.A(_08050_),
    .X(_01591_));
 sky130_fd_sc_hd__buf_1 _23796_ (.A(\execute.io_target_pc[1] ),
    .X(_08051_));
 sky130_fd_sc_hd__mux2_2 _23797_ (.A0(_08051_),
    .A1(\fetch.bht.bhtTable_target_pc[15][1] ),
    .S(_07952_),
    .X(_08052_));
 sky130_fd_sc_hd__buf_1 _23798_ (.A(_08052_),
    .X(_01592_));
 sky130_fd_sc_hd__buf_1 _23799_ (.A(\execute.io_target_pc[2] ),
    .X(_08053_));
 sky130_fd_sc_hd__mux2_2 _23800_ (.A0(_08053_),
    .A1(\fetch.bht.bhtTable_target_pc[15][2] ),
    .S(_07952_),
    .X(_08054_));
 sky130_fd_sc_hd__buf_1 _23801_ (.A(_08054_),
    .X(_01593_));
 sky130_fd_sc_hd__buf_1 _23802_ (.A(\execute.io_target_pc[3] ),
    .X(_08055_));
 sky130_fd_sc_hd__mux2_2 _23803_ (.A0(_08055_),
    .A1(\fetch.bht.bhtTable_target_pc[15][3] ),
    .S(_07952_),
    .X(_08056_));
 sky130_fd_sc_hd__buf_1 _23804_ (.A(_08056_),
    .X(_01594_));
 sky130_fd_sc_hd__buf_1 _23805_ (.A(\execute.io_target_pc[4] ),
    .X(_08057_));
 sky130_fd_sc_hd__buf_1 _23806_ (.A(_07929_),
    .X(_08058_));
 sky130_fd_sc_hd__mux2_2 _23807_ (.A0(_08057_),
    .A1(\fetch.bht.bhtTable_target_pc[15][4] ),
    .S(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__buf_1 _23808_ (.A(_08059_),
    .X(_01595_));
 sky130_fd_sc_hd__buf_1 _23809_ (.A(\execute.io_target_pc[5] ),
    .X(_08060_));
 sky130_fd_sc_hd__mux2_2 _23810_ (.A0(_08060_),
    .A1(\fetch.bht.bhtTable_target_pc[15][5] ),
    .S(_08058_),
    .X(_08061_));
 sky130_fd_sc_hd__buf_1 _23811_ (.A(_08061_),
    .X(_01596_));
 sky130_fd_sc_hd__buf_1 _23812_ (.A(\execute.io_target_pc[6] ),
    .X(_08062_));
 sky130_fd_sc_hd__mux2_2 _23813_ (.A0(_08062_),
    .A1(\fetch.bht.bhtTable_target_pc[15][6] ),
    .S(_08058_),
    .X(_08063_));
 sky130_fd_sc_hd__buf_1 _23814_ (.A(_08063_),
    .X(_01597_));
 sky130_fd_sc_hd__buf_1 _23815_ (.A(\execute.io_target_pc[7] ),
    .X(_08064_));
 sky130_fd_sc_hd__mux2_2 _23816_ (.A0(_08064_),
    .A1(\fetch.bht.bhtTable_target_pc[15][7] ),
    .S(_08058_),
    .X(_08065_));
 sky130_fd_sc_hd__buf_1 _23817_ (.A(_08065_),
    .X(_01598_));
 sky130_fd_sc_hd__buf_1 _23818_ (.A(\execute.io_target_pc[8] ),
    .X(_08066_));
 sky130_fd_sc_hd__mux2_2 _23819_ (.A0(_08066_),
    .A1(\fetch.bht.bhtTable_target_pc[15][8] ),
    .S(_08058_),
    .X(_08067_));
 sky130_fd_sc_hd__buf_1 _23820_ (.A(_08067_),
    .X(_01599_));
 sky130_fd_sc_hd__buf_1 _23821_ (.A(\execute.io_target_pc[9] ),
    .X(_08068_));
 sky130_fd_sc_hd__mux2_2 _23822_ (.A0(_08068_),
    .A1(\fetch.bht.bhtTable_target_pc[15][9] ),
    .S(_08058_),
    .X(_08069_));
 sky130_fd_sc_hd__buf_1 _23823_ (.A(_08069_),
    .X(_01600_));
 sky130_fd_sc_hd__buf_1 _23824_ (.A(\execute.io_target_pc[10] ),
    .X(_08070_));
 sky130_fd_sc_hd__mux2_2 _23825_ (.A0(_08070_),
    .A1(\fetch.bht.bhtTable_target_pc[15][10] ),
    .S(_08058_),
    .X(_08071_));
 sky130_fd_sc_hd__buf_1 _23826_ (.A(_08071_),
    .X(_01601_));
 sky130_fd_sc_hd__buf_1 _23827_ (.A(\execute.io_target_pc[11] ),
    .X(_08072_));
 sky130_fd_sc_hd__mux2_2 _23828_ (.A0(_08072_),
    .A1(\fetch.bht.bhtTable_target_pc[15][11] ),
    .S(_08058_),
    .X(_08073_));
 sky130_fd_sc_hd__buf_1 _23829_ (.A(_08073_),
    .X(_01602_));
 sky130_fd_sc_hd__buf_1 _23830_ (.A(\execute.io_target_pc[12] ),
    .X(_08074_));
 sky130_fd_sc_hd__mux2_2 _23831_ (.A0(_08074_),
    .A1(\fetch.bht.bhtTable_target_pc[15][12] ),
    .S(_08058_),
    .X(_08075_));
 sky130_fd_sc_hd__buf_1 _23832_ (.A(_08075_),
    .X(_01603_));
 sky130_fd_sc_hd__buf_1 _23833_ (.A(\execute.io_target_pc[13] ),
    .X(_08076_));
 sky130_fd_sc_hd__mux2_2 _23834_ (.A0(_08076_),
    .A1(\fetch.bht.bhtTable_target_pc[15][13] ),
    .S(_08058_),
    .X(_08077_));
 sky130_fd_sc_hd__buf_1 _23835_ (.A(_08077_),
    .X(_01604_));
 sky130_fd_sc_hd__buf_1 _23836_ (.A(\execute.io_target_pc[14] ),
    .X(_08078_));
 sky130_fd_sc_hd__buf_1 _23837_ (.A(_07929_),
    .X(_08079_));
 sky130_fd_sc_hd__mux2_2 _23838_ (.A0(_08078_),
    .A1(\fetch.bht.bhtTable_target_pc[15][14] ),
    .S(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__buf_1 _23839_ (.A(_08080_),
    .X(_01605_));
 sky130_fd_sc_hd__buf_1 _23840_ (.A(\execute.io_target_pc[15] ),
    .X(_08081_));
 sky130_fd_sc_hd__mux2_2 _23841_ (.A0(_08081_),
    .A1(\fetch.bht.bhtTable_target_pc[15][15] ),
    .S(_08079_),
    .X(_08082_));
 sky130_fd_sc_hd__buf_1 _23842_ (.A(_08082_),
    .X(_01606_));
 sky130_fd_sc_hd__buf_1 _23843_ (.A(\execute.io_target_pc[16] ),
    .X(_08083_));
 sky130_fd_sc_hd__mux2_2 _23844_ (.A0(_08083_),
    .A1(\fetch.bht.bhtTable_target_pc[15][16] ),
    .S(_08079_),
    .X(_08084_));
 sky130_fd_sc_hd__buf_1 _23845_ (.A(_08084_),
    .X(_01607_));
 sky130_fd_sc_hd__buf_1 _23846_ (.A(\execute.io_target_pc[17] ),
    .X(_08085_));
 sky130_fd_sc_hd__mux2_2 _23847_ (.A0(_08085_),
    .A1(\fetch.bht.bhtTable_target_pc[15][17] ),
    .S(_08079_),
    .X(_08086_));
 sky130_fd_sc_hd__buf_1 _23848_ (.A(_08086_),
    .X(_01608_));
 sky130_fd_sc_hd__buf_1 _23849_ (.A(\execute.io_target_pc[18] ),
    .X(_08087_));
 sky130_fd_sc_hd__mux2_2 _23850_ (.A0(_08087_),
    .A1(\fetch.bht.bhtTable_target_pc[15][18] ),
    .S(_08079_),
    .X(_08088_));
 sky130_fd_sc_hd__buf_1 _23851_ (.A(_08088_),
    .X(_01609_));
 sky130_fd_sc_hd__buf_1 _23852_ (.A(\execute.io_target_pc[19] ),
    .X(_08089_));
 sky130_fd_sc_hd__mux2_2 _23853_ (.A0(_08089_),
    .A1(\fetch.bht.bhtTable_target_pc[15][19] ),
    .S(_08079_),
    .X(_08090_));
 sky130_fd_sc_hd__buf_1 _23854_ (.A(_08090_),
    .X(_01610_));
 sky130_fd_sc_hd__buf_1 _23855_ (.A(\execute.io_target_pc[20] ),
    .X(_08091_));
 sky130_fd_sc_hd__mux2_2 _23856_ (.A0(_08091_),
    .A1(\fetch.bht.bhtTable_target_pc[15][20] ),
    .S(_08079_),
    .X(_08092_));
 sky130_fd_sc_hd__buf_1 _23857_ (.A(_08092_),
    .X(_01611_));
 sky130_fd_sc_hd__buf_1 _23858_ (.A(\execute.io_target_pc[21] ),
    .X(_08093_));
 sky130_fd_sc_hd__mux2_2 _23859_ (.A0(_08093_),
    .A1(\fetch.bht.bhtTable_target_pc[15][21] ),
    .S(_08079_),
    .X(_08094_));
 sky130_fd_sc_hd__buf_1 _23860_ (.A(_08094_),
    .X(_01612_));
 sky130_fd_sc_hd__buf_1 _23861_ (.A(\execute.io_target_pc[22] ),
    .X(_08095_));
 sky130_fd_sc_hd__mux2_2 _23862_ (.A0(_08095_),
    .A1(\fetch.bht.bhtTable_target_pc[15][22] ),
    .S(_08079_),
    .X(_08096_));
 sky130_fd_sc_hd__buf_1 _23863_ (.A(_08096_),
    .X(_01613_));
 sky130_fd_sc_hd__buf_1 _23864_ (.A(\execute.io_target_pc[23] ),
    .X(_08097_));
 sky130_fd_sc_hd__mux2_2 _23865_ (.A0(_08097_),
    .A1(\fetch.bht.bhtTable_target_pc[15][23] ),
    .S(_08079_),
    .X(_08098_));
 sky130_fd_sc_hd__buf_1 _23866_ (.A(_08098_),
    .X(_01614_));
 sky130_fd_sc_hd__buf_1 _23867_ (.A(\execute.io_target_pc[24] ),
    .X(_08099_));
 sky130_fd_sc_hd__mux2_2 _23868_ (.A0(_08099_),
    .A1(\fetch.bht.bhtTable_target_pc[15][24] ),
    .S(_07940_),
    .X(_08100_));
 sky130_fd_sc_hd__buf_1 _23869_ (.A(_08100_),
    .X(_01615_));
 sky130_fd_sc_hd__buf_1 _23870_ (.A(\execute.io_target_pc[25] ),
    .X(_08101_));
 sky130_fd_sc_hd__mux2_2 _23871_ (.A0(_08101_),
    .A1(\fetch.bht.bhtTable_target_pc[15][25] ),
    .S(_07940_),
    .X(_08102_));
 sky130_fd_sc_hd__buf_1 _23872_ (.A(_08102_),
    .X(_01616_));
 sky130_fd_sc_hd__buf_1 _23873_ (.A(\execute.io_target_pc[26] ),
    .X(_08103_));
 sky130_fd_sc_hd__mux2_2 _23874_ (.A0(_08103_),
    .A1(\fetch.bht.bhtTable_target_pc[15][26] ),
    .S(_07940_),
    .X(_08104_));
 sky130_fd_sc_hd__buf_1 _23875_ (.A(_08104_),
    .X(_01617_));
 sky130_fd_sc_hd__buf_1 _23876_ (.A(\execute.io_target_pc[27] ),
    .X(_08105_));
 sky130_fd_sc_hd__mux2_2 _23877_ (.A0(_08105_),
    .A1(\fetch.bht.bhtTable_target_pc[15][27] ),
    .S(_07940_),
    .X(_08106_));
 sky130_fd_sc_hd__buf_1 _23878_ (.A(_08106_),
    .X(_01618_));
 sky130_fd_sc_hd__buf_1 _23879_ (.A(\execute.io_target_pc[28] ),
    .X(_08107_));
 sky130_fd_sc_hd__mux2_2 _23880_ (.A0(_08107_),
    .A1(\fetch.bht.bhtTable_target_pc[15][28] ),
    .S(_07940_),
    .X(_08108_));
 sky130_fd_sc_hd__buf_1 _23881_ (.A(_08108_),
    .X(_01619_));
 sky130_fd_sc_hd__buf_1 _23882_ (.A(\execute.io_target_pc[29] ),
    .X(_08109_));
 sky130_fd_sc_hd__mux2_2 _23883_ (.A0(_08109_),
    .A1(\fetch.bht.bhtTable_target_pc[15][29] ),
    .S(_07940_),
    .X(_08110_));
 sky130_fd_sc_hd__buf_1 _23884_ (.A(_08110_),
    .X(_01620_));
 sky130_fd_sc_hd__buf_1 _23885_ (.A(\execute.io_target_pc[30] ),
    .X(_08111_));
 sky130_fd_sc_hd__mux2_2 _23886_ (.A0(_08111_),
    .A1(\fetch.bht.bhtTable_target_pc[15][30] ),
    .S(_07940_),
    .X(_08112_));
 sky130_fd_sc_hd__buf_1 _23887_ (.A(_08112_),
    .X(_01621_));
 sky130_fd_sc_hd__buf_1 _23888_ (.A(\execute.io_target_pc[31] ),
    .X(_08113_));
 sky130_fd_sc_hd__mux2_2 _23889_ (.A0(_08113_),
    .A1(\fetch.bht.bhtTable_target_pc[15][31] ),
    .S(_07940_),
    .X(_08114_));
 sky130_fd_sc_hd__buf_1 _23890_ (.A(_08114_),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_2 _23891_ (.A0(\fetch.bht.bhtTable_target_pc[1][0] ),
    .A1(_08049_),
    .S(_06179_),
    .X(_08115_));
 sky130_fd_sc_hd__buf_1 _23892_ (.A(_08115_),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_2 _23893_ (.A0(\fetch.bht.bhtTable_target_pc[1][1] ),
    .A1(_08051_),
    .S(_06179_),
    .X(_08116_));
 sky130_fd_sc_hd__buf_1 _23894_ (.A(_08116_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_2 _23895_ (.A0(\fetch.bht.bhtTable_target_pc[1][2] ),
    .A1(_08053_),
    .S(_06179_),
    .X(_08117_));
 sky130_fd_sc_hd__buf_1 _23896_ (.A(_08117_),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_2 _23897_ (.A0(\fetch.bht.bhtTable_target_pc[1][3] ),
    .A1(_08055_),
    .S(_06179_),
    .X(_08118_));
 sky130_fd_sc_hd__buf_1 _23898_ (.A(_08118_),
    .X(_01626_));
 sky130_fd_sc_hd__buf_1 _23899_ (.A(_06155_),
    .X(_08119_));
 sky130_fd_sc_hd__mux2_2 _23900_ (.A0(\fetch.bht.bhtTable_target_pc[1][4] ),
    .A1(_08057_),
    .S(_08119_),
    .X(_08120_));
 sky130_fd_sc_hd__buf_1 _23901_ (.A(_08120_),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_2 _23902_ (.A0(\fetch.bht.bhtTable_target_pc[1][5] ),
    .A1(_08060_),
    .S(_08119_),
    .X(_08121_));
 sky130_fd_sc_hd__buf_1 _23903_ (.A(_08121_),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_2 _23904_ (.A0(\fetch.bht.bhtTable_target_pc[1][6] ),
    .A1(_08062_),
    .S(_08119_),
    .X(_08122_));
 sky130_fd_sc_hd__buf_1 _23905_ (.A(_08122_),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_2 _23906_ (.A0(\fetch.bht.bhtTable_target_pc[1][7] ),
    .A1(_08064_),
    .S(_08119_),
    .X(_08123_));
 sky130_fd_sc_hd__buf_1 _23907_ (.A(_08123_),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_2 _23908_ (.A0(\fetch.bht.bhtTable_target_pc[1][8] ),
    .A1(_08066_),
    .S(_08119_),
    .X(_08124_));
 sky130_fd_sc_hd__buf_1 _23909_ (.A(_08124_),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_2 _23910_ (.A0(\fetch.bht.bhtTable_target_pc[1][9] ),
    .A1(_08068_),
    .S(_08119_),
    .X(_08125_));
 sky130_fd_sc_hd__buf_1 _23911_ (.A(_08125_),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_2 _23912_ (.A0(\fetch.bht.bhtTable_target_pc[1][10] ),
    .A1(_08070_),
    .S(_08119_),
    .X(_08126_));
 sky130_fd_sc_hd__buf_1 _23913_ (.A(_08126_),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_2 _23914_ (.A0(\fetch.bht.bhtTable_target_pc[1][11] ),
    .A1(_08072_),
    .S(_08119_),
    .X(_08127_));
 sky130_fd_sc_hd__buf_1 _23915_ (.A(_08127_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_2 _23916_ (.A0(\fetch.bht.bhtTable_target_pc[1][12] ),
    .A1(_08074_),
    .S(_08119_),
    .X(_08128_));
 sky130_fd_sc_hd__buf_1 _23917_ (.A(_08128_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_2 _23918_ (.A0(\fetch.bht.bhtTable_target_pc[1][13] ),
    .A1(_08076_),
    .S(_08119_),
    .X(_08129_));
 sky130_fd_sc_hd__buf_1 _23919_ (.A(_08129_),
    .X(_01636_));
 sky130_fd_sc_hd__buf_1 _23920_ (.A(_06155_),
    .X(_08130_));
 sky130_fd_sc_hd__mux2_2 _23921_ (.A0(\fetch.bht.bhtTable_target_pc[1][14] ),
    .A1(_08078_),
    .S(_08130_),
    .X(_08131_));
 sky130_fd_sc_hd__buf_1 _23922_ (.A(_08131_),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_2 _23923_ (.A0(\fetch.bht.bhtTable_target_pc[1][15] ),
    .A1(_08081_),
    .S(_08130_),
    .X(_08132_));
 sky130_fd_sc_hd__buf_1 _23924_ (.A(_08132_),
    .X(_01638_));
 sky130_fd_sc_hd__mux2_2 _23925_ (.A0(\fetch.bht.bhtTable_target_pc[1][16] ),
    .A1(_08083_),
    .S(_08130_),
    .X(_08133_));
 sky130_fd_sc_hd__buf_1 _23926_ (.A(_08133_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_2 _23927_ (.A0(\fetch.bht.bhtTable_target_pc[1][17] ),
    .A1(_08085_),
    .S(_08130_),
    .X(_08134_));
 sky130_fd_sc_hd__buf_1 _23928_ (.A(_08134_),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_2 _23929_ (.A0(\fetch.bht.bhtTable_target_pc[1][18] ),
    .A1(_08087_),
    .S(_08130_),
    .X(_08135_));
 sky130_fd_sc_hd__buf_1 _23930_ (.A(_08135_),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_2 _23931_ (.A0(\fetch.bht.bhtTable_target_pc[1][19] ),
    .A1(_08089_),
    .S(_08130_),
    .X(_08136_));
 sky130_fd_sc_hd__buf_1 _23932_ (.A(_08136_),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_2 _23933_ (.A0(\fetch.bht.bhtTable_target_pc[1][20] ),
    .A1(_08091_),
    .S(_08130_),
    .X(_08137_));
 sky130_fd_sc_hd__buf_1 _23934_ (.A(_08137_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_2 _23935_ (.A0(\fetch.bht.bhtTable_target_pc[1][21] ),
    .A1(_08093_),
    .S(_08130_),
    .X(_08138_));
 sky130_fd_sc_hd__buf_1 _23936_ (.A(_08138_),
    .X(_01644_));
 sky130_fd_sc_hd__mux2_2 _23937_ (.A0(\fetch.bht.bhtTable_target_pc[1][22] ),
    .A1(_08095_),
    .S(_08130_),
    .X(_08139_));
 sky130_fd_sc_hd__buf_1 _23938_ (.A(_08139_),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_2 _23939_ (.A0(\fetch.bht.bhtTable_target_pc[1][23] ),
    .A1(_08097_),
    .S(_08130_),
    .X(_08140_));
 sky130_fd_sc_hd__buf_1 _23940_ (.A(_08140_),
    .X(_01646_));
 sky130_fd_sc_hd__mux2_2 _23941_ (.A0(\fetch.bht.bhtTable_target_pc[1][24] ),
    .A1(_08099_),
    .S(_06156_),
    .X(_08141_));
 sky130_fd_sc_hd__buf_1 _23942_ (.A(_08141_),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_2 _23943_ (.A0(\fetch.bht.bhtTable_target_pc[1][25] ),
    .A1(_08101_),
    .S(_06156_),
    .X(_08142_));
 sky130_fd_sc_hd__buf_1 _23944_ (.A(_08142_),
    .X(_01648_));
 sky130_fd_sc_hd__mux2_2 _23945_ (.A0(\fetch.bht.bhtTable_target_pc[1][26] ),
    .A1(_08103_),
    .S(_06156_),
    .X(_08143_));
 sky130_fd_sc_hd__buf_1 _23946_ (.A(_08143_),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_2 _23947_ (.A0(\fetch.bht.bhtTable_target_pc[1][27] ),
    .A1(_08105_),
    .S(_06156_),
    .X(_08144_));
 sky130_fd_sc_hd__buf_1 _23948_ (.A(_08144_),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_2 _23949_ (.A0(\fetch.bht.bhtTable_target_pc[1][28] ),
    .A1(_08107_),
    .S(_06156_),
    .X(_08145_));
 sky130_fd_sc_hd__buf_1 _23950_ (.A(_08145_),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_2 _23951_ (.A0(\fetch.bht.bhtTable_target_pc[1][29] ),
    .A1(_08109_),
    .S(_06156_),
    .X(_08146_));
 sky130_fd_sc_hd__buf_1 _23952_ (.A(_08146_),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_2 _23953_ (.A0(\fetch.bht.bhtTable_target_pc[1][30] ),
    .A1(_08111_),
    .S(_06156_),
    .X(_08147_));
 sky130_fd_sc_hd__buf_1 _23954_ (.A(_08147_),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_2 _23955_ (.A0(\fetch.bht.bhtTable_target_pc[1][31] ),
    .A1(_08113_),
    .S(_06156_),
    .X(_08148_));
 sky130_fd_sc_hd__buf_1 _23956_ (.A(_08148_),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_2 _23957_ (.A0(\fetch.bht.bhtTable_target_pc[2][0] ),
    .A1(\execute.io_target_pc[0] ),
    .S(_07983_),
    .X(_08149_));
 sky130_fd_sc_hd__buf_1 _23958_ (.A(_08149_),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_2 _23959_ (.A0(\fetch.bht.bhtTable_target_pc[2][1] ),
    .A1(\execute.io_target_pc[1] ),
    .S(_07983_),
    .X(_08150_));
 sky130_fd_sc_hd__buf_1 _23960_ (.A(_08150_),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_2 _23961_ (.A0(\fetch.bht.bhtTable_target_pc[2][2] ),
    .A1(\execute.io_target_pc[2] ),
    .S(_07983_),
    .X(_08151_));
 sky130_fd_sc_hd__buf_1 _23962_ (.A(_08151_),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_2 _23963_ (.A0(\fetch.bht.bhtTable_target_pc[2][3] ),
    .A1(\execute.io_target_pc[3] ),
    .S(_07983_),
    .X(_08152_));
 sky130_fd_sc_hd__buf_1 _23964_ (.A(_08152_),
    .X(_01658_));
 sky130_fd_sc_hd__buf_1 _23965_ (.A(_07959_),
    .X(_08153_));
 sky130_fd_sc_hd__mux2_2 _23966_ (.A0(\fetch.bht.bhtTable_target_pc[2][4] ),
    .A1(\execute.io_target_pc[4] ),
    .S(_08153_),
    .X(_08154_));
 sky130_fd_sc_hd__buf_1 _23967_ (.A(_08154_),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_2 _23968_ (.A0(\fetch.bht.bhtTable_target_pc[2][5] ),
    .A1(\execute.io_target_pc[5] ),
    .S(_08153_),
    .X(_08155_));
 sky130_fd_sc_hd__buf_1 _23969_ (.A(_08155_),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_2 _23970_ (.A0(\fetch.bht.bhtTable_target_pc[2][6] ),
    .A1(\execute.io_target_pc[6] ),
    .S(_08153_),
    .X(_08156_));
 sky130_fd_sc_hd__buf_1 _23971_ (.A(_08156_),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_2 _23972_ (.A0(\fetch.bht.bhtTable_target_pc[2][7] ),
    .A1(\execute.io_target_pc[7] ),
    .S(_08153_),
    .X(_08157_));
 sky130_fd_sc_hd__buf_1 _23973_ (.A(_08157_),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_2 _23974_ (.A0(\fetch.bht.bhtTable_target_pc[2][8] ),
    .A1(\execute.io_target_pc[8] ),
    .S(_08153_),
    .X(_08158_));
 sky130_fd_sc_hd__buf_1 _23975_ (.A(_08158_),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_2 _23976_ (.A0(\fetch.bht.bhtTable_target_pc[2][9] ),
    .A1(\execute.io_target_pc[9] ),
    .S(_08153_),
    .X(_08159_));
 sky130_fd_sc_hd__buf_1 _23977_ (.A(_08159_),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_2 _23978_ (.A0(\fetch.bht.bhtTable_target_pc[2][10] ),
    .A1(\execute.io_target_pc[10] ),
    .S(_08153_),
    .X(_08160_));
 sky130_fd_sc_hd__buf_1 _23979_ (.A(_08160_),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_2 _23980_ (.A0(\fetch.bht.bhtTable_target_pc[2][11] ),
    .A1(\execute.io_target_pc[11] ),
    .S(_08153_),
    .X(_08161_));
 sky130_fd_sc_hd__buf_1 _23981_ (.A(_08161_),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_2 _23982_ (.A0(\fetch.bht.bhtTable_target_pc[2][12] ),
    .A1(\execute.io_target_pc[12] ),
    .S(_08153_),
    .X(_08162_));
 sky130_fd_sc_hd__buf_1 _23983_ (.A(_08162_),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_2 _23984_ (.A0(\fetch.bht.bhtTable_target_pc[2][13] ),
    .A1(\execute.io_target_pc[13] ),
    .S(_08153_),
    .X(_08163_));
 sky130_fd_sc_hd__buf_1 _23985_ (.A(_08163_),
    .X(_01668_));
 sky130_fd_sc_hd__buf_1 _23986_ (.A(_07959_),
    .X(_08164_));
 sky130_fd_sc_hd__mux2_2 _23987_ (.A0(\fetch.bht.bhtTable_target_pc[2][14] ),
    .A1(\execute.io_target_pc[14] ),
    .S(_08164_),
    .X(_08165_));
 sky130_fd_sc_hd__buf_1 _23988_ (.A(_08165_),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_2 _23989_ (.A0(\fetch.bht.bhtTable_target_pc[2][15] ),
    .A1(\execute.io_target_pc[15] ),
    .S(_08164_),
    .X(_08166_));
 sky130_fd_sc_hd__buf_1 _23990_ (.A(_08166_),
    .X(_01670_));
 sky130_fd_sc_hd__mux2_2 _23991_ (.A0(\fetch.bht.bhtTable_target_pc[2][16] ),
    .A1(\execute.io_target_pc[16] ),
    .S(_08164_),
    .X(_08167_));
 sky130_fd_sc_hd__buf_1 _23992_ (.A(_08167_),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_2 _23993_ (.A0(\fetch.bht.bhtTable_target_pc[2][17] ),
    .A1(\execute.io_target_pc[17] ),
    .S(_08164_),
    .X(_08168_));
 sky130_fd_sc_hd__buf_1 _23994_ (.A(_08168_),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_2 _23995_ (.A0(\fetch.bht.bhtTable_target_pc[2][18] ),
    .A1(\execute.io_target_pc[18] ),
    .S(_08164_),
    .X(_08169_));
 sky130_fd_sc_hd__buf_1 _23996_ (.A(_08169_),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_2 _23997_ (.A0(\fetch.bht.bhtTable_target_pc[2][19] ),
    .A1(\execute.io_target_pc[19] ),
    .S(_08164_),
    .X(_08170_));
 sky130_fd_sc_hd__buf_1 _23998_ (.A(_08170_),
    .X(_01674_));
 sky130_fd_sc_hd__mux2_2 _23999_ (.A0(\fetch.bht.bhtTable_target_pc[2][20] ),
    .A1(\execute.io_target_pc[20] ),
    .S(_08164_),
    .X(_08171_));
 sky130_fd_sc_hd__buf_1 _24000_ (.A(_08171_),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_2 _24001_ (.A0(\fetch.bht.bhtTable_target_pc[2][21] ),
    .A1(\execute.io_target_pc[21] ),
    .S(_08164_),
    .X(_08172_));
 sky130_fd_sc_hd__buf_1 _24002_ (.A(_08172_),
    .X(_01676_));
 sky130_fd_sc_hd__mux2_2 _24003_ (.A0(\fetch.bht.bhtTable_target_pc[2][22] ),
    .A1(\execute.io_target_pc[22] ),
    .S(_08164_),
    .X(_08173_));
 sky130_fd_sc_hd__buf_1 _24004_ (.A(_08173_),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_2 _24005_ (.A0(\fetch.bht.bhtTable_target_pc[2][23] ),
    .A1(\execute.io_target_pc[23] ),
    .S(_08164_),
    .X(_08174_));
 sky130_fd_sc_hd__buf_1 _24006_ (.A(_08174_),
    .X(_01678_));
 sky130_fd_sc_hd__mux2_2 _24007_ (.A0(\fetch.bht.bhtTable_target_pc[2][24] ),
    .A1(\execute.io_target_pc[24] ),
    .S(_07960_),
    .X(_08175_));
 sky130_fd_sc_hd__buf_1 _24008_ (.A(_08175_),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_2 _24009_ (.A0(\fetch.bht.bhtTable_target_pc[2][25] ),
    .A1(\execute.io_target_pc[25] ),
    .S(_07960_),
    .X(_08176_));
 sky130_fd_sc_hd__buf_1 _24010_ (.A(_08176_),
    .X(_01680_));
 sky130_fd_sc_hd__mux2_2 _24011_ (.A0(\fetch.bht.bhtTable_target_pc[2][26] ),
    .A1(\execute.io_target_pc[26] ),
    .S(_07960_),
    .X(_08177_));
 sky130_fd_sc_hd__buf_1 _24012_ (.A(_08177_),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_2 _24013_ (.A0(\fetch.bht.bhtTable_target_pc[2][27] ),
    .A1(\execute.io_target_pc[27] ),
    .S(_07960_),
    .X(_08178_));
 sky130_fd_sc_hd__buf_1 _24014_ (.A(_08178_),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_2 _24015_ (.A0(\fetch.bht.bhtTable_target_pc[2][28] ),
    .A1(\execute.io_target_pc[28] ),
    .S(_07960_),
    .X(_08179_));
 sky130_fd_sc_hd__buf_1 _24016_ (.A(_08179_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_2 _24017_ (.A0(\fetch.bht.bhtTable_target_pc[2][29] ),
    .A1(\execute.io_target_pc[29] ),
    .S(_07960_),
    .X(_08180_));
 sky130_fd_sc_hd__buf_1 _24018_ (.A(_08180_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_2 _24019_ (.A0(\fetch.bht.bhtTable_target_pc[2][30] ),
    .A1(\execute.io_target_pc[30] ),
    .S(_07960_),
    .X(_08181_));
 sky130_fd_sc_hd__buf_1 _24020_ (.A(_08181_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_2 _24021_ (.A0(\fetch.bht.bhtTable_target_pc[2][31] ),
    .A1(\execute.io_target_pc[31] ),
    .S(_07960_),
    .X(_08182_));
 sky130_fd_sc_hd__buf_1 _24022_ (.A(_08182_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_2 _24023_ (.A0(\fetch.bht.bhtTable_target_pc[3][0] ),
    .A1(\execute.io_target_pc[0] ),
    .S(_08014_),
    .X(_08183_));
 sky130_fd_sc_hd__buf_1 _24024_ (.A(_08183_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_2 _24025_ (.A0(\fetch.bht.bhtTable_target_pc[3][1] ),
    .A1(\execute.io_target_pc[1] ),
    .S(_08014_),
    .X(_08184_));
 sky130_fd_sc_hd__buf_1 _24026_ (.A(_08184_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_2 _24027_ (.A0(\fetch.bht.bhtTable_target_pc[3][2] ),
    .A1(\execute.io_target_pc[2] ),
    .S(_08014_),
    .X(_08185_));
 sky130_fd_sc_hd__buf_1 _24028_ (.A(_08185_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_2 _24029_ (.A0(\fetch.bht.bhtTable_target_pc[3][3] ),
    .A1(\execute.io_target_pc[3] ),
    .S(_08014_),
    .X(_08186_));
 sky130_fd_sc_hd__buf_1 _24030_ (.A(_08186_),
    .X(_01690_));
 sky130_fd_sc_hd__buf_1 _24031_ (.A(_07990_),
    .X(_08187_));
 sky130_fd_sc_hd__mux2_2 _24032_ (.A0(\fetch.bht.bhtTable_target_pc[3][4] ),
    .A1(\execute.io_target_pc[4] ),
    .S(_08187_),
    .X(_08188_));
 sky130_fd_sc_hd__buf_1 _24033_ (.A(_08188_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_2 _24034_ (.A0(\fetch.bht.bhtTable_target_pc[3][5] ),
    .A1(\execute.io_target_pc[5] ),
    .S(_08187_),
    .X(_08189_));
 sky130_fd_sc_hd__buf_1 _24035_ (.A(_08189_),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_2 _24036_ (.A0(\fetch.bht.bhtTable_target_pc[3][6] ),
    .A1(\execute.io_target_pc[6] ),
    .S(_08187_),
    .X(_08190_));
 sky130_fd_sc_hd__buf_1 _24037_ (.A(_08190_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_2 _24038_ (.A0(\fetch.bht.bhtTable_target_pc[3][7] ),
    .A1(\execute.io_target_pc[7] ),
    .S(_08187_),
    .X(_08191_));
 sky130_fd_sc_hd__buf_1 _24039_ (.A(_08191_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_2 _24040_ (.A0(\fetch.bht.bhtTable_target_pc[3][8] ),
    .A1(\execute.io_target_pc[8] ),
    .S(_08187_),
    .X(_08192_));
 sky130_fd_sc_hd__buf_1 _24041_ (.A(_08192_),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_2 _24042_ (.A0(\fetch.bht.bhtTable_target_pc[3][9] ),
    .A1(\execute.io_target_pc[9] ),
    .S(_08187_),
    .X(_08193_));
 sky130_fd_sc_hd__buf_1 _24043_ (.A(_08193_),
    .X(_01696_));
 sky130_fd_sc_hd__mux2_2 _24044_ (.A0(\fetch.bht.bhtTable_target_pc[3][10] ),
    .A1(\execute.io_target_pc[10] ),
    .S(_08187_),
    .X(_08194_));
 sky130_fd_sc_hd__buf_1 _24045_ (.A(_08194_),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_2 _24046_ (.A0(\fetch.bht.bhtTable_target_pc[3][11] ),
    .A1(\execute.io_target_pc[11] ),
    .S(_08187_),
    .X(_08195_));
 sky130_fd_sc_hd__buf_1 _24047_ (.A(_08195_),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_2 _24048_ (.A0(\fetch.bht.bhtTable_target_pc[3][12] ),
    .A1(\execute.io_target_pc[12] ),
    .S(_08187_),
    .X(_08196_));
 sky130_fd_sc_hd__buf_1 _24049_ (.A(_08196_),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_2 _24050_ (.A0(\fetch.bht.bhtTable_target_pc[3][13] ),
    .A1(\execute.io_target_pc[13] ),
    .S(_08187_),
    .X(_08197_));
 sky130_fd_sc_hd__buf_1 _24051_ (.A(_08197_),
    .X(_01700_));
 sky130_fd_sc_hd__buf_1 _24052_ (.A(_07990_),
    .X(_08198_));
 sky130_fd_sc_hd__mux2_2 _24053_ (.A0(\fetch.bht.bhtTable_target_pc[3][14] ),
    .A1(\execute.io_target_pc[14] ),
    .S(_08198_),
    .X(_08199_));
 sky130_fd_sc_hd__buf_1 _24054_ (.A(_08199_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_2 _24055_ (.A0(\fetch.bht.bhtTable_target_pc[3][15] ),
    .A1(\execute.io_target_pc[15] ),
    .S(_08198_),
    .X(_08200_));
 sky130_fd_sc_hd__buf_1 _24056_ (.A(_08200_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_2 _24057_ (.A0(\fetch.bht.bhtTable_target_pc[3][16] ),
    .A1(\execute.io_target_pc[16] ),
    .S(_08198_),
    .X(_08201_));
 sky130_fd_sc_hd__buf_1 _24058_ (.A(_08201_),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_2 _24059_ (.A0(\fetch.bht.bhtTable_target_pc[3][17] ),
    .A1(\execute.io_target_pc[17] ),
    .S(_08198_),
    .X(_08202_));
 sky130_fd_sc_hd__buf_1 _24060_ (.A(_08202_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_2 _24061_ (.A0(\fetch.bht.bhtTable_target_pc[3][18] ),
    .A1(\execute.io_target_pc[18] ),
    .S(_08198_),
    .X(_08203_));
 sky130_fd_sc_hd__buf_1 _24062_ (.A(_08203_),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_2 _24063_ (.A0(\fetch.bht.bhtTable_target_pc[3][19] ),
    .A1(\execute.io_target_pc[19] ),
    .S(_08198_),
    .X(_08204_));
 sky130_fd_sc_hd__buf_1 _24064_ (.A(_08204_),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_2 _24065_ (.A0(\fetch.bht.bhtTable_target_pc[3][20] ),
    .A1(\execute.io_target_pc[20] ),
    .S(_08198_),
    .X(_08205_));
 sky130_fd_sc_hd__buf_1 _24066_ (.A(_08205_),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_2 _24067_ (.A0(\fetch.bht.bhtTable_target_pc[3][21] ),
    .A1(\execute.io_target_pc[21] ),
    .S(_08198_),
    .X(_08206_));
 sky130_fd_sc_hd__buf_1 _24068_ (.A(_08206_),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_2 _24069_ (.A0(\fetch.bht.bhtTable_target_pc[3][22] ),
    .A1(\execute.io_target_pc[22] ),
    .S(_08198_),
    .X(_08207_));
 sky130_fd_sc_hd__buf_1 _24070_ (.A(_08207_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_2 _24071_ (.A0(\fetch.bht.bhtTable_target_pc[3][23] ),
    .A1(\execute.io_target_pc[23] ),
    .S(_08198_),
    .X(_08208_));
 sky130_fd_sc_hd__buf_1 _24072_ (.A(_08208_),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_2 _24073_ (.A0(\fetch.bht.bhtTable_target_pc[3][24] ),
    .A1(\execute.io_target_pc[24] ),
    .S(_07991_),
    .X(_08209_));
 sky130_fd_sc_hd__buf_1 _24074_ (.A(_08209_),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_2 _24075_ (.A0(\fetch.bht.bhtTable_target_pc[3][25] ),
    .A1(\execute.io_target_pc[25] ),
    .S(_07991_),
    .X(_08210_));
 sky130_fd_sc_hd__buf_1 _24076_ (.A(_08210_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_2 _24077_ (.A0(\fetch.bht.bhtTable_target_pc[3][26] ),
    .A1(\execute.io_target_pc[26] ),
    .S(_07991_),
    .X(_08211_));
 sky130_fd_sc_hd__buf_1 _24078_ (.A(_08211_),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_2 _24079_ (.A0(\fetch.bht.bhtTable_target_pc[3][27] ),
    .A1(\execute.io_target_pc[27] ),
    .S(_07991_),
    .X(_08212_));
 sky130_fd_sc_hd__buf_1 _24080_ (.A(_08212_),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_2 _24081_ (.A0(\fetch.bht.bhtTable_target_pc[3][28] ),
    .A1(\execute.io_target_pc[28] ),
    .S(_07991_),
    .X(_08213_));
 sky130_fd_sc_hd__buf_1 _24082_ (.A(_08213_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_2 _24083_ (.A0(\fetch.bht.bhtTable_target_pc[3][29] ),
    .A1(\execute.io_target_pc[29] ),
    .S(_07991_),
    .X(_08214_));
 sky130_fd_sc_hd__buf_1 _24084_ (.A(_08214_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_2 _24085_ (.A0(\fetch.bht.bhtTable_target_pc[3][30] ),
    .A1(\execute.io_target_pc[30] ),
    .S(_07991_),
    .X(_08215_));
 sky130_fd_sc_hd__buf_1 _24086_ (.A(_08215_),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_2 _24087_ (.A0(\fetch.bht.bhtTable_target_pc[3][31] ),
    .A1(\execute.io_target_pc[31] ),
    .S(_07991_),
    .X(_08216_));
 sky130_fd_sc_hd__buf_1 _24088_ (.A(_08216_),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_2 _24089_ (.A0(\fetch.bht.bhtTable_target_pc[4][0] ),
    .A1(\execute.io_target_pc[0] ),
    .S(_06450_),
    .X(_08217_));
 sky130_fd_sc_hd__buf_1 _24090_ (.A(_08217_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_2 _24091_ (.A0(\fetch.bht.bhtTable_target_pc[4][1] ),
    .A1(\execute.io_target_pc[1] ),
    .S(_06450_),
    .X(_08218_));
 sky130_fd_sc_hd__buf_1 _24092_ (.A(_08218_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_2 _24093_ (.A0(\fetch.bht.bhtTable_target_pc[4][2] ),
    .A1(\execute.io_target_pc[2] ),
    .S(_06450_),
    .X(_08219_));
 sky130_fd_sc_hd__buf_1 _24094_ (.A(_08219_),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_2 _24095_ (.A0(\fetch.bht.bhtTable_target_pc[4][3] ),
    .A1(\execute.io_target_pc[3] ),
    .S(_06450_),
    .X(_08220_));
 sky130_fd_sc_hd__buf_1 _24096_ (.A(_08220_),
    .X(_01722_));
 sky130_fd_sc_hd__buf_1 _24097_ (.A(_06426_),
    .X(_08221_));
 sky130_fd_sc_hd__mux2_2 _24098_ (.A0(\fetch.bht.bhtTable_target_pc[4][4] ),
    .A1(\execute.io_target_pc[4] ),
    .S(_08221_),
    .X(_08222_));
 sky130_fd_sc_hd__buf_1 _24099_ (.A(_08222_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_2 _24100_ (.A0(\fetch.bht.bhtTable_target_pc[4][5] ),
    .A1(\execute.io_target_pc[5] ),
    .S(_08221_),
    .X(_08223_));
 sky130_fd_sc_hd__buf_1 _24101_ (.A(_08223_),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_2 _24102_ (.A0(\fetch.bht.bhtTable_target_pc[4][6] ),
    .A1(\execute.io_target_pc[6] ),
    .S(_08221_),
    .X(_08224_));
 sky130_fd_sc_hd__buf_1 _24103_ (.A(_08224_),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_2 _24104_ (.A0(\fetch.bht.bhtTable_target_pc[4][7] ),
    .A1(\execute.io_target_pc[7] ),
    .S(_08221_),
    .X(_08225_));
 sky130_fd_sc_hd__buf_1 _24105_ (.A(_08225_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_2 _24106_ (.A0(\fetch.bht.bhtTable_target_pc[4][8] ),
    .A1(\execute.io_target_pc[8] ),
    .S(_08221_),
    .X(_08226_));
 sky130_fd_sc_hd__buf_1 _24107_ (.A(_08226_),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_2 _24108_ (.A0(\fetch.bht.bhtTable_target_pc[4][9] ),
    .A1(\execute.io_target_pc[9] ),
    .S(_08221_),
    .X(_08227_));
 sky130_fd_sc_hd__buf_1 _24109_ (.A(_08227_),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_2 _24110_ (.A0(\fetch.bht.bhtTable_target_pc[4][10] ),
    .A1(\execute.io_target_pc[10] ),
    .S(_08221_),
    .X(_08228_));
 sky130_fd_sc_hd__buf_1 _24111_ (.A(_08228_),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_2 _24112_ (.A0(\fetch.bht.bhtTable_target_pc[4][11] ),
    .A1(\execute.io_target_pc[11] ),
    .S(_08221_),
    .X(_08229_));
 sky130_fd_sc_hd__buf_1 _24113_ (.A(_08229_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_2 _24114_ (.A0(\fetch.bht.bhtTable_target_pc[4][12] ),
    .A1(\execute.io_target_pc[12] ),
    .S(_08221_),
    .X(_08230_));
 sky130_fd_sc_hd__buf_1 _24115_ (.A(_08230_),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_2 _24116_ (.A0(\fetch.bht.bhtTable_target_pc[4][13] ),
    .A1(\execute.io_target_pc[13] ),
    .S(_08221_),
    .X(_08231_));
 sky130_fd_sc_hd__buf_1 _24117_ (.A(_08231_),
    .X(_01732_));
 sky130_fd_sc_hd__buf_1 _24118_ (.A(_06426_),
    .X(_08232_));
 sky130_fd_sc_hd__mux2_2 _24119_ (.A0(\fetch.bht.bhtTable_target_pc[4][14] ),
    .A1(\execute.io_target_pc[14] ),
    .S(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__buf_1 _24120_ (.A(_08233_),
    .X(_01733_));
 sky130_fd_sc_hd__mux2_2 _24121_ (.A0(\fetch.bht.bhtTable_target_pc[4][15] ),
    .A1(\execute.io_target_pc[15] ),
    .S(_08232_),
    .X(_08234_));
 sky130_fd_sc_hd__buf_1 _24122_ (.A(_08234_),
    .X(_01734_));
 sky130_fd_sc_hd__mux2_2 _24123_ (.A0(\fetch.bht.bhtTable_target_pc[4][16] ),
    .A1(\execute.io_target_pc[16] ),
    .S(_08232_),
    .X(_08235_));
 sky130_fd_sc_hd__buf_1 _24124_ (.A(_08235_),
    .X(_01735_));
 sky130_fd_sc_hd__mux2_2 _24125_ (.A0(\fetch.bht.bhtTable_target_pc[4][17] ),
    .A1(\execute.io_target_pc[17] ),
    .S(_08232_),
    .X(_08236_));
 sky130_fd_sc_hd__buf_1 _24126_ (.A(_08236_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_2 _24127_ (.A0(\fetch.bht.bhtTable_target_pc[4][18] ),
    .A1(\execute.io_target_pc[18] ),
    .S(_08232_),
    .X(_08237_));
 sky130_fd_sc_hd__buf_1 _24128_ (.A(_08237_),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_2 _24129_ (.A0(\fetch.bht.bhtTable_target_pc[4][19] ),
    .A1(\execute.io_target_pc[19] ),
    .S(_08232_),
    .X(_08238_));
 sky130_fd_sc_hd__buf_1 _24130_ (.A(_08238_),
    .X(_01738_));
 sky130_fd_sc_hd__mux2_2 _24131_ (.A0(\fetch.bht.bhtTable_target_pc[4][20] ),
    .A1(\execute.io_target_pc[20] ),
    .S(_08232_),
    .X(_08239_));
 sky130_fd_sc_hd__buf_1 _24132_ (.A(_08239_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_2 _24133_ (.A0(\fetch.bht.bhtTable_target_pc[4][21] ),
    .A1(\execute.io_target_pc[21] ),
    .S(_08232_),
    .X(_08240_));
 sky130_fd_sc_hd__buf_1 _24134_ (.A(_08240_),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_2 _24135_ (.A0(\fetch.bht.bhtTable_target_pc[4][22] ),
    .A1(\execute.io_target_pc[22] ),
    .S(_08232_),
    .X(_08241_));
 sky130_fd_sc_hd__buf_1 _24136_ (.A(_08241_),
    .X(_01741_));
 sky130_fd_sc_hd__mux2_2 _24137_ (.A0(\fetch.bht.bhtTable_target_pc[4][23] ),
    .A1(\execute.io_target_pc[23] ),
    .S(_08232_),
    .X(_08242_));
 sky130_fd_sc_hd__buf_1 _24138_ (.A(_08242_),
    .X(_01742_));
 sky130_fd_sc_hd__mux2_2 _24139_ (.A0(\fetch.bht.bhtTable_target_pc[4][24] ),
    .A1(\execute.io_target_pc[24] ),
    .S(_06427_),
    .X(_08243_));
 sky130_fd_sc_hd__buf_1 _24140_ (.A(_08243_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_2 _24141_ (.A0(\fetch.bht.bhtTable_target_pc[4][25] ),
    .A1(\execute.io_target_pc[25] ),
    .S(_06427_),
    .X(_08244_));
 sky130_fd_sc_hd__buf_1 _24142_ (.A(_08244_),
    .X(_01744_));
 sky130_fd_sc_hd__mux2_2 _24143_ (.A0(\fetch.bht.bhtTable_target_pc[4][26] ),
    .A1(\execute.io_target_pc[26] ),
    .S(_06427_),
    .X(_08245_));
 sky130_fd_sc_hd__buf_1 _24144_ (.A(_08245_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_2 _24145_ (.A0(\fetch.bht.bhtTable_target_pc[4][27] ),
    .A1(\execute.io_target_pc[27] ),
    .S(_06427_),
    .X(_08246_));
 sky130_fd_sc_hd__buf_1 _24146_ (.A(_08246_),
    .X(_01746_));
 sky130_fd_sc_hd__mux2_2 _24147_ (.A0(\fetch.bht.bhtTable_target_pc[4][28] ),
    .A1(\execute.io_target_pc[28] ),
    .S(_06427_),
    .X(_08247_));
 sky130_fd_sc_hd__buf_1 _24148_ (.A(_08247_),
    .X(_01747_));
 sky130_fd_sc_hd__mux2_2 _24149_ (.A0(\fetch.bht.bhtTable_target_pc[4][29] ),
    .A1(\execute.io_target_pc[29] ),
    .S(_06427_),
    .X(_08248_));
 sky130_fd_sc_hd__buf_1 _24150_ (.A(_08248_),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_2 _24151_ (.A0(\fetch.bht.bhtTable_target_pc[4][30] ),
    .A1(\execute.io_target_pc[30] ),
    .S(_06427_),
    .X(_08249_));
 sky130_fd_sc_hd__buf_1 _24152_ (.A(_08249_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_2 _24153_ (.A0(\fetch.bht.bhtTable_target_pc[4][31] ),
    .A1(\execute.io_target_pc[31] ),
    .S(_06427_),
    .X(_08250_));
 sky130_fd_sc_hd__buf_1 _24154_ (.A(_08250_),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_2 _24155_ (.A0(_08049_),
    .A1(\fetch.bht.bhtTable_target_pc[5][0] ),
    .S(_06274_),
    .X(_08251_));
 sky130_fd_sc_hd__buf_1 _24156_ (.A(_08251_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_2 _24157_ (.A0(_08051_),
    .A1(\fetch.bht.bhtTable_target_pc[5][1] ),
    .S(_06274_),
    .X(_08252_));
 sky130_fd_sc_hd__buf_1 _24158_ (.A(_08252_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_2 _24159_ (.A0(_08053_),
    .A1(\fetch.bht.bhtTable_target_pc[5][2] ),
    .S(_06274_),
    .X(_08253_));
 sky130_fd_sc_hd__buf_1 _24160_ (.A(_08253_),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_2 _24161_ (.A0(_08055_),
    .A1(\fetch.bht.bhtTable_target_pc[5][3] ),
    .S(_06274_),
    .X(_08254_));
 sky130_fd_sc_hd__buf_1 _24162_ (.A(_08254_),
    .X(_01754_));
 sky130_fd_sc_hd__buf_1 _24163_ (.A(_06250_),
    .X(_08255_));
 sky130_fd_sc_hd__mux2_2 _24164_ (.A0(_08057_),
    .A1(\fetch.bht.bhtTable_target_pc[5][4] ),
    .S(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__buf_1 _24165_ (.A(_08256_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_2 _24166_ (.A0(_08060_),
    .A1(\fetch.bht.bhtTable_target_pc[5][5] ),
    .S(_08255_),
    .X(_08257_));
 sky130_fd_sc_hd__buf_1 _24167_ (.A(_08257_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_2 _24168_ (.A0(_08062_),
    .A1(\fetch.bht.bhtTable_target_pc[5][6] ),
    .S(_08255_),
    .X(_08258_));
 sky130_fd_sc_hd__buf_1 _24169_ (.A(_08258_),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_2 _24170_ (.A0(_08064_),
    .A1(\fetch.bht.bhtTable_target_pc[5][7] ),
    .S(_08255_),
    .X(_08259_));
 sky130_fd_sc_hd__buf_1 _24171_ (.A(_08259_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_2 _24172_ (.A0(_08066_),
    .A1(\fetch.bht.bhtTable_target_pc[5][8] ),
    .S(_08255_),
    .X(_08260_));
 sky130_fd_sc_hd__buf_1 _24173_ (.A(_08260_),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_2 _24174_ (.A0(_08068_),
    .A1(\fetch.bht.bhtTable_target_pc[5][9] ),
    .S(_08255_),
    .X(_08261_));
 sky130_fd_sc_hd__buf_1 _24175_ (.A(_08261_),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_2 _24176_ (.A0(_08070_),
    .A1(\fetch.bht.bhtTable_target_pc[5][10] ),
    .S(_08255_),
    .X(_08262_));
 sky130_fd_sc_hd__buf_1 _24177_ (.A(_08262_),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_2 _24178_ (.A0(_08072_),
    .A1(\fetch.bht.bhtTable_target_pc[5][11] ),
    .S(_08255_),
    .X(_08263_));
 sky130_fd_sc_hd__buf_1 _24179_ (.A(_08263_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_2 _24180_ (.A0(_08074_),
    .A1(\fetch.bht.bhtTable_target_pc[5][12] ),
    .S(_08255_),
    .X(_08264_));
 sky130_fd_sc_hd__buf_1 _24181_ (.A(_08264_),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_2 _24182_ (.A0(_08076_),
    .A1(\fetch.bht.bhtTable_target_pc[5][13] ),
    .S(_08255_),
    .X(_08265_));
 sky130_fd_sc_hd__buf_1 _24183_ (.A(_08265_),
    .X(_01764_));
 sky130_fd_sc_hd__buf_1 _24184_ (.A(_06250_),
    .X(_08266_));
 sky130_fd_sc_hd__mux2_2 _24185_ (.A0(_08078_),
    .A1(\fetch.bht.bhtTable_target_pc[5][14] ),
    .S(_08266_),
    .X(_08267_));
 sky130_fd_sc_hd__buf_1 _24186_ (.A(_08267_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_2 _24187_ (.A0(_08081_),
    .A1(\fetch.bht.bhtTable_target_pc[5][15] ),
    .S(_08266_),
    .X(_08268_));
 sky130_fd_sc_hd__buf_1 _24188_ (.A(_08268_),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_2 _24189_ (.A0(_08083_),
    .A1(\fetch.bht.bhtTable_target_pc[5][16] ),
    .S(_08266_),
    .X(_08269_));
 sky130_fd_sc_hd__buf_1 _24190_ (.A(_08269_),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_2 _24191_ (.A0(_08085_),
    .A1(\fetch.bht.bhtTable_target_pc[5][17] ),
    .S(_08266_),
    .X(_08270_));
 sky130_fd_sc_hd__buf_1 _24192_ (.A(_08270_),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_2 _24193_ (.A0(_08087_),
    .A1(\fetch.bht.bhtTable_target_pc[5][18] ),
    .S(_08266_),
    .X(_08271_));
 sky130_fd_sc_hd__buf_1 _24194_ (.A(_08271_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_2 _24195_ (.A0(_08089_),
    .A1(\fetch.bht.bhtTable_target_pc[5][19] ),
    .S(_08266_),
    .X(_08272_));
 sky130_fd_sc_hd__buf_1 _24196_ (.A(_08272_),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_2 _24197_ (.A0(_08091_),
    .A1(\fetch.bht.bhtTable_target_pc[5][20] ),
    .S(_08266_),
    .X(_08273_));
 sky130_fd_sc_hd__buf_1 _24198_ (.A(_08273_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_2 _24199_ (.A0(_08093_),
    .A1(\fetch.bht.bhtTable_target_pc[5][21] ),
    .S(_08266_),
    .X(_08274_));
 sky130_fd_sc_hd__buf_1 _24200_ (.A(_08274_),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_2 _24201_ (.A0(_08095_),
    .A1(\fetch.bht.bhtTable_target_pc[5][22] ),
    .S(_08266_),
    .X(_08275_));
 sky130_fd_sc_hd__buf_1 _24202_ (.A(_08275_),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_2 _24203_ (.A0(_08097_),
    .A1(\fetch.bht.bhtTable_target_pc[5][23] ),
    .S(_08266_),
    .X(_08276_));
 sky130_fd_sc_hd__buf_1 _24204_ (.A(_08276_),
    .X(_01774_));
 sky130_fd_sc_hd__mux2_2 _24205_ (.A0(_08099_),
    .A1(\fetch.bht.bhtTable_target_pc[5][24] ),
    .S(_06251_),
    .X(_08277_));
 sky130_fd_sc_hd__buf_1 _24206_ (.A(_08277_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_2 _24207_ (.A0(_08101_),
    .A1(\fetch.bht.bhtTable_target_pc[5][25] ),
    .S(_06251_),
    .X(_08278_));
 sky130_fd_sc_hd__buf_1 _24208_ (.A(_08278_),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_2 _24209_ (.A0(_08103_),
    .A1(\fetch.bht.bhtTable_target_pc[5][26] ),
    .S(_06251_),
    .X(_08279_));
 sky130_fd_sc_hd__buf_1 _24210_ (.A(_08279_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_2 _24211_ (.A0(_08105_),
    .A1(\fetch.bht.bhtTable_target_pc[5][27] ),
    .S(_06251_),
    .X(_08280_));
 sky130_fd_sc_hd__buf_1 _24212_ (.A(_08280_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_2 _24213_ (.A0(_08107_),
    .A1(\fetch.bht.bhtTable_target_pc[5][28] ),
    .S(_06251_),
    .X(_08281_));
 sky130_fd_sc_hd__buf_1 _24214_ (.A(_08281_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_2 _24215_ (.A0(_08109_),
    .A1(\fetch.bht.bhtTable_target_pc[5][29] ),
    .S(_06251_),
    .X(_08282_));
 sky130_fd_sc_hd__buf_1 _24216_ (.A(_08282_),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_2 _24217_ (.A0(_08111_),
    .A1(\fetch.bht.bhtTable_target_pc[5][30] ),
    .S(_06251_),
    .X(_08283_));
 sky130_fd_sc_hd__buf_1 _24218_ (.A(_08283_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_2 _24219_ (.A0(_08113_),
    .A1(\fetch.bht.bhtTable_target_pc[5][31] ),
    .S(_06251_),
    .X(_08284_));
 sky130_fd_sc_hd__buf_1 _24220_ (.A(_08284_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_2 _24221_ (.A0(_08049_),
    .A1(\fetch.bht.bhtTable_target_pc[6][0] ),
    .S(_06241_),
    .X(_08285_));
 sky130_fd_sc_hd__buf_1 _24222_ (.A(_08285_),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_2 _24223_ (.A0(_08051_),
    .A1(\fetch.bht.bhtTable_target_pc[6][1] ),
    .S(_06241_),
    .X(_08286_));
 sky130_fd_sc_hd__buf_1 _24224_ (.A(_08286_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_2 _24225_ (.A0(_08053_),
    .A1(\fetch.bht.bhtTable_target_pc[6][2] ),
    .S(_06241_),
    .X(_08287_));
 sky130_fd_sc_hd__buf_1 _24226_ (.A(_08287_),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_2 _24227_ (.A0(_08055_),
    .A1(\fetch.bht.bhtTable_target_pc[6][3] ),
    .S(_06241_),
    .X(_08288_));
 sky130_fd_sc_hd__buf_1 _24228_ (.A(_08288_),
    .X(_01786_));
 sky130_fd_sc_hd__buf_1 _24229_ (.A(_06217_),
    .X(_08289_));
 sky130_fd_sc_hd__mux2_2 _24230_ (.A0(_08057_),
    .A1(\fetch.bht.bhtTable_target_pc[6][4] ),
    .S(_08289_),
    .X(_08290_));
 sky130_fd_sc_hd__buf_1 _24231_ (.A(_08290_),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_2 _24232_ (.A0(_08060_),
    .A1(\fetch.bht.bhtTable_target_pc[6][5] ),
    .S(_08289_),
    .X(_08291_));
 sky130_fd_sc_hd__buf_1 _24233_ (.A(_08291_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_2 _24234_ (.A0(_08062_),
    .A1(\fetch.bht.bhtTable_target_pc[6][6] ),
    .S(_08289_),
    .X(_08292_));
 sky130_fd_sc_hd__buf_1 _24235_ (.A(_08292_),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_2 _24236_ (.A0(_08064_),
    .A1(\fetch.bht.bhtTable_target_pc[6][7] ),
    .S(_08289_),
    .X(_08293_));
 sky130_fd_sc_hd__buf_1 _24237_ (.A(_08293_),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_2 _24238_ (.A0(_08066_),
    .A1(\fetch.bht.bhtTable_target_pc[6][8] ),
    .S(_08289_),
    .X(_08294_));
 sky130_fd_sc_hd__buf_1 _24239_ (.A(_08294_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_2 _24240_ (.A0(_08068_),
    .A1(\fetch.bht.bhtTable_target_pc[6][9] ),
    .S(_08289_),
    .X(_08295_));
 sky130_fd_sc_hd__buf_1 _24241_ (.A(_08295_),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_2 _24242_ (.A0(_08070_),
    .A1(\fetch.bht.bhtTable_target_pc[6][10] ),
    .S(_08289_),
    .X(_08296_));
 sky130_fd_sc_hd__buf_1 _24243_ (.A(_08296_),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_2 _24244_ (.A0(_08072_),
    .A1(\fetch.bht.bhtTable_target_pc[6][11] ),
    .S(_08289_),
    .X(_08297_));
 sky130_fd_sc_hd__buf_1 _24245_ (.A(_08297_),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_2 _24246_ (.A0(_08074_),
    .A1(\fetch.bht.bhtTable_target_pc[6][12] ),
    .S(_08289_),
    .X(_08298_));
 sky130_fd_sc_hd__buf_1 _24247_ (.A(_08298_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_2 _24248_ (.A0(_08076_),
    .A1(\fetch.bht.bhtTable_target_pc[6][13] ),
    .S(_08289_),
    .X(_08299_));
 sky130_fd_sc_hd__buf_1 _24249_ (.A(_08299_),
    .X(_01796_));
 sky130_fd_sc_hd__buf_1 _24250_ (.A(_06217_),
    .X(_08300_));
 sky130_fd_sc_hd__mux2_2 _24251_ (.A0(_08078_),
    .A1(\fetch.bht.bhtTable_target_pc[6][14] ),
    .S(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__buf_1 _24252_ (.A(_08301_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_2 _24253_ (.A0(_08081_),
    .A1(\fetch.bht.bhtTable_target_pc[6][15] ),
    .S(_08300_),
    .X(_08302_));
 sky130_fd_sc_hd__buf_1 _24254_ (.A(_08302_),
    .X(_01798_));
 sky130_fd_sc_hd__mux2_2 _24255_ (.A0(_08083_),
    .A1(\fetch.bht.bhtTable_target_pc[6][16] ),
    .S(_08300_),
    .X(_08303_));
 sky130_fd_sc_hd__buf_1 _24256_ (.A(_08303_),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_2 _24257_ (.A0(_08085_),
    .A1(\fetch.bht.bhtTable_target_pc[6][17] ),
    .S(_08300_),
    .X(_08304_));
 sky130_fd_sc_hd__buf_1 _24258_ (.A(_08304_),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_2 _24259_ (.A0(_08087_),
    .A1(\fetch.bht.bhtTable_target_pc[6][18] ),
    .S(_08300_),
    .X(_08305_));
 sky130_fd_sc_hd__buf_1 _24260_ (.A(_08305_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_2 _24261_ (.A0(_08089_),
    .A1(\fetch.bht.bhtTable_target_pc[6][19] ),
    .S(_08300_),
    .X(_08306_));
 sky130_fd_sc_hd__buf_1 _24262_ (.A(_08306_),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_2 _24263_ (.A0(_08091_),
    .A1(\fetch.bht.bhtTable_target_pc[6][20] ),
    .S(_08300_),
    .X(_08307_));
 sky130_fd_sc_hd__buf_1 _24264_ (.A(_08307_),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_2 _24265_ (.A0(_08093_),
    .A1(\fetch.bht.bhtTable_target_pc[6][21] ),
    .S(_08300_),
    .X(_08308_));
 sky130_fd_sc_hd__buf_1 _24266_ (.A(_08308_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_2 _24267_ (.A0(_08095_),
    .A1(\fetch.bht.bhtTable_target_pc[6][22] ),
    .S(_08300_),
    .X(_08309_));
 sky130_fd_sc_hd__buf_1 _24268_ (.A(_08309_),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_2 _24269_ (.A0(_08097_),
    .A1(\fetch.bht.bhtTable_target_pc[6][23] ),
    .S(_08300_),
    .X(_08310_));
 sky130_fd_sc_hd__buf_1 _24270_ (.A(_08310_),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_2 _24271_ (.A0(_08099_),
    .A1(\fetch.bht.bhtTable_target_pc[6][24] ),
    .S(_06218_),
    .X(_08311_));
 sky130_fd_sc_hd__buf_1 _24272_ (.A(_08311_),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_2 _24273_ (.A0(_08101_),
    .A1(\fetch.bht.bhtTable_target_pc[6][25] ),
    .S(_06218_),
    .X(_08312_));
 sky130_fd_sc_hd__buf_1 _24274_ (.A(_08312_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_2 _24275_ (.A0(_08103_),
    .A1(\fetch.bht.bhtTable_target_pc[6][26] ),
    .S(_06218_),
    .X(_08313_));
 sky130_fd_sc_hd__buf_1 _24276_ (.A(_08313_),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_2 _24277_ (.A0(_08105_),
    .A1(\fetch.bht.bhtTable_target_pc[6][27] ),
    .S(_06218_),
    .X(_08314_));
 sky130_fd_sc_hd__buf_1 _24278_ (.A(_08314_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_2 _24279_ (.A0(_08107_),
    .A1(\fetch.bht.bhtTable_target_pc[6][28] ),
    .S(_06218_),
    .X(_08315_));
 sky130_fd_sc_hd__buf_1 _24280_ (.A(_08315_),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_2 _24281_ (.A0(_08109_),
    .A1(\fetch.bht.bhtTable_target_pc[6][29] ),
    .S(_06218_),
    .X(_08316_));
 sky130_fd_sc_hd__buf_1 _24282_ (.A(_08316_),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_2 _24283_ (.A0(_08111_),
    .A1(\fetch.bht.bhtTable_target_pc[6][30] ),
    .S(_06218_),
    .X(_08317_));
 sky130_fd_sc_hd__buf_1 _24284_ (.A(_08317_),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_2 _24285_ (.A0(_08113_),
    .A1(\fetch.bht.bhtTable_target_pc[6][31] ),
    .S(_06218_),
    .X(_08318_));
 sky130_fd_sc_hd__buf_1 _24286_ (.A(_08318_),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_2 _24287_ (.A0(_08049_),
    .A1(\fetch.bht.bhtTable_target_pc[7][0] ),
    .S(_06210_),
    .X(_08319_));
 sky130_fd_sc_hd__buf_1 _24288_ (.A(_08319_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_2 _24289_ (.A0(_08051_),
    .A1(\fetch.bht.bhtTable_target_pc[7][1] ),
    .S(_06210_),
    .X(_08320_));
 sky130_fd_sc_hd__buf_1 _24290_ (.A(_08320_),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_2 _24291_ (.A0(_08053_),
    .A1(\fetch.bht.bhtTable_target_pc[7][2] ),
    .S(_06210_),
    .X(_08321_));
 sky130_fd_sc_hd__buf_1 _24292_ (.A(_08321_),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_2 _24293_ (.A0(_08055_),
    .A1(\fetch.bht.bhtTable_target_pc[7][3] ),
    .S(_06210_),
    .X(_08322_));
 sky130_fd_sc_hd__buf_1 _24294_ (.A(_08322_),
    .X(_01818_));
 sky130_fd_sc_hd__buf_1 _24295_ (.A(_06186_),
    .X(_08323_));
 sky130_fd_sc_hd__mux2_2 _24296_ (.A0(_08057_),
    .A1(\fetch.bht.bhtTable_target_pc[7][4] ),
    .S(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__buf_1 _24297_ (.A(_08324_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_2 _24298_ (.A0(_08060_),
    .A1(\fetch.bht.bhtTable_target_pc[7][5] ),
    .S(_08323_),
    .X(_08325_));
 sky130_fd_sc_hd__buf_1 _24299_ (.A(_08325_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_2 _24300_ (.A0(_08062_),
    .A1(\fetch.bht.bhtTable_target_pc[7][6] ),
    .S(_08323_),
    .X(_08326_));
 sky130_fd_sc_hd__buf_1 _24301_ (.A(_08326_),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_2 _24302_ (.A0(_08064_),
    .A1(\fetch.bht.bhtTable_target_pc[7][7] ),
    .S(_08323_),
    .X(_08327_));
 sky130_fd_sc_hd__buf_1 _24303_ (.A(_08327_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_2 _24304_ (.A0(_08066_),
    .A1(\fetch.bht.bhtTable_target_pc[7][8] ),
    .S(_08323_),
    .X(_08328_));
 sky130_fd_sc_hd__buf_1 _24305_ (.A(_08328_),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_2 _24306_ (.A0(_08068_),
    .A1(\fetch.bht.bhtTable_target_pc[7][9] ),
    .S(_08323_),
    .X(_08329_));
 sky130_fd_sc_hd__buf_1 _24307_ (.A(_08329_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_2 _24308_ (.A0(_08070_),
    .A1(\fetch.bht.bhtTable_target_pc[7][10] ),
    .S(_08323_),
    .X(_08330_));
 sky130_fd_sc_hd__buf_1 _24309_ (.A(_08330_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_2 _24310_ (.A0(_08072_),
    .A1(\fetch.bht.bhtTable_target_pc[7][11] ),
    .S(_08323_),
    .X(_08331_));
 sky130_fd_sc_hd__buf_1 _24311_ (.A(_08331_),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_2 _24312_ (.A0(_08074_),
    .A1(\fetch.bht.bhtTable_target_pc[7][12] ),
    .S(_08323_),
    .X(_08332_));
 sky130_fd_sc_hd__buf_1 _24313_ (.A(_08332_),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_2 _24314_ (.A0(_08076_),
    .A1(\fetch.bht.bhtTable_target_pc[7][13] ),
    .S(_08323_),
    .X(_08333_));
 sky130_fd_sc_hd__buf_1 _24315_ (.A(_08333_),
    .X(_01828_));
 sky130_fd_sc_hd__buf_1 _24316_ (.A(_06186_),
    .X(_08334_));
 sky130_fd_sc_hd__mux2_2 _24317_ (.A0(_08078_),
    .A1(\fetch.bht.bhtTable_target_pc[7][14] ),
    .S(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__buf_1 _24318_ (.A(_08335_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_2 _24319_ (.A0(_08081_),
    .A1(\fetch.bht.bhtTable_target_pc[7][15] ),
    .S(_08334_),
    .X(_08336_));
 sky130_fd_sc_hd__buf_1 _24320_ (.A(_08336_),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_2 _24321_ (.A0(_08083_),
    .A1(\fetch.bht.bhtTable_target_pc[7][16] ),
    .S(_08334_),
    .X(_08337_));
 sky130_fd_sc_hd__buf_1 _24322_ (.A(_08337_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_2 _24323_ (.A0(_08085_),
    .A1(\fetch.bht.bhtTable_target_pc[7][17] ),
    .S(_08334_),
    .X(_08338_));
 sky130_fd_sc_hd__buf_1 _24324_ (.A(_08338_),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_2 _24325_ (.A0(_08087_),
    .A1(\fetch.bht.bhtTable_target_pc[7][18] ),
    .S(_08334_),
    .X(_08339_));
 sky130_fd_sc_hd__buf_1 _24326_ (.A(_08339_),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_2 _24327_ (.A0(_08089_),
    .A1(\fetch.bht.bhtTable_target_pc[7][19] ),
    .S(_08334_),
    .X(_08340_));
 sky130_fd_sc_hd__buf_1 _24328_ (.A(_08340_),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_2 _24329_ (.A0(_08091_),
    .A1(\fetch.bht.bhtTable_target_pc[7][20] ),
    .S(_08334_),
    .X(_08341_));
 sky130_fd_sc_hd__buf_1 _24330_ (.A(_08341_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_2 _24331_ (.A0(_08093_),
    .A1(\fetch.bht.bhtTable_target_pc[7][21] ),
    .S(_08334_),
    .X(_08342_));
 sky130_fd_sc_hd__buf_1 _24332_ (.A(_08342_),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_2 _24333_ (.A0(_08095_),
    .A1(\fetch.bht.bhtTable_target_pc[7][22] ),
    .S(_08334_),
    .X(_08343_));
 sky130_fd_sc_hd__buf_1 _24334_ (.A(_08343_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_2 _24335_ (.A0(_08097_),
    .A1(\fetch.bht.bhtTable_target_pc[7][23] ),
    .S(_08334_),
    .X(_08344_));
 sky130_fd_sc_hd__buf_1 _24336_ (.A(_08344_),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_2 _24337_ (.A0(_08099_),
    .A1(\fetch.bht.bhtTable_target_pc[7][24] ),
    .S(_06187_),
    .X(_08345_));
 sky130_fd_sc_hd__buf_1 _24338_ (.A(_08345_),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_2 _24339_ (.A0(_08101_),
    .A1(\fetch.bht.bhtTable_target_pc[7][25] ),
    .S(_06187_),
    .X(_08346_));
 sky130_fd_sc_hd__buf_1 _24340_ (.A(_08346_),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_2 _24341_ (.A0(_08103_),
    .A1(\fetch.bht.bhtTable_target_pc[7][26] ),
    .S(_06187_),
    .X(_08347_));
 sky130_fd_sc_hd__buf_1 _24342_ (.A(_08347_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_2 _24343_ (.A0(_08105_),
    .A1(\fetch.bht.bhtTable_target_pc[7][27] ),
    .S(_06187_),
    .X(_08348_));
 sky130_fd_sc_hd__buf_1 _24344_ (.A(_08348_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_2 _24345_ (.A0(_08107_),
    .A1(\fetch.bht.bhtTable_target_pc[7][28] ),
    .S(_06187_),
    .X(_08349_));
 sky130_fd_sc_hd__buf_1 _24346_ (.A(_08349_),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_2 _24347_ (.A0(_08109_),
    .A1(\fetch.bht.bhtTable_target_pc[7][29] ),
    .S(_06187_),
    .X(_08350_));
 sky130_fd_sc_hd__buf_1 _24348_ (.A(_08350_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_2 _24349_ (.A0(_08111_),
    .A1(\fetch.bht.bhtTable_target_pc[7][30] ),
    .S(_06187_),
    .X(_08351_));
 sky130_fd_sc_hd__buf_1 _24350_ (.A(_08351_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_2 _24351_ (.A0(_08113_),
    .A1(\fetch.bht.bhtTable_target_pc[7][31] ),
    .S(_06187_),
    .X(_08352_));
 sky130_fd_sc_hd__buf_1 _24352_ (.A(_08352_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_2 _24353_ (.A0(\fetch.bht.bhtTable_target_pc[8][0] ),
    .A1(\execute.io_target_pc[0] ),
    .S(_06141_),
    .X(_08353_));
 sky130_fd_sc_hd__buf_1 _24354_ (.A(_08353_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_2 _24355_ (.A0(\fetch.bht.bhtTable_target_pc[8][1] ),
    .A1(\execute.io_target_pc[1] ),
    .S(_06141_),
    .X(_08354_));
 sky130_fd_sc_hd__buf_1 _24356_ (.A(_08354_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_2 _24357_ (.A0(\fetch.bht.bhtTable_target_pc[8][2] ),
    .A1(\execute.io_target_pc[2] ),
    .S(_06141_),
    .X(_08355_));
 sky130_fd_sc_hd__buf_1 _24358_ (.A(_08355_),
    .X(_01849_));
 sky130_fd_sc_hd__buf_1 _24359_ (.A(_09910_),
    .X(_08356_));
 sky130_fd_sc_hd__mux2_2 _24360_ (.A0(\fetch.bht.bhtTable_target_pc[8][3] ),
    .A1(\execute.io_target_pc[3] ),
    .S(_08356_),
    .X(_08357_));
 sky130_fd_sc_hd__buf_1 _24361_ (.A(_08357_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_2 _24362_ (.A0(\fetch.bht.bhtTable_target_pc[8][4] ),
    .A1(\execute.io_target_pc[4] ),
    .S(_08356_),
    .X(_08358_));
 sky130_fd_sc_hd__buf_1 _24363_ (.A(_08358_),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_2 _24364_ (.A0(\fetch.bht.bhtTable_target_pc[8][5] ),
    .A1(\execute.io_target_pc[5] ),
    .S(_08356_),
    .X(_08359_));
 sky130_fd_sc_hd__buf_1 _24365_ (.A(_08359_),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_2 _24366_ (.A0(\fetch.bht.bhtTable_target_pc[8][6] ),
    .A1(\execute.io_target_pc[6] ),
    .S(_08356_),
    .X(_08360_));
 sky130_fd_sc_hd__buf_1 _24367_ (.A(_08360_),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_2 _24368_ (.A0(\fetch.bht.bhtTable_target_pc[8][7] ),
    .A1(\execute.io_target_pc[7] ),
    .S(_08356_),
    .X(_08361_));
 sky130_fd_sc_hd__buf_1 _24369_ (.A(_08361_),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_2 _24370_ (.A0(\fetch.bht.bhtTable_target_pc[8][8] ),
    .A1(\execute.io_target_pc[8] ),
    .S(_08356_),
    .X(_08362_));
 sky130_fd_sc_hd__buf_1 _24371_ (.A(_08362_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_2 _24372_ (.A0(\fetch.bht.bhtTable_target_pc[8][9] ),
    .A1(\execute.io_target_pc[9] ),
    .S(_08356_),
    .X(_08363_));
 sky130_fd_sc_hd__buf_1 _24373_ (.A(_08363_),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_2 _24374_ (.A0(\fetch.bht.bhtTable_target_pc[8][10] ),
    .A1(\execute.io_target_pc[10] ),
    .S(_08356_),
    .X(_08364_));
 sky130_fd_sc_hd__buf_1 _24375_ (.A(_08364_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_2 _24376_ (.A0(\fetch.bht.bhtTable_target_pc[8][11] ),
    .A1(\execute.io_target_pc[11] ),
    .S(_08356_),
    .X(_08365_));
 sky130_fd_sc_hd__buf_1 _24377_ (.A(_08365_),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_2 _24378_ (.A0(\fetch.bht.bhtTable_target_pc[8][12] ),
    .A1(\execute.io_target_pc[12] ),
    .S(_08356_),
    .X(_08366_));
 sky130_fd_sc_hd__buf_1 _24379_ (.A(_08366_),
    .X(_01859_));
 sky130_fd_sc_hd__buf_1 _24380_ (.A(_09910_),
    .X(_08367_));
 sky130_fd_sc_hd__mux2_2 _24381_ (.A0(\fetch.bht.bhtTable_target_pc[8][13] ),
    .A1(\execute.io_target_pc[13] ),
    .S(_08367_),
    .X(_08368_));
 sky130_fd_sc_hd__buf_1 _24382_ (.A(_08368_),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_2 _24383_ (.A0(\fetch.bht.bhtTable_target_pc[8][14] ),
    .A1(\execute.io_target_pc[14] ),
    .S(_08367_),
    .X(_08369_));
 sky130_fd_sc_hd__buf_1 _24384_ (.A(_08369_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_2 _24385_ (.A0(\fetch.bht.bhtTable_target_pc[8][15] ),
    .A1(\execute.io_target_pc[15] ),
    .S(_08367_),
    .X(_08370_));
 sky130_fd_sc_hd__buf_1 _24386_ (.A(_08370_),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_2 _24387_ (.A0(\fetch.bht.bhtTable_target_pc[8][16] ),
    .A1(\execute.io_target_pc[16] ),
    .S(_08367_),
    .X(_08371_));
 sky130_fd_sc_hd__buf_1 _24388_ (.A(_08371_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_2 _24389_ (.A0(\fetch.bht.bhtTable_target_pc[8][17] ),
    .A1(\execute.io_target_pc[17] ),
    .S(_08367_),
    .X(_08372_));
 sky130_fd_sc_hd__buf_1 _24390_ (.A(_08372_),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_2 _24391_ (.A0(\fetch.bht.bhtTable_target_pc[8][18] ),
    .A1(\execute.io_target_pc[18] ),
    .S(_08367_),
    .X(_08373_));
 sky130_fd_sc_hd__buf_1 _24392_ (.A(_08373_),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_2 _24393_ (.A0(\fetch.bht.bhtTable_target_pc[8][19] ),
    .A1(\execute.io_target_pc[19] ),
    .S(_08367_),
    .X(_08374_));
 sky130_fd_sc_hd__buf_1 _24394_ (.A(_08374_),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_2 _24395_ (.A0(\fetch.bht.bhtTable_target_pc[8][20] ),
    .A1(\execute.io_target_pc[20] ),
    .S(_08367_),
    .X(_08375_));
 sky130_fd_sc_hd__buf_1 _24396_ (.A(_08375_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_2 _24397_ (.A0(\fetch.bht.bhtTable_target_pc[8][21] ),
    .A1(\execute.io_target_pc[21] ),
    .S(_08367_),
    .X(_08376_));
 sky130_fd_sc_hd__buf_1 _24398_ (.A(_08376_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_2 _24399_ (.A0(\fetch.bht.bhtTable_target_pc[8][22] ),
    .A1(\execute.io_target_pc[22] ),
    .S(_08367_),
    .X(_08377_));
 sky130_fd_sc_hd__buf_1 _24400_ (.A(_08377_),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_2 _24401_ (.A0(\fetch.bht.bhtTable_target_pc[8][23] ),
    .A1(\execute.io_target_pc[23] ),
    .S(_09911_),
    .X(_08378_));
 sky130_fd_sc_hd__buf_1 _24402_ (.A(_08378_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_2 _24403_ (.A0(\fetch.bht.bhtTable_target_pc[8][24] ),
    .A1(\execute.io_target_pc[24] ),
    .S(_09911_),
    .X(_08379_));
 sky130_fd_sc_hd__buf_1 _24404_ (.A(_08379_),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_2 _24405_ (.A0(\fetch.bht.bhtTable_target_pc[8][25] ),
    .A1(\execute.io_target_pc[25] ),
    .S(_09911_),
    .X(_08380_));
 sky130_fd_sc_hd__buf_1 _24406_ (.A(_08380_),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_2 _24407_ (.A0(\fetch.bht.bhtTable_target_pc[8][26] ),
    .A1(\execute.io_target_pc[26] ),
    .S(_09911_),
    .X(_08381_));
 sky130_fd_sc_hd__buf_1 _24408_ (.A(_08381_),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_2 _24409_ (.A0(\fetch.bht.bhtTable_target_pc[8][27] ),
    .A1(\execute.io_target_pc[27] ),
    .S(_09911_),
    .X(_08382_));
 sky130_fd_sc_hd__buf_1 _24410_ (.A(_08382_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_2 _24411_ (.A0(\fetch.bht.bhtTable_target_pc[8][28] ),
    .A1(\execute.io_target_pc[28] ),
    .S(_09911_),
    .X(_08383_));
 sky130_fd_sc_hd__buf_1 _24412_ (.A(_08383_),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_2 _24413_ (.A0(\fetch.bht.bhtTable_target_pc[8][29] ),
    .A1(\execute.io_target_pc[29] ),
    .S(_09911_),
    .X(_08384_));
 sky130_fd_sc_hd__buf_1 _24414_ (.A(_08384_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_2 _24415_ (.A0(\fetch.bht.bhtTable_target_pc[8][30] ),
    .A1(\execute.io_target_pc[30] ),
    .S(_09911_),
    .X(_08385_));
 sky130_fd_sc_hd__buf_1 _24416_ (.A(_08385_),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_2 _24417_ (.A0(\fetch.bht.bhtTable_target_pc[8][31] ),
    .A1(\execute.io_target_pc[31] ),
    .S(_09911_),
    .X(_08386_));
 sky130_fd_sc_hd__buf_1 _24418_ (.A(_08386_),
    .X(_01878_));
 sky130_fd_sc_hd__or4b_2 _24419_ (.A(_10556_),
    .B(_10557_),
    .C(_09900_),
    .D_N(_09917_),
    .X(_08387_));
 sky130_fd_sc_hd__buf_1 _24420_ (.A(_08387_),
    .X(_08388_));
 sky130_fd_sc_hd__buf_1 _24421_ (.A(_08388_),
    .X(_08389_));
 sky130_fd_sc_hd__mux2_2 _24422_ (.A0(_08049_),
    .A1(\fetch.bht.bhtTable_target_pc[0][0] ),
    .S(_08389_),
    .X(_08390_));
 sky130_fd_sc_hd__buf_1 _24423_ (.A(_08390_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_2 _24424_ (.A0(_08051_),
    .A1(\fetch.bht.bhtTable_target_pc[0][1] ),
    .S(_08389_),
    .X(_08391_));
 sky130_fd_sc_hd__buf_1 _24425_ (.A(_08391_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_2 _24426_ (.A0(_08053_),
    .A1(\fetch.bht.bhtTable_target_pc[0][2] ),
    .S(_08389_),
    .X(_08392_));
 sky130_fd_sc_hd__buf_1 _24427_ (.A(_08392_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_2 _24428_ (.A0(_08055_),
    .A1(\fetch.bht.bhtTable_target_pc[0][3] ),
    .S(_08389_),
    .X(_08393_));
 sky130_fd_sc_hd__buf_1 _24429_ (.A(_08393_),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_2 _24430_ (.A0(_08057_),
    .A1(\fetch.bht.bhtTable_target_pc[0][4] ),
    .S(_08389_),
    .X(_08394_));
 sky130_fd_sc_hd__buf_1 _24431_ (.A(_08394_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_2 _24432_ (.A0(_08060_),
    .A1(\fetch.bht.bhtTable_target_pc[0][5] ),
    .S(_08389_),
    .X(_08395_));
 sky130_fd_sc_hd__buf_1 _24433_ (.A(_08395_),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_2 _24434_ (.A0(_08062_),
    .A1(\fetch.bht.bhtTable_target_pc[0][6] ),
    .S(_08389_),
    .X(_08396_));
 sky130_fd_sc_hd__buf_1 _24435_ (.A(_08396_),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_2 _24436_ (.A0(_08064_),
    .A1(\fetch.bht.bhtTable_target_pc[0][7] ),
    .S(_08389_),
    .X(_08397_));
 sky130_fd_sc_hd__buf_1 _24437_ (.A(_08397_),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_2 _24438_ (.A0(_08066_),
    .A1(\fetch.bht.bhtTable_target_pc[0][8] ),
    .S(_08389_),
    .X(_08398_));
 sky130_fd_sc_hd__buf_1 _24439_ (.A(_08398_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_2 _24440_ (.A0(_08068_),
    .A1(\fetch.bht.bhtTable_target_pc[0][9] ),
    .S(_08389_),
    .X(_08399_));
 sky130_fd_sc_hd__buf_1 _24441_ (.A(_08399_),
    .X(_01888_));
 sky130_fd_sc_hd__buf_1 _24442_ (.A(_08388_),
    .X(_08400_));
 sky130_fd_sc_hd__mux2_2 _24443_ (.A0(_08070_),
    .A1(\fetch.bht.bhtTable_target_pc[0][10] ),
    .S(_08400_),
    .X(_08401_));
 sky130_fd_sc_hd__buf_1 _24444_ (.A(_08401_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_2 _24445_ (.A0(_08072_),
    .A1(\fetch.bht.bhtTable_target_pc[0][11] ),
    .S(_08400_),
    .X(_08402_));
 sky130_fd_sc_hd__buf_1 _24446_ (.A(_08402_),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_2 _24447_ (.A0(_08074_),
    .A1(\fetch.bht.bhtTable_target_pc[0][12] ),
    .S(_08400_),
    .X(_08403_));
 sky130_fd_sc_hd__buf_1 _24448_ (.A(_08403_),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_2 _24449_ (.A0(_08076_),
    .A1(\fetch.bht.bhtTable_target_pc[0][13] ),
    .S(_08400_),
    .X(_08404_));
 sky130_fd_sc_hd__buf_1 _24450_ (.A(_08404_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_2 _24451_ (.A0(_08078_),
    .A1(\fetch.bht.bhtTable_target_pc[0][14] ),
    .S(_08400_),
    .X(_08405_));
 sky130_fd_sc_hd__buf_1 _24452_ (.A(_08405_),
    .X(_01893_));
 sky130_fd_sc_hd__mux2_2 _24453_ (.A0(_08081_),
    .A1(\fetch.bht.bhtTable_target_pc[0][15] ),
    .S(_08400_),
    .X(_08406_));
 sky130_fd_sc_hd__buf_1 _24454_ (.A(_08406_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_2 _24455_ (.A0(_08083_),
    .A1(\fetch.bht.bhtTable_target_pc[0][16] ),
    .S(_08400_),
    .X(_08407_));
 sky130_fd_sc_hd__buf_1 _24456_ (.A(_08407_),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_2 _24457_ (.A0(_08085_),
    .A1(\fetch.bht.bhtTable_target_pc[0][17] ),
    .S(_08400_),
    .X(_08408_));
 sky130_fd_sc_hd__buf_1 _24458_ (.A(_08408_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_2 _24459_ (.A0(_08087_),
    .A1(\fetch.bht.bhtTable_target_pc[0][18] ),
    .S(_08400_),
    .X(_08409_));
 sky130_fd_sc_hd__buf_1 _24460_ (.A(_08409_),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_2 _24461_ (.A0(_08089_),
    .A1(\fetch.bht.bhtTable_target_pc[0][19] ),
    .S(_08400_),
    .X(_08410_));
 sky130_fd_sc_hd__buf_1 _24462_ (.A(_08410_),
    .X(_01898_));
 sky130_fd_sc_hd__buf_1 _24463_ (.A(_08387_),
    .X(_08411_));
 sky130_fd_sc_hd__mux2_2 _24464_ (.A0(_08091_),
    .A1(\fetch.bht.bhtTable_target_pc[0][20] ),
    .S(_08411_),
    .X(_08412_));
 sky130_fd_sc_hd__buf_1 _24465_ (.A(_08412_),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_2 _24466_ (.A0(_08093_),
    .A1(\fetch.bht.bhtTable_target_pc[0][21] ),
    .S(_08411_),
    .X(_08413_));
 sky130_fd_sc_hd__buf_1 _24467_ (.A(_08413_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_2 _24468_ (.A0(_08095_),
    .A1(\fetch.bht.bhtTable_target_pc[0][22] ),
    .S(_08411_),
    .X(_08414_));
 sky130_fd_sc_hd__buf_1 _24469_ (.A(_08414_),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_2 _24470_ (.A0(_08097_),
    .A1(\fetch.bht.bhtTable_target_pc[0][23] ),
    .S(_08411_),
    .X(_08415_));
 sky130_fd_sc_hd__buf_1 _24471_ (.A(_08415_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_2 _24472_ (.A0(_08099_),
    .A1(\fetch.bht.bhtTable_target_pc[0][24] ),
    .S(_08411_),
    .X(_08416_));
 sky130_fd_sc_hd__buf_1 _24473_ (.A(_08416_),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_2 _24474_ (.A0(_08101_),
    .A1(\fetch.bht.bhtTable_target_pc[0][25] ),
    .S(_08411_),
    .X(_08417_));
 sky130_fd_sc_hd__buf_1 _24475_ (.A(_08417_),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_2 _24476_ (.A0(_08103_),
    .A1(\fetch.bht.bhtTable_target_pc[0][26] ),
    .S(_08411_),
    .X(_08418_));
 sky130_fd_sc_hd__buf_1 _24477_ (.A(_08418_),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_2 _24478_ (.A0(_08105_),
    .A1(\fetch.bht.bhtTable_target_pc[0][27] ),
    .S(_08411_),
    .X(_08419_));
 sky130_fd_sc_hd__buf_1 _24479_ (.A(_08419_),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_2 _24480_ (.A0(_08107_),
    .A1(\fetch.bht.bhtTable_target_pc[0][28] ),
    .S(_08411_),
    .X(_08420_));
 sky130_fd_sc_hd__buf_1 _24481_ (.A(_08420_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_2 _24482_ (.A0(_08109_),
    .A1(\fetch.bht.bhtTable_target_pc[0][29] ),
    .S(_08411_),
    .X(_08421_));
 sky130_fd_sc_hd__buf_1 _24483_ (.A(_08421_),
    .X(_01908_));
 sky130_fd_sc_hd__buf_1 _24484_ (.A(_08387_),
    .X(_08422_));
 sky130_fd_sc_hd__mux2_2 _24485_ (.A0(_08111_),
    .A1(\fetch.bht.bhtTable_target_pc[0][30] ),
    .S(_08422_),
    .X(_08423_));
 sky130_fd_sc_hd__buf_1 _24486_ (.A(_08423_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_2 _24487_ (.A0(_08113_),
    .A1(\fetch.bht.bhtTable_target_pc[0][31] ),
    .S(_08422_),
    .X(_08424_));
 sky130_fd_sc_hd__buf_1 _24488_ (.A(_08424_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_2 _24489_ (.A0(_08049_),
    .A1(\fetch.bht.bhtTable_target_pc[10][0] ),
    .S(_07276_),
    .X(_08425_));
 sky130_fd_sc_hd__buf_1 _24490_ (.A(_08425_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_2 _24491_ (.A0(_08051_),
    .A1(\fetch.bht.bhtTable_target_pc[10][1] ),
    .S(_07276_),
    .X(_08426_));
 sky130_fd_sc_hd__buf_1 _24492_ (.A(_08426_),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_2 _24493_ (.A0(_08053_),
    .A1(\fetch.bht.bhtTable_target_pc[10][2] ),
    .S(_07276_),
    .X(_08427_));
 sky130_fd_sc_hd__buf_1 _24494_ (.A(_08427_),
    .X(_01913_));
 sky130_fd_sc_hd__buf_1 _24495_ (.A(_09901_),
    .X(_08428_));
 sky130_fd_sc_hd__mux2_2 _24496_ (.A0(_08055_),
    .A1(\fetch.bht.bhtTable_target_pc[10][3] ),
    .S(_08428_),
    .X(_08429_));
 sky130_fd_sc_hd__buf_1 _24497_ (.A(_08429_),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_2 _24498_ (.A0(_08057_),
    .A1(\fetch.bht.bhtTable_target_pc[10][4] ),
    .S(_08428_),
    .X(_08430_));
 sky130_fd_sc_hd__buf_1 _24499_ (.A(_08430_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_2 _24500_ (.A0(_08060_),
    .A1(\fetch.bht.bhtTable_target_pc[10][5] ),
    .S(_08428_),
    .X(_08431_));
 sky130_fd_sc_hd__buf_1 _24501_ (.A(_08431_),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_2 _24502_ (.A0(_08062_),
    .A1(\fetch.bht.bhtTable_target_pc[10][6] ),
    .S(_08428_),
    .X(_08432_));
 sky130_fd_sc_hd__buf_1 _24503_ (.A(_08432_),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_2 _24504_ (.A0(_08064_),
    .A1(\fetch.bht.bhtTable_target_pc[10][7] ),
    .S(_08428_),
    .X(_08433_));
 sky130_fd_sc_hd__buf_1 _24505_ (.A(_08433_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_2 _24506_ (.A0(_08066_),
    .A1(\fetch.bht.bhtTable_target_pc[10][8] ),
    .S(_08428_),
    .X(_08434_));
 sky130_fd_sc_hd__buf_1 _24507_ (.A(_08434_),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_2 _24508_ (.A0(_08068_),
    .A1(\fetch.bht.bhtTable_target_pc[10][9] ),
    .S(_08428_),
    .X(_08435_));
 sky130_fd_sc_hd__buf_1 _24509_ (.A(_08435_),
    .X(_01920_));
 sky130_fd_sc_hd__mux2_2 _24510_ (.A0(_08070_),
    .A1(\fetch.bht.bhtTable_target_pc[10][10] ),
    .S(_08428_),
    .X(_08436_));
 sky130_fd_sc_hd__buf_1 _24511_ (.A(_08436_),
    .X(_01921_));
 sky130_fd_sc_hd__mux2_2 _24512_ (.A0(_08072_),
    .A1(\fetch.bht.bhtTable_target_pc[10][11] ),
    .S(_08428_),
    .X(_08437_));
 sky130_fd_sc_hd__buf_1 _24513_ (.A(_08437_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_2 _24514_ (.A0(_08074_),
    .A1(\fetch.bht.bhtTable_target_pc[10][12] ),
    .S(_08428_),
    .X(_08438_));
 sky130_fd_sc_hd__buf_1 _24515_ (.A(_08438_),
    .X(_01923_));
 sky130_fd_sc_hd__buf_1 _24516_ (.A(_09901_),
    .X(_08439_));
 sky130_fd_sc_hd__mux2_2 _24517_ (.A0(_08076_),
    .A1(\fetch.bht.bhtTable_target_pc[10][13] ),
    .S(_08439_),
    .X(_08440_));
 sky130_fd_sc_hd__buf_1 _24518_ (.A(_08440_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_2 _24519_ (.A0(_08078_),
    .A1(\fetch.bht.bhtTable_target_pc[10][14] ),
    .S(_08439_),
    .X(_08441_));
 sky130_fd_sc_hd__buf_1 _24520_ (.A(_08441_),
    .X(_01925_));
 sky130_fd_sc_hd__mux2_2 _24521_ (.A0(_08081_),
    .A1(\fetch.bht.bhtTable_target_pc[10][15] ),
    .S(_08439_),
    .X(_08442_));
 sky130_fd_sc_hd__buf_1 _24522_ (.A(_08442_),
    .X(_01926_));
 sky130_fd_sc_hd__mux2_2 _24523_ (.A0(_08083_),
    .A1(\fetch.bht.bhtTable_target_pc[10][16] ),
    .S(_08439_),
    .X(_08443_));
 sky130_fd_sc_hd__buf_1 _24524_ (.A(_08443_),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_2 _24525_ (.A0(_08085_),
    .A1(\fetch.bht.bhtTable_target_pc[10][17] ),
    .S(_08439_),
    .X(_08444_));
 sky130_fd_sc_hd__buf_1 _24526_ (.A(_08444_),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_2 _24527_ (.A0(_08087_),
    .A1(\fetch.bht.bhtTable_target_pc[10][18] ),
    .S(_08439_),
    .X(_08445_));
 sky130_fd_sc_hd__buf_1 _24528_ (.A(_08445_),
    .X(_01929_));
 sky130_fd_sc_hd__mux2_2 _24529_ (.A0(_08089_),
    .A1(\fetch.bht.bhtTable_target_pc[10][19] ),
    .S(_08439_),
    .X(_08446_));
 sky130_fd_sc_hd__buf_1 _24530_ (.A(_08446_),
    .X(_01930_));
 sky130_fd_sc_hd__mux2_2 _24531_ (.A0(_08091_),
    .A1(\fetch.bht.bhtTable_target_pc[10][20] ),
    .S(_08439_),
    .X(_08447_));
 sky130_fd_sc_hd__buf_1 _24532_ (.A(_08447_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_2 _24533_ (.A0(_08093_),
    .A1(\fetch.bht.bhtTable_target_pc[10][21] ),
    .S(_08439_),
    .X(_08448_));
 sky130_fd_sc_hd__buf_1 _24534_ (.A(_08448_),
    .X(_01932_));
 sky130_fd_sc_hd__mux2_2 _24535_ (.A0(_08095_),
    .A1(\fetch.bht.bhtTable_target_pc[10][22] ),
    .S(_08439_),
    .X(_08449_));
 sky130_fd_sc_hd__buf_1 _24536_ (.A(_08449_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_2 _24537_ (.A0(_08097_),
    .A1(\fetch.bht.bhtTable_target_pc[10][23] ),
    .S(_09902_),
    .X(_08450_));
 sky130_fd_sc_hd__buf_1 _24538_ (.A(_08450_),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_2 _24539_ (.A0(_08099_),
    .A1(\fetch.bht.bhtTable_target_pc[10][24] ),
    .S(_09902_),
    .X(_08451_));
 sky130_fd_sc_hd__buf_1 _24540_ (.A(_08451_),
    .X(_01935_));
 sky130_fd_sc_hd__mux2_2 _24541_ (.A0(_08101_),
    .A1(\fetch.bht.bhtTable_target_pc[10][25] ),
    .S(_09902_),
    .X(_08452_));
 sky130_fd_sc_hd__buf_1 _24542_ (.A(_08452_),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_2 _24543_ (.A0(_08103_),
    .A1(\fetch.bht.bhtTable_target_pc[10][26] ),
    .S(_09902_),
    .X(_08453_));
 sky130_fd_sc_hd__buf_1 _24544_ (.A(_08453_),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_2 _24545_ (.A0(_08105_),
    .A1(\fetch.bht.bhtTable_target_pc[10][27] ),
    .S(_09902_),
    .X(_08454_));
 sky130_fd_sc_hd__buf_1 _24546_ (.A(_08454_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_2 _24547_ (.A0(_08107_),
    .A1(\fetch.bht.bhtTable_target_pc[10][28] ),
    .S(_09902_),
    .X(_08455_));
 sky130_fd_sc_hd__buf_1 _24548_ (.A(_08455_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_2 _24549_ (.A0(_08109_),
    .A1(\fetch.bht.bhtTable_target_pc[10][29] ),
    .S(_09902_),
    .X(_08456_));
 sky130_fd_sc_hd__buf_1 _24550_ (.A(_08456_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_2 _24551_ (.A0(_08111_),
    .A1(\fetch.bht.bhtTable_target_pc[10][30] ),
    .S(_09902_),
    .X(_08457_));
 sky130_fd_sc_hd__buf_1 _24552_ (.A(_08457_),
    .X(_01941_));
 sky130_fd_sc_hd__mux2_2 _24553_ (.A0(_08113_),
    .A1(\fetch.bht.bhtTable_target_pc[10][31] ),
    .S(_09902_),
    .X(_08458_));
 sky130_fd_sc_hd__buf_1 _24554_ (.A(_08458_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_2 _24555_ (.A0(\fetch.bht.bhtTable_target_pc[11][0] ),
    .A1(\execute.io_target_pc[0] ),
    .S(_07335_),
    .X(_08459_));
 sky130_fd_sc_hd__buf_1 _24556_ (.A(_08459_),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_2 _24557_ (.A0(\fetch.bht.bhtTable_target_pc[11][1] ),
    .A1(\execute.io_target_pc[1] ),
    .S(_07335_),
    .X(_08460_));
 sky130_fd_sc_hd__buf_1 _24558_ (.A(_08460_),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_2 _24559_ (.A0(\fetch.bht.bhtTable_target_pc[11][2] ),
    .A1(\execute.io_target_pc[2] ),
    .S(_07335_),
    .X(_08461_));
 sky130_fd_sc_hd__buf_1 _24560_ (.A(_08461_),
    .X(_01945_));
 sky130_fd_sc_hd__buf_1 _24561_ (.A(_09896_),
    .X(_08462_));
 sky130_fd_sc_hd__mux2_2 _24562_ (.A0(\fetch.bht.bhtTable_target_pc[11][3] ),
    .A1(\execute.io_target_pc[3] ),
    .S(_08462_),
    .X(_08463_));
 sky130_fd_sc_hd__buf_1 _24563_ (.A(_08463_),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_2 _24564_ (.A0(\fetch.bht.bhtTable_target_pc[11][4] ),
    .A1(\execute.io_target_pc[4] ),
    .S(_08462_),
    .X(_08464_));
 sky130_fd_sc_hd__buf_1 _24565_ (.A(_08464_),
    .X(_01947_));
 sky130_fd_sc_hd__mux2_2 _24566_ (.A0(\fetch.bht.bhtTable_target_pc[11][5] ),
    .A1(\execute.io_target_pc[5] ),
    .S(_08462_),
    .X(_08465_));
 sky130_fd_sc_hd__buf_1 _24567_ (.A(_08465_),
    .X(_01948_));
 sky130_fd_sc_hd__mux2_2 _24568_ (.A0(\fetch.bht.bhtTable_target_pc[11][6] ),
    .A1(\execute.io_target_pc[6] ),
    .S(_08462_),
    .X(_08466_));
 sky130_fd_sc_hd__buf_1 _24569_ (.A(_08466_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_2 _24570_ (.A0(\fetch.bht.bhtTable_target_pc[11][7] ),
    .A1(\execute.io_target_pc[7] ),
    .S(_08462_),
    .X(_08467_));
 sky130_fd_sc_hd__buf_1 _24571_ (.A(_08467_),
    .X(_01950_));
 sky130_fd_sc_hd__mux2_2 _24572_ (.A0(\fetch.bht.bhtTable_target_pc[11][8] ),
    .A1(\execute.io_target_pc[8] ),
    .S(_08462_),
    .X(_08468_));
 sky130_fd_sc_hd__buf_1 _24573_ (.A(_08468_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_2 _24574_ (.A0(\fetch.bht.bhtTable_target_pc[11][9] ),
    .A1(\execute.io_target_pc[9] ),
    .S(_08462_),
    .X(_08469_));
 sky130_fd_sc_hd__buf_1 _24575_ (.A(_08469_),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_2 _24576_ (.A0(\fetch.bht.bhtTable_target_pc[11][10] ),
    .A1(\execute.io_target_pc[10] ),
    .S(_08462_),
    .X(_08470_));
 sky130_fd_sc_hd__buf_1 _24577_ (.A(_08470_),
    .X(_01953_));
 sky130_fd_sc_hd__mux2_2 _24578_ (.A0(\fetch.bht.bhtTable_target_pc[11][11] ),
    .A1(\execute.io_target_pc[11] ),
    .S(_08462_),
    .X(_08471_));
 sky130_fd_sc_hd__buf_1 _24579_ (.A(_08471_),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_2 _24580_ (.A0(\fetch.bht.bhtTable_target_pc[11][12] ),
    .A1(\execute.io_target_pc[12] ),
    .S(_08462_),
    .X(_08472_));
 sky130_fd_sc_hd__buf_1 _24581_ (.A(_08472_),
    .X(_01955_));
 sky130_fd_sc_hd__buf_1 _24582_ (.A(_09896_),
    .X(_08473_));
 sky130_fd_sc_hd__mux2_2 _24583_ (.A0(\fetch.bht.bhtTable_target_pc[11][13] ),
    .A1(\execute.io_target_pc[13] ),
    .S(_08473_),
    .X(_08474_));
 sky130_fd_sc_hd__buf_1 _24584_ (.A(_08474_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_2 _24585_ (.A0(\fetch.bht.bhtTable_target_pc[11][14] ),
    .A1(\execute.io_target_pc[14] ),
    .S(_08473_),
    .X(_08475_));
 sky130_fd_sc_hd__buf_1 _24586_ (.A(_08475_),
    .X(_01957_));
 sky130_fd_sc_hd__mux2_2 _24587_ (.A0(\fetch.bht.bhtTable_target_pc[11][15] ),
    .A1(\execute.io_target_pc[15] ),
    .S(_08473_),
    .X(_08476_));
 sky130_fd_sc_hd__buf_1 _24588_ (.A(_08476_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_2 _24589_ (.A0(\fetch.bht.bhtTable_target_pc[11][16] ),
    .A1(\execute.io_target_pc[16] ),
    .S(_08473_),
    .X(_08477_));
 sky130_fd_sc_hd__buf_1 _24590_ (.A(_08477_),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_2 _24591_ (.A0(\fetch.bht.bhtTable_target_pc[11][17] ),
    .A1(\execute.io_target_pc[17] ),
    .S(_08473_),
    .X(_08478_));
 sky130_fd_sc_hd__buf_1 _24592_ (.A(_08478_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_2 _24593_ (.A0(\fetch.bht.bhtTable_target_pc[11][18] ),
    .A1(\execute.io_target_pc[18] ),
    .S(_08473_),
    .X(_08479_));
 sky130_fd_sc_hd__buf_1 _24594_ (.A(_08479_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_2 _24595_ (.A0(\fetch.bht.bhtTable_target_pc[11][19] ),
    .A1(\execute.io_target_pc[19] ),
    .S(_08473_),
    .X(_08480_));
 sky130_fd_sc_hd__buf_1 _24596_ (.A(_08480_),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_2 _24597_ (.A0(\fetch.bht.bhtTable_target_pc[11][20] ),
    .A1(\execute.io_target_pc[20] ),
    .S(_08473_),
    .X(_08481_));
 sky130_fd_sc_hd__buf_1 _24598_ (.A(_08481_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_2 _24599_ (.A0(\fetch.bht.bhtTable_target_pc[11][21] ),
    .A1(\execute.io_target_pc[21] ),
    .S(_08473_),
    .X(_08482_));
 sky130_fd_sc_hd__buf_1 _24600_ (.A(_08482_),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_2 _24601_ (.A0(\fetch.bht.bhtTable_target_pc[11][22] ),
    .A1(\execute.io_target_pc[22] ),
    .S(_08473_),
    .X(_08483_));
 sky130_fd_sc_hd__buf_1 _24602_ (.A(_08483_),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_2 _24603_ (.A0(\fetch.bht.bhtTable_target_pc[11][23] ),
    .A1(\execute.io_target_pc[23] ),
    .S(_09897_),
    .X(_08484_));
 sky130_fd_sc_hd__buf_1 _24604_ (.A(_08484_),
    .X(_01966_));
 sky130_fd_sc_hd__mux2_2 _24605_ (.A0(\fetch.bht.bhtTable_target_pc[11][24] ),
    .A1(\execute.io_target_pc[24] ),
    .S(_09897_),
    .X(_08485_));
 sky130_fd_sc_hd__buf_1 _24606_ (.A(_08485_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_2 _24607_ (.A0(\fetch.bht.bhtTable_target_pc[11][25] ),
    .A1(\execute.io_target_pc[25] ),
    .S(_09897_),
    .X(_08486_));
 sky130_fd_sc_hd__buf_1 _24608_ (.A(_08486_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_2 _24609_ (.A0(\fetch.bht.bhtTable_target_pc[11][26] ),
    .A1(\execute.io_target_pc[26] ),
    .S(_09897_),
    .X(_08487_));
 sky130_fd_sc_hd__buf_1 _24610_ (.A(_08487_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_2 _24611_ (.A0(\fetch.bht.bhtTable_target_pc[11][27] ),
    .A1(\execute.io_target_pc[27] ),
    .S(_09897_),
    .X(_08488_));
 sky130_fd_sc_hd__buf_1 _24612_ (.A(_08488_),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_2 _24613_ (.A0(\fetch.bht.bhtTable_target_pc[11][28] ),
    .A1(\execute.io_target_pc[28] ),
    .S(_09897_),
    .X(_08489_));
 sky130_fd_sc_hd__buf_1 _24614_ (.A(_08489_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_2 _24615_ (.A0(\fetch.bht.bhtTable_target_pc[11][29] ),
    .A1(\execute.io_target_pc[29] ),
    .S(_09897_),
    .X(_08490_));
 sky130_fd_sc_hd__buf_1 _24616_ (.A(_08490_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_2 _24617_ (.A0(\fetch.bht.bhtTable_target_pc[11][30] ),
    .A1(\execute.io_target_pc[30] ),
    .S(_09897_),
    .X(_08491_));
 sky130_fd_sc_hd__buf_1 _24618_ (.A(_08491_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_2 _24619_ (.A0(\fetch.bht.bhtTable_target_pc[11][31] ),
    .A1(\execute.io_target_pc[31] ),
    .S(_09897_),
    .X(_08492_));
 sky130_fd_sc_hd__buf_1 _24620_ (.A(_08492_),
    .X(_01974_));
 sky130_fd_sc_hd__mux2_2 _24621_ (.A0(\fetch.bht.bhtTable_target_pc[12][0] ),
    .A1(\execute.io_target_pc[0] ),
    .S(_07308_),
    .X(_08493_));
 sky130_fd_sc_hd__buf_1 _24622_ (.A(_08493_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_2 _24623_ (.A0(\fetch.bht.bhtTable_target_pc[12][1] ),
    .A1(\execute.io_target_pc[1] ),
    .S(_07308_),
    .X(_08494_));
 sky130_fd_sc_hd__buf_1 _24624_ (.A(_08494_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_2 _24625_ (.A0(\fetch.bht.bhtTable_target_pc[12][2] ),
    .A1(\execute.io_target_pc[2] ),
    .S(_07308_),
    .X(_08495_));
 sky130_fd_sc_hd__buf_1 _24626_ (.A(_08495_),
    .X(_01977_));
 sky130_fd_sc_hd__mux2_2 _24627_ (.A0(\fetch.bht.bhtTable_target_pc[12][3] ),
    .A1(\execute.io_target_pc[3] ),
    .S(_07308_),
    .X(_08496_));
 sky130_fd_sc_hd__buf_1 _24628_ (.A(_08496_),
    .X(_01978_));
 sky130_fd_sc_hd__buf_1 _24629_ (.A(_07284_),
    .X(_08497_));
 sky130_fd_sc_hd__mux2_2 _24630_ (.A0(\fetch.bht.bhtTable_target_pc[12][4] ),
    .A1(\execute.io_target_pc[4] ),
    .S(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__buf_1 _24631_ (.A(_08498_),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_2 _24632_ (.A0(\fetch.bht.bhtTable_target_pc[12][5] ),
    .A1(\execute.io_target_pc[5] ),
    .S(_08497_),
    .X(_08499_));
 sky130_fd_sc_hd__buf_1 _24633_ (.A(_08499_),
    .X(_01980_));
 sky130_fd_sc_hd__mux2_2 _24634_ (.A0(\fetch.bht.bhtTable_target_pc[12][6] ),
    .A1(\execute.io_target_pc[6] ),
    .S(_08497_),
    .X(_08500_));
 sky130_fd_sc_hd__buf_1 _24635_ (.A(_08500_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_2 _24636_ (.A0(\fetch.bht.bhtTable_target_pc[12][7] ),
    .A1(\execute.io_target_pc[7] ),
    .S(_08497_),
    .X(_08501_));
 sky130_fd_sc_hd__buf_1 _24637_ (.A(_08501_),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_2 _24638_ (.A0(\fetch.bht.bhtTable_target_pc[12][8] ),
    .A1(\execute.io_target_pc[8] ),
    .S(_08497_),
    .X(_08502_));
 sky130_fd_sc_hd__buf_1 _24639_ (.A(_08502_),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_2 _24640_ (.A0(\fetch.bht.bhtTable_target_pc[12][9] ),
    .A1(\execute.io_target_pc[9] ),
    .S(_08497_),
    .X(_08503_));
 sky130_fd_sc_hd__buf_1 _24641_ (.A(_08503_),
    .X(_01984_));
 sky130_fd_sc_hd__mux2_2 _24642_ (.A0(\fetch.bht.bhtTable_target_pc[12][10] ),
    .A1(\execute.io_target_pc[10] ),
    .S(_08497_),
    .X(_08504_));
 sky130_fd_sc_hd__buf_1 _24643_ (.A(_08504_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_2 _24644_ (.A0(\fetch.bht.bhtTable_target_pc[12][11] ),
    .A1(\execute.io_target_pc[11] ),
    .S(_08497_),
    .X(_08505_));
 sky130_fd_sc_hd__buf_1 _24645_ (.A(_08505_),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_2 _24646_ (.A0(\fetch.bht.bhtTable_target_pc[12][12] ),
    .A1(\execute.io_target_pc[12] ),
    .S(_08497_),
    .X(_08506_));
 sky130_fd_sc_hd__buf_1 _24647_ (.A(_08506_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_2 _24648_ (.A0(\fetch.bht.bhtTable_target_pc[12][13] ),
    .A1(\execute.io_target_pc[13] ),
    .S(_08497_),
    .X(_08507_));
 sky130_fd_sc_hd__buf_1 _24649_ (.A(_08507_),
    .X(_01988_));
 sky130_fd_sc_hd__buf_1 _24650_ (.A(_07284_),
    .X(_08508_));
 sky130_fd_sc_hd__mux2_2 _24651_ (.A0(\fetch.bht.bhtTable_target_pc[12][14] ),
    .A1(\execute.io_target_pc[14] ),
    .S(_08508_),
    .X(_08509_));
 sky130_fd_sc_hd__buf_1 _24652_ (.A(_08509_),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_2 _24653_ (.A0(\fetch.bht.bhtTable_target_pc[12][15] ),
    .A1(\execute.io_target_pc[15] ),
    .S(_08508_),
    .X(_08510_));
 sky130_fd_sc_hd__buf_1 _24654_ (.A(_08510_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_2 _24655_ (.A0(\fetch.bht.bhtTable_target_pc[12][16] ),
    .A1(\execute.io_target_pc[16] ),
    .S(_08508_),
    .X(_08511_));
 sky130_fd_sc_hd__buf_1 _24656_ (.A(_08511_),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_2 _24657_ (.A0(\fetch.bht.bhtTable_target_pc[12][17] ),
    .A1(\execute.io_target_pc[17] ),
    .S(_08508_),
    .X(_08512_));
 sky130_fd_sc_hd__buf_1 _24658_ (.A(_08512_),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_2 _24659_ (.A0(\fetch.bht.bhtTable_target_pc[12][18] ),
    .A1(\execute.io_target_pc[18] ),
    .S(_08508_),
    .X(_08513_));
 sky130_fd_sc_hd__buf_1 _24660_ (.A(_08513_),
    .X(_01993_));
 sky130_fd_sc_hd__mux2_2 _24661_ (.A0(\fetch.bht.bhtTable_target_pc[12][19] ),
    .A1(\execute.io_target_pc[19] ),
    .S(_08508_),
    .X(_08514_));
 sky130_fd_sc_hd__buf_1 _24662_ (.A(_08514_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_2 _24663_ (.A0(\fetch.bht.bhtTable_target_pc[12][20] ),
    .A1(\execute.io_target_pc[20] ),
    .S(_08508_),
    .X(_08515_));
 sky130_fd_sc_hd__buf_1 _24664_ (.A(_08515_),
    .X(_01995_));
 sky130_fd_sc_hd__mux2_2 _24665_ (.A0(\fetch.bht.bhtTable_target_pc[12][21] ),
    .A1(\execute.io_target_pc[21] ),
    .S(_08508_),
    .X(_08516_));
 sky130_fd_sc_hd__buf_1 _24666_ (.A(_08516_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_2 _24667_ (.A0(\fetch.bht.bhtTable_target_pc[12][22] ),
    .A1(\execute.io_target_pc[22] ),
    .S(_08508_),
    .X(_08517_));
 sky130_fd_sc_hd__buf_1 _24668_ (.A(_08517_),
    .X(_01997_));
 sky130_fd_sc_hd__mux2_2 _24669_ (.A0(\fetch.bht.bhtTable_target_pc[12][23] ),
    .A1(\execute.io_target_pc[23] ),
    .S(_08508_),
    .X(_08518_));
 sky130_fd_sc_hd__buf_1 _24670_ (.A(_08518_),
    .X(_01998_));
 sky130_fd_sc_hd__mux2_2 _24671_ (.A0(\fetch.bht.bhtTable_target_pc[12][24] ),
    .A1(\execute.io_target_pc[24] ),
    .S(_07285_),
    .X(_08519_));
 sky130_fd_sc_hd__buf_1 _24672_ (.A(_08519_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_2 _24673_ (.A0(\fetch.bht.bhtTable_target_pc[12][25] ),
    .A1(\execute.io_target_pc[25] ),
    .S(_07285_),
    .X(_08520_));
 sky130_fd_sc_hd__buf_1 _24674_ (.A(_08520_),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_2 _24675_ (.A0(\fetch.bht.bhtTable_target_pc[12][26] ),
    .A1(\execute.io_target_pc[26] ),
    .S(_07285_),
    .X(_08521_));
 sky130_fd_sc_hd__buf_1 _24676_ (.A(_08521_),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_2 _24677_ (.A0(\fetch.bht.bhtTable_target_pc[12][27] ),
    .A1(\execute.io_target_pc[27] ),
    .S(_07285_),
    .X(_08522_));
 sky130_fd_sc_hd__buf_1 _24678_ (.A(_08522_),
    .X(_02002_));
 sky130_fd_sc_hd__mux2_2 _24679_ (.A0(\fetch.bht.bhtTable_target_pc[12][28] ),
    .A1(\execute.io_target_pc[28] ),
    .S(_07285_),
    .X(_08523_));
 sky130_fd_sc_hd__buf_1 _24680_ (.A(_08523_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_2 _24681_ (.A0(\fetch.bht.bhtTable_target_pc[12][29] ),
    .A1(\execute.io_target_pc[29] ),
    .S(_07285_),
    .X(_08524_));
 sky130_fd_sc_hd__buf_1 _24682_ (.A(_08524_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_2 _24683_ (.A0(\fetch.bht.bhtTable_target_pc[12][30] ),
    .A1(\execute.io_target_pc[30] ),
    .S(_07285_),
    .X(_08525_));
 sky130_fd_sc_hd__buf_1 _24684_ (.A(_08525_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_2 _24685_ (.A0(\fetch.bht.bhtTable_target_pc[12][31] ),
    .A1(\execute.io_target_pc[31] ),
    .S(_07285_),
    .X(_08526_));
 sky130_fd_sc_hd__buf_1 _24686_ (.A(_08526_),
    .X(_02006_));
 sky130_fd_sc_hd__mux2_2 _24687_ (.A0(_08049_),
    .A1(\fetch.bht.bhtTable_target_pc[13][0] ),
    .S(_06306_),
    .X(_08527_));
 sky130_fd_sc_hd__buf_1 _24688_ (.A(_08527_),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_2 _24689_ (.A0(_08051_),
    .A1(\fetch.bht.bhtTable_target_pc[13][1] ),
    .S(_06306_),
    .X(_08528_));
 sky130_fd_sc_hd__buf_1 _24690_ (.A(_08528_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_2 _24691_ (.A0(_08053_),
    .A1(\fetch.bht.bhtTable_target_pc[13][2] ),
    .S(_06306_),
    .X(_08529_));
 sky130_fd_sc_hd__buf_1 _24692_ (.A(_08529_),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_2 _24693_ (.A0(_08055_),
    .A1(\fetch.bht.bhtTable_target_pc[13][3] ),
    .S(_06306_),
    .X(_08530_));
 sky130_fd_sc_hd__buf_1 _24694_ (.A(_08530_),
    .X(_02010_));
 sky130_fd_sc_hd__buf_1 _24695_ (.A(_06282_),
    .X(_08531_));
 sky130_fd_sc_hd__mux2_2 _24696_ (.A0(_08057_),
    .A1(\fetch.bht.bhtTable_target_pc[13][4] ),
    .S(_08531_),
    .X(_08532_));
 sky130_fd_sc_hd__buf_1 _24697_ (.A(_08532_),
    .X(_02011_));
 sky130_fd_sc_hd__mux2_2 _24698_ (.A0(_08060_),
    .A1(\fetch.bht.bhtTable_target_pc[13][5] ),
    .S(_08531_),
    .X(_08533_));
 sky130_fd_sc_hd__buf_1 _24699_ (.A(_08533_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_2 _24700_ (.A0(_08062_),
    .A1(\fetch.bht.bhtTable_target_pc[13][6] ),
    .S(_08531_),
    .X(_08534_));
 sky130_fd_sc_hd__buf_1 _24701_ (.A(_08534_),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_2 _24702_ (.A0(_08064_),
    .A1(\fetch.bht.bhtTable_target_pc[13][7] ),
    .S(_08531_),
    .X(_08535_));
 sky130_fd_sc_hd__buf_1 _24703_ (.A(_08535_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_2 _24704_ (.A0(_08066_),
    .A1(\fetch.bht.bhtTable_target_pc[13][8] ),
    .S(_08531_),
    .X(_08536_));
 sky130_fd_sc_hd__buf_1 _24705_ (.A(_08536_),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_2 _24706_ (.A0(_08068_),
    .A1(\fetch.bht.bhtTable_target_pc[13][9] ),
    .S(_08531_),
    .X(_08537_));
 sky130_fd_sc_hd__buf_1 _24707_ (.A(_08537_),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_2 _24708_ (.A0(_08070_),
    .A1(\fetch.bht.bhtTable_target_pc[13][10] ),
    .S(_08531_),
    .X(_08538_));
 sky130_fd_sc_hd__buf_1 _24709_ (.A(_08538_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_2 _24710_ (.A0(_08072_),
    .A1(\fetch.bht.bhtTable_target_pc[13][11] ),
    .S(_08531_),
    .X(_08539_));
 sky130_fd_sc_hd__buf_1 _24711_ (.A(_08539_),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_2 _24712_ (.A0(_08074_),
    .A1(\fetch.bht.bhtTable_target_pc[13][12] ),
    .S(_08531_),
    .X(_08540_));
 sky130_fd_sc_hd__buf_1 _24713_ (.A(_08540_),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_2 _24714_ (.A0(_08076_),
    .A1(\fetch.bht.bhtTable_target_pc[13][13] ),
    .S(_08531_),
    .X(_08541_));
 sky130_fd_sc_hd__buf_1 _24715_ (.A(_08541_),
    .X(_02020_));
 sky130_fd_sc_hd__buf_1 _24716_ (.A(_06282_),
    .X(_08542_));
 sky130_fd_sc_hd__mux2_2 _24717_ (.A0(_08078_),
    .A1(\fetch.bht.bhtTable_target_pc[13][14] ),
    .S(_08542_),
    .X(_08543_));
 sky130_fd_sc_hd__buf_1 _24718_ (.A(_08543_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_2 _24719_ (.A0(_08081_),
    .A1(\fetch.bht.bhtTable_target_pc[13][15] ),
    .S(_08542_),
    .X(_08544_));
 sky130_fd_sc_hd__buf_1 _24720_ (.A(_08544_),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_2 _24721_ (.A0(_08083_),
    .A1(\fetch.bht.bhtTable_target_pc[13][16] ),
    .S(_08542_),
    .X(_08545_));
 sky130_fd_sc_hd__buf_1 _24722_ (.A(_08545_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_2 _24723_ (.A0(_08085_),
    .A1(\fetch.bht.bhtTable_target_pc[13][17] ),
    .S(_08542_),
    .X(_08546_));
 sky130_fd_sc_hd__buf_1 _24724_ (.A(_08546_),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_2 _24725_ (.A0(_08087_),
    .A1(\fetch.bht.bhtTable_target_pc[13][18] ),
    .S(_08542_),
    .X(_08547_));
 sky130_fd_sc_hd__buf_1 _24726_ (.A(_08547_),
    .X(_02025_));
 sky130_fd_sc_hd__mux2_2 _24727_ (.A0(_08089_),
    .A1(\fetch.bht.bhtTable_target_pc[13][19] ),
    .S(_08542_),
    .X(_08548_));
 sky130_fd_sc_hd__buf_1 _24728_ (.A(_08548_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_2 _24729_ (.A0(_08091_),
    .A1(\fetch.bht.bhtTable_target_pc[13][20] ),
    .S(_08542_),
    .X(_08549_));
 sky130_fd_sc_hd__buf_1 _24730_ (.A(_08549_),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_2 _24731_ (.A0(_08093_),
    .A1(\fetch.bht.bhtTable_target_pc[13][21] ),
    .S(_08542_),
    .X(_08550_));
 sky130_fd_sc_hd__buf_1 _24732_ (.A(_08550_),
    .X(_02028_));
 sky130_fd_sc_hd__mux2_2 _24733_ (.A0(_08095_),
    .A1(\fetch.bht.bhtTable_target_pc[13][22] ),
    .S(_08542_),
    .X(_08551_));
 sky130_fd_sc_hd__buf_1 _24734_ (.A(_08551_),
    .X(_02029_));
 sky130_fd_sc_hd__mux2_2 _24735_ (.A0(_08097_),
    .A1(\fetch.bht.bhtTable_target_pc[13][23] ),
    .S(_08542_),
    .X(_08552_));
 sky130_fd_sc_hd__buf_1 _24736_ (.A(_08552_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_2 _24737_ (.A0(_08099_),
    .A1(\fetch.bht.bhtTable_target_pc[13][24] ),
    .S(_06283_),
    .X(_08553_));
 sky130_fd_sc_hd__buf_1 _24738_ (.A(_08553_),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_2 _24739_ (.A0(_08101_),
    .A1(\fetch.bht.bhtTable_target_pc[13][25] ),
    .S(_06283_),
    .X(_08554_));
 sky130_fd_sc_hd__buf_1 _24740_ (.A(_08554_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_2 _24741_ (.A0(_08103_),
    .A1(\fetch.bht.bhtTable_target_pc[13][26] ),
    .S(_06283_),
    .X(_08555_));
 sky130_fd_sc_hd__buf_1 _24742_ (.A(_08555_),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_2 _24743_ (.A0(_08105_),
    .A1(\fetch.bht.bhtTable_target_pc[13][27] ),
    .S(_06283_),
    .X(_08556_));
 sky130_fd_sc_hd__buf_1 _24744_ (.A(_08556_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_2 _24745_ (.A0(_08107_),
    .A1(\fetch.bht.bhtTable_target_pc[13][28] ),
    .S(_06283_),
    .X(_08557_));
 sky130_fd_sc_hd__buf_1 _24746_ (.A(_08557_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_2 _24747_ (.A0(_08109_),
    .A1(\fetch.bht.bhtTable_target_pc[13][29] ),
    .S(_06283_),
    .X(_08558_));
 sky130_fd_sc_hd__buf_1 _24748_ (.A(_08558_),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_2 _24749_ (.A0(_08111_),
    .A1(\fetch.bht.bhtTable_target_pc[13][30] ),
    .S(_06283_),
    .X(_08559_));
 sky130_fd_sc_hd__buf_1 _24750_ (.A(_08559_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_2 _24751_ (.A0(_08113_),
    .A1(\fetch.bht.bhtTable_target_pc[13][31] ),
    .S(_06283_),
    .X(_08560_));
 sky130_fd_sc_hd__buf_1 _24752_ (.A(_08560_),
    .X(_02038_));
 sky130_fd_sc_hd__or3b_2 _24753_ (.A(_09900_),
    .B(_06281_),
    .C_N(_09887_),
    .X(_08561_));
 sky130_fd_sc_hd__buf_1 _24754_ (.A(_08561_),
    .X(_08562_));
 sky130_fd_sc_hd__buf_1 _24755_ (.A(_08562_),
    .X(_08563_));
 sky130_fd_sc_hd__mux2_2 _24756_ (.A0(_08049_),
    .A1(\fetch.bht.bhtTable_target_pc[14][0] ),
    .S(_08563_),
    .X(_08564_));
 sky130_fd_sc_hd__buf_1 _24757_ (.A(_08564_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_2 _24758_ (.A0(_08051_),
    .A1(\fetch.bht.bhtTable_target_pc[14][1] ),
    .S(_08563_),
    .X(_08565_));
 sky130_fd_sc_hd__buf_1 _24759_ (.A(_08565_),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_2 _24760_ (.A0(_08053_),
    .A1(\fetch.bht.bhtTable_target_pc[14][2] ),
    .S(_08563_),
    .X(_08566_));
 sky130_fd_sc_hd__buf_1 _24761_ (.A(_08566_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_2 _24762_ (.A0(_08055_),
    .A1(\fetch.bht.bhtTable_target_pc[14][3] ),
    .S(_08563_),
    .X(_08567_));
 sky130_fd_sc_hd__buf_1 _24763_ (.A(_08567_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_2 _24764_ (.A0(_08057_),
    .A1(\fetch.bht.bhtTable_target_pc[14][4] ),
    .S(_08563_),
    .X(_08568_));
 sky130_fd_sc_hd__buf_1 _24765_ (.A(_08568_),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_2 _24766_ (.A0(_08060_),
    .A1(\fetch.bht.bhtTable_target_pc[14][5] ),
    .S(_08563_),
    .X(_08569_));
 sky130_fd_sc_hd__buf_1 _24767_ (.A(_08569_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_2 _24768_ (.A0(_08062_),
    .A1(\fetch.bht.bhtTable_target_pc[14][6] ),
    .S(_08563_),
    .X(_08570_));
 sky130_fd_sc_hd__buf_1 _24769_ (.A(_08570_),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_2 _24770_ (.A0(_08064_),
    .A1(\fetch.bht.bhtTable_target_pc[14][7] ),
    .S(_08563_),
    .X(_08571_));
 sky130_fd_sc_hd__buf_1 _24771_ (.A(_08571_),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_2 _24772_ (.A0(_08066_),
    .A1(\fetch.bht.bhtTable_target_pc[14][8] ),
    .S(_08563_),
    .X(_08572_));
 sky130_fd_sc_hd__buf_1 _24773_ (.A(_08572_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_2 _24774_ (.A0(_08068_),
    .A1(\fetch.bht.bhtTable_target_pc[14][9] ),
    .S(_08563_),
    .X(_08573_));
 sky130_fd_sc_hd__buf_1 _24775_ (.A(_08573_),
    .X(_02048_));
 sky130_fd_sc_hd__buf_1 _24776_ (.A(_08562_),
    .X(_08574_));
 sky130_fd_sc_hd__mux2_2 _24777_ (.A0(_08070_),
    .A1(\fetch.bht.bhtTable_target_pc[14][10] ),
    .S(_08574_),
    .X(_08575_));
 sky130_fd_sc_hd__buf_1 _24778_ (.A(_08575_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_2 _24779_ (.A0(_08072_),
    .A1(\fetch.bht.bhtTable_target_pc[14][11] ),
    .S(_08574_),
    .X(_08576_));
 sky130_fd_sc_hd__buf_1 _24780_ (.A(_08576_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_2 _24781_ (.A0(_08074_),
    .A1(\fetch.bht.bhtTable_target_pc[14][12] ),
    .S(_08574_),
    .X(_08577_));
 sky130_fd_sc_hd__buf_1 _24782_ (.A(_08577_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_2 _24783_ (.A0(_08076_),
    .A1(\fetch.bht.bhtTable_target_pc[14][13] ),
    .S(_08574_),
    .X(_08578_));
 sky130_fd_sc_hd__buf_1 _24784_ (.A(_08578_),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_2 _24785_ (.A0(_08078_),
    .A1(\fetch.bht.bhtTable_target_pc[14][14] ),
    .S(_08574_),
    .X(_08579_));
 sky130_fd_sc_hd__buf_1 _24786_ (.A(_08579_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_2 _24787_ (.A0(_08081_),
    .A1(\fetch.bht.bhtTable_target_pc[14][15] ),
    .S(_08574_),
    .X(_08580_));
 sky130_fd_sc_hd__buf_1 _24788_ (.A(_08580_),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_2 _24789_ (.A0(_08083_),
    .A1(\fetch.bht.bhtTable_target_pc[14][16] ),
    .S(_08574_),
    .X(_08581_));
 sky130_fd_sc_hd__buf_1 _24790_ (.A(_08581_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_2 _24791_ (.A0(_08085_),
    .A1(\fetch.bht.bhtTable_target_pc[14][17] ),
    .S(_08574_),
    .X(_08582_));
 sky130_fd_sc_hd__buf_1 _24792_ (.A(_08582_),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_2 _24793_ (.A0(_08087_),
    .A1(\fetch.bht.bhtTable_target_pc[14][18] ),
    .S(_08574_),
    .X(_08583_));
 sky130_fd_sc_hd__buf_1 _24794_ (.A(_08583_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_2 _24795_ (.A0(_08089_),
    .A1(\fetch.bht.bhtTable_target_pc[14][19] ),
    .S(_08574_),
    .X(_08584_));
 sky130_fd_sc_hd__buf_1 _24796_ (.A(_08584_),
    .X(_02058_));
 sky130_fd_sc_hd__buf_1 _24797_ (.A(_08561_),
    .X(_08585_));
 sky130_fd_sc_hd__mux2_2 _24798_ (.A0(_08091_),
    .A1(\fetch.bht.bhtTable_target_pc[14][20] ),
    .S(_08585_),
    .X(_08586_));
 sky130_fd_sc_hd__buf_1 _24799_ (.A(_08586_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_2 _24800_ (.A0(_08093_),
    .A1(\fetch.bht.bhtTable_target_pc[14][21] ),
    .S(_08585_),
    .X(_08587_));
 sky130_fd_sc_hd__buf_1 _24801_ (.A(_08587_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_2 _24802_ (.A0(_08095_),
    .A1(\fetch.bht.bhtTable_target_pc[14][22] ),
    .S(_08585_),
    .X(_08588_));
 sky130_fd_sc_hd__buf_1 _24803_ (.A(_08588_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_2 _24804_ (.A0(_08097_),
    .A1(\fetch.bht.bhtTable_target_pc[14][23] ),
    .S(_08585_),
    .X(_08589_));
 sky130_fd_sc_hd__buf_1 _24805_ (.A(_08589_),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_2 _24806_ (.A0(_08099_),
    .A1(\fetch.bht.bhtTable_target_pc[14][24] ),
    .S(_08585_),
    .X(_08590_));
 sky130_fd_sc_hd__buf_1 _24807_ (.A(_08590_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_2 _24808_ (.A0(_08101_),
    .A1(\fetch.bht.bhtTable_target_pc[14][25] ),
    .S(_08585_),
    .X(_08591_));
 sky130_fd_sc_hd__buf_1 _24809_ (.A(_08591_),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_2 _24810_ (.A0(_08103_),
    .A1(\fetch.bht.bhtTable_target_pc[14][26] ),
    .S(_08585_),
    .X(_08592_));
 sky130_fd_sc_hd__buf_1 _24811_ (.A(_08592_),
    .X(_02065_));
 sky130_fd_sc_hd__mux2_2 _24812_ (.A0(_08105_),
    .A1(\fetch.bht.bhtTable_target_pc[14][27] ),
    .S(_08585_),
    .X(_08593_));
 sky130_fd_sc_hd__buf_1 _24813_ (.A(_08593_),
    .X(_02066_));
 sky130_fd_sc_hd__mux2_2 _24814_ (.A0(_08107_),
    .A1(\fetch.bht.bhtTable_target_pc[14][28] ),
    .S(_08585_),
    .X(_08594_));
 sky130_fd_sc_hd__buf_1 _24815_ (.A(_08594_),
    .X(_02067_));
 sky130_fd_sc_hd__mux2_2 _24816_ (.A0(_08109_),
    .A1(\fetch.bht.bhtTable_target_pc[14][29] ),
    .S(_08585_),
    .X(_08595_));
 sky130_fd_sc_hd__buf_1 _24817_ (.A(_08595_),
    .X(_02068_));
 sky130_fd_sc_hd__buf_1 _24818_ (.A(_08561_),
    .X(_08596_));
 sky130_fd_sc_hd__mux2_2 _24819_ (.A0(_08111_),
    .A1(\fetch.bht.bhtTable_target_pc[14][30] ),
    .S(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__buf_1 _24820_ (.A(_08597_),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_2 _24821_ (.A0(_08113_),
    .A1(\fetch.bht.bhtTable_target_pc[14][31] ),
    .S(_08596_),
    .X(_08598_));
 sky130_fd_sc_hd__buf_1 _24822_ (.A(_08598_),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_2 _24823_ (.A0(_06101_),
    .A1(\fetch.bht.bhtTable_tag[0][0] ),
    .S(_08422_),
    .X(_08599_));
 sky130_fd_sc_hd__buf_1 _24824_ (.A(_08599_),
    .X(_02071_));
 sky130_fd_sc_hd__mux2_2 _24825_ (.A0(_06103_),
    .A1(\fetch.bht.bhtTable_tag[0][1] ),
    .S(_08422_),
    .X(_08600_));
 sky130_fd_sc_hd__buf_1 _24826_ (.A(_08600_),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_2 _24827_ (.A0(_06105_),
    .A1(\fetch.bht.bhtTable_tag[0][2] ),
    .S(_08422_),
    .X(_08601_));
 sky130_fd_sc_hd__buf_1 _24828_ (.A(_08601_),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_2 _24829_ (.A0(_06107_),
    .A1(\fetch.bht.bhtTable_tag[0][3] ),
    .S(_08422_),
    .X(_08602_));
 sky130_fd_sc_hd__buf_1 _24830_ (.A(_08602_),
    .X(_02074_));
 sky130_fd_sc_hd__mux2_2 _24831_ (.A0(_06109_),
    .A1(\fetch.bht.bhtTable_tag[0][4] ),
    .S(_08422_),
    .X(_08603_));
 sky130_fd_sc_hd__buf_1 _24832_ (.A(_08603_),
    .X(_02075_));
 sky130_fd_sc_hd__mux2_2 _24833_ (.A0(_06111_),
    .A1(\fetch.bht.bhtTable_tag[0][5] ),
    .S(_08422_),
    .X(_08604_));
 sky130_fd_sc_hd__buf_1 _24834_ (.A(_08604_),
    .X(_02076_));
 sky130_fd_sc_hd__mux2_2 _24835_ (.A0(_06113_),
    .A1(\fetch.bht.bhtTable_tag[0][6] ),
    .S(_08422_),
    .X(_08605_));
 sky130_fd_sc_hd__buf_1 _24836_ (.A(_08605_),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_2 _24837_ (.A0(_06115_),
    .A1(\fetch.bht.bhtTable_tag[0][7] ),
    .S(_08422_),
    .X(_08606_));
 sky130_fd_sc_hd__buf_1 _24838_ (.A(_08606_),
    .X(_02078_));
 sky130_fd_sc_hd__buf_1 _24839_ (.A(_08387_),
    .X(_08607_));
 sky130_fd_sc_hd__mux2_2 _24840_ (.A0(_06117_),
    .A1(\fetch.bht.bhtTable_tag[0][8] ),
    .S(_08607_),
    .X(_08608_));
 sky130_fd_sc_hd__buf_1 _24841_ (.A(_08608_),
    .X(_02079_));
 sky130_fd_sc_hd__mux2_2 _24842_ (.A0(_06119_),
    .A1(\fetch.bht.bhtTable_tag[0][9] ),
    .S(_08607_),
    .X(_08609_));
 sky130_fd_sc_hd__buf_1 _24843_ (.A(_08609_),
    .X(_02080_));
 sky130_fd_sc_hd__mux2_2 _24844_ (.A0(_06122_),
    .A1(\fetch.bht.bhtTable_tag[0][10] ),
    .S(_08607_),
    .X(_08610_));
 sky130_fd_sc_hd__buf_1 _24845_ (.A(_08610_),
    .X(_02081_));
 sky130_fd_sc_hd__mux2_2 _24846_ (.A0(_06124_),
    .A1(\fetch.bht.bhtTable_tag[0][11] ),
    .S(_08607_),
    .X(_08611_));
 sky130_fd_sc_hd__buf_1 _24847_ (.A(_08611_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_2 _24848_ (.A0(_06126_),
    .A1(\fetch.bht.bhtTable_tag[0][12] ),
    .S(_08607_),
    .X(_08612_));
 sky130_fd_sc_hd__buf_1 _24849_ (.A(_08612_),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_2 _24850_ (.A0(_06128_),
    .A1(\fetch.bht.bhtTable_tag[0][13] ),
    .S(_08607_),
    .X(_08613_));
 sky130_fd_sc_hd__buf_1 _24851_ (.A(_08613_),
    .X(_02084_));
 sky130_fd_sc_hd__mux2_2 _24852_ (.A0(_06130_),
    .A1(\fetch.bht.bhtTable_tag[0][14] ),
    .S(_08607_),
    .X(_08614_));
 sky130_fd_sc_hd__buf_1 _24853_ (.A(_08614_),
    .X(_02085_));
 sky130_fd_sc_hd__mux2_2 _24854_ (.A0(_06132_),
    .A1(\fetch.bht.bhtTable_tag[0][15] ),
    .S(_08607_),
    .X(_08615_));
 sky130_fd_sc_hd__buf_1 _24855_ (.A(_08615_),
    .X(_02086_));
 sky130_fd_sc_hd__mux2_2 _24856_ (.A0(_06134_),
    .A1(\fetch.bht.bhtTable_tag[0][16] ),
    .S(_08607_),
    .X(_08616_));
 sky130_fd_sc_hd__buf_1 _24857_ (.A(_08616_),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_2 _24858_ (.A0(_06136_),
    .A1(\fetch.bht.bhtTable_tag[0][17] ),
    .S(_08607_),
    .X(_08617_));
 sky130_fd_sc_hd__buf_1 _24859_ (.A(_08617_),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_2 _24860_ (.A0(_06138_),
    .A1(\fetch.bht.bhtTable_tag[0][18] ),
    .S(_08388_),
    .X(_08618_));
 sky130_fd_sc_hd__buf_1 _24861_ (.A(_08618_),
    .X(_02089_));
 sky130_fd_sc_hd__mux2_2 _24862_ (.A0(_06140_),
    .A1(\fetch.bht.bhtTable_tag[0][19] ),
    .S(_08388_),
    .X(_08619_));
 sky130_fd_sc_hd__buf_1 _24863_ (.A(_08619_),
    .X(_02090_));
 sky130_fd_sc_hd__mux2_2 _24864_ (.A0(_06143_),
    .A1(\fetch.bht.bhtTable_tag[0][20] ),
    .S(_08388_),
    .X(_08620_));
 sky130_fd_sc_hd__buf_1 _24865_ (.A(_08620_),
    .X(_02091_));
 sky130_fd_sc_hd__mux2_2 _24866_ (.A0(_06145_),
    .A1(\fetch.bht.bhtTable_tag[0][21] ),
    .S(_08388_),
    .X(_08621_));
 sky130_fd_sc_hd__buf_1 _24867_ (.A(_08621_),
    .X(_02092_));
 sky130_fd_sc_hd__mux2_2 _24868_ (.A0(_06147_),
    .A1(\fetch.bht.bhtTable_tag[0][22] ),
    .S(_08388_),
    .X(_08622_));
 sky130_fd_sc_hd__buf_1 _24869_ (.A(_08622_),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_2 _24870_ (.A0(_06149_),
    .A1(\fetch.bht.bhtTable_tag[0][23] ),
    .S(_08388_),
    .X(_08623_));
 sky130_fd_sc_hd__buf_1 _24871_ (.A(_08623_),
    .X(_02094_));
 sky130_fd_sc_hd__mux2_2 _24872_ (.A0(_06151_),
    .A1(\fetch.bht.bhtTable_tag[0][24] ),
    .S(_08388_),
    .X(_08624_));
 sky130_fd_sc_hd__buf_1 _24873_ (.A(_08624_),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_2 _24874_ (.A0(_06153_),
    .A1(\fetch.bht.bhtTable_tag[0][25] ),
    .S(_08388_),
    .X(_08625_));
 sky130_fd_sc_hd__buf_1 _24875_ (.A(_08625_),
    .X(_02096_));
 sky130_fd_sc_hd__and4_2 _24876_ (.A(\csr.mcycle[14] ),
    .B(\csr.mcycle[13] ),
    .C(\csr.mcycle[18] ),
    .D(\csr.mcycle[17] ),
    .X(_08626_));
 sky130_fd_sc_hd__and4_2 _24877_ (.A(\csr.mcycle[10] ),
    .B(\csr.mcycle[9] ),
    .C(\csr.mcycle[12] ),
    .D(\csr.mcycle[11] ),
    .X(_08627_));
 sky130_fd_sc_hd__and4_2 _24878_ (.A(\csr.mcycle[16] ),
    .B(\csr.mcycle[15] ),
    .C(_08626_),
    .D(_08627_),
    .X(_08628_));
 sky130_fd_sc_hd__and4_2 _24879_ (.A(\csr.mcycle[19] ),
    .B(\csr.mcycle[22] ),
    .C(\csr.mcycle[21] ),
    .D(\csr.mcycle[24] ),
    .X(_08629_));
 sky130_fd_sc_hd__and4_2 _24880_ (.A(\csr.mcycle[23] ),
    .B(\csr.mcycle[26] ),
    .C(\csr.mcycle[25] ),
    .D(\csr.mcycle[30] ),
    .X(_08630_));
 sky130_fd_sc_hd__and4_2 _24881_ (.A(\csr.mcycle[28] ),
    .B(\csr.mcycle[27] ),
    .C(\csr.mcycle[29] ),
    .D(_08630_),
    .X(_08631_));
 sky130_fd_sc_hd__and4_2 _24882_ (.A(\csr.mcycle[8] ),
    .B(\csr.mcycle[20] ),
    .C(_08629_),
    .D(_08631_),
    .X(_08632_));
 sky130_fd_sc_hd__nand4_2 _24883_ (.A(\csr.io_csr_write_address[11] ),
    .B(_06313_),
    .C(_06314_),
    .D(_06459_),
    .Y(_08633_));
 sky130_fd_sc_hd__and4_2 _24884_ (.A(_08633_),
    .B(_03558_),
    .C(\csr.mcycle[7] ),
    .D(\csr.mcycle[6] ),
    .X(_08634_));
 sky130_fd_sc_hd__buf_1 _24885_ (.A(_08634_),
    .X(_08635_));
 sky130_fd_sc_hd__and4_2 _24886_ (.A(\csr.mcycle[31] ),
    .B(_08628_),
    .C(_08632_),
    .D(_08635_),
    .X(_08636_));
 sky130_fd_sc_hd__a21oi_2 _24887_ (.A1(\csr._mcycle_T_3[32] ),
    .A2(_08636_),
    .B1(_07179_),
    .Y(_08637_));
 sky130_fd_sc_hd__o21a_2 _24888_ (.A1(\csr._mcycle_T_3[32] ),
    .A2(_08636_),
    .B1(_08637_),
    .X(_02097_));
 sky130_fd_sc_hd__a21oi_2 _24889_ (.A1(\csr._mcycle_T_3[32] ),
    .A2(_08636_),
    .B1(\csr._mcycle_T_3[33] ),
    .Y(_08638_));
 sky130_fd_sc_hd__and4_2 _24890_ (.A(\csr.mcycle[28] ),
    .B(\csr.mcycle[27] ),
    .C(\csr.mcycle[30] ),
    .D(\csr.mcycle[29] ),
    .X(_08639_));
 sky130_fd_sc_hd__and4_2 _24891_ (.A(_03555_),
    .B(\csr.mcycle[23] ),
    .C(\csr.mcycle[26] ),
    .D(\csr.mcycle[25] ),
    .X(_08640_));
 sky130_fd_sc_hd__and3_2 _24892_ (.A(\csr.mcycle[21] ),
    .B(\csr.mcycle[24] ),
    .C(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__and4_2 _24893_ (.A(\csr.mcycle[10] ),
    .B(\csr.mcycle[9] ),
    .C(\csr.mcycle[12] ),
    .D(\csr.mcycle[13] ),
    .X(_08642_));
 sky130_fd_sc_hd__and3_2 _24894_ (.A(\csr.mcycle[11] ),
    .B(_03559_),
    .C(_08642_),
    .X(_08643_));
 sky130_fd_sc_hd__and4_2 _24895_ (.A(_08633_),
    .B(_08643_),
    .C(_03556_),
    .D(\csr.mcycle[18] ),
    .X(_08644_));
 sky130_fd_sc_hd__and3_2 _24896_ (.A(\csr.mcycle[20] ),
    .B(_03554_),
    .C(_08644_),
    .X(_08645_));
 sky130_fd_sc_hd__and3_2 _24897_ (.A(_08639_),
    .B(_08641_),
    .C(_08645_),
    .X(_08646_));
 sky130_fd_sc_hd__and4_2 _24898_ (.A(\csr._mcycle_T_3[33] ),
    .B(\csr._mcycle_T_3[32] ),
    .C(\csr.mcycle[31] ),
    .D(_08646_),
    .X(_08647_));
 sky130_fd_sc_hd__nor3_2 _24899_ (.A(_07199_),
    .B(_08638_),
    .C(_08647_),
    .Y(_02098_));
 sky130_fd_sc_hd__a21oi_2 _24900_ (.A1(\csr._mcycle_T_3[34] ),
    .A2(_08647_),
    .B1(_07179_),
    .Y(_08648_));
 sky130_fd_sc_hd__o21a_2 _24901_ (.A1(\csr._mcycle_T_3[34] ),
    .A2(_08647_),
    .B1(_08648_),
    .X(_02099_));
 sky130_fd_sc_hd__and4_2 _24902_ (.A(\csr._mcycle_T_3[34] ),
    .B(\csr._mcycle_T_3[33] ),
    .C(\csr._mcycle_T_3[32] ),
    .D(_08636_),
    .X(_08649_));
 sky130_fd_sc_hd__a21oi_2 _24903_ (.A1(\csr._mcycle_T_3[35] ),
    .A2(_08649_),
    .B1(_07179_),
    .Y(_08650_));
 sky130_fd_sc_hd__o21a_2 _24904_ (.A1(\csr._mcycle_T_3[35] ),
    .A2(_08649_),
    .B1(_08650_),
    .X(_02100_));
 sky130_fd_sc_hd__a21oi_2 _24905_ (.A1(\csr._mcycle_T_3[35] ),
    .A2(_08649_),
    .B1(\csr._mcycle_T_3[36] ),
    .Y(_08651_));
 sky130_fd_sc_hd__and4_2 _24906_ (.A(\csr._mcycle_T_3[36] ),
    .B(\csr._mcycle_T_3[35] ),
    .C(\csr._mcycle_T_3[34] ),
    .D(_08647_),
    .X(_08652_));
 sky130_fd_sc_hd__nor3_2 _24907_ (.A(_07199_),
    .B(_08651_),
    .C(_08652_),
    .Y(_02101_));
 sky130_fd_sc_hd__a21oi_2 _24908_ (.A1(\csr._mcycle_T_3[37] ),
    .A2(_08652_),
    .B1(_07179_),
    .Y(_08653_));
 sky130_fd_sc_hd__o21a_2 _24909_ (.A1(\csr._mcycle_T_3[37] ),
    .A2(_08652_),
    .B1(_08653_),
    .X(_02102_));
 sky130_fd_sc_hd__and4_2 _24910_ (.A(\csr._mcycle_T_3[37] ),
    .B(\csr._mcycle_T_3[36] ),
    .C(\csr._mcycle_T_3[35] ),
    .D(_08649_),
    .X(_08654_));
 sky130_fd_sc_hd__a21oi_2 _24911_ (.A1(\csr._mcycle_T_3[38] ),
    .A2(_08654_),
    .B1(_07179_),
    .Y(_08655_));
 sky130_fd_sc_hd__o21a_2 _24912_ (.A1(\csr._mcycle_T_3[38] ),
    .A2(_08654_),
    .B1(_08655_),
    .X(_02103_));
 sky130_fd_sc_hd__and3_2 _24913_ (.A(\csr._mcycle_T_3[38] ),
    .B(\csr._mcycle_T_3[37] ),
    .C(_08652_),
    .X(_08656_));
 sky130_fd_sc_hd__a31o_2 _24914_ (.A1(\csr._mcycle_T_3[39] ),
    .A2(\csr._mcycle_T_3[38] ),
    .A3(_08654_),
    .B1(_06422_),
    .X(_08657_));
 sky130_fd_sc_hd__o21ba_2 _24915_ (.A1(\csr._mcycle_T_3[39] ),
    .A2(_08656_),
    .B1_N(_08657_),
    .X(_02104_));
 sky130_fd_sc_hd__a21oi_2 _24916_ (.A1(\csr._mcycle_T_3[39] ),
    .A2(_08656_),
    .B1(\csr._mcycle_T_3[40] ),
    .Y(_08658_));
 sky130_fd_sc_hd__and4_2 _24917_ (.A(\csr._mcycle_T_3[40] ),
    .B(\csr._mcycle_T_3[39] ),
    .C(\csr._mcycle_T_3[38] ),
    .D(_08654_),
    .X(_08659_));
 sky130_fd_sc_hd__nor3_2 _24918_ (.A(_07199_),
    .B(_08658_),
    .C(_08659_),
    .Y(_02105_));
 sky130_fd_sc_hd__a41o_2 _24919_ (.A1(\csr._mcycle_T_3[41] ),
    .A2(\csr._mcycle_T_3[40] ),
    .A3(\csr._mcycle_T_3[39] ),
    .A4(_08656_),
    .B1(_07148_),
    .X(_08660_));
 sky130_fd_sc_hd__o21ba_2 _24920_ (.A1(\csr._mcycle_T_3[41] ),
    .A2(_08659_),
    .B1_N(_08660_),
    .X(_02106_));
 sky130_fd_sc_hd__and4_2 _24921_ (.A(\csr._mcycle_T_3[41] ),
    .B(\csr._mcycle_T_3[40] ),
    .C(\csr._mcycle_T_3[39] ),
    .D(_08656_),
    .X(_08661_));
 sky130_fd_sc_hd__and3_2 _24922_ (.A(\csr._mcycle_T_3[42] ),
    .B(\csr._mcycle_T_3[41] ),
    .C(_08659_),
    .X(_08662_));
 sky130_fd_sc_hd__nor2_2 _24923_ (.A(_06318_),
    .B(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__o21a_2 _24924_ (.A1(\csr._mcycle_T_3[42] ),
    .A2(_08661_),
    .B1(_08663_),
    .X(_02107_));
 sky130_fd_sc_hd__a21oi_2 _24925_ (.A1(\csr._mcycle_T_3[43] ),
    .A2(_08662_),
    .B1(_06318_),
    .Y(_08664_));
 sky130_fd_sc_hd__o21a_2 _24926_ (.A1(\csr._mcycle_T_3[43] ),
    .A2(_08662_),
    .B1(_08664_),
    .X(_02108_));
 sky130_fd_sc_hd__and3_2 _24927_ (.A(\csr._mcycle_T_3[43] ),
    .B(\csr._mcycle_T_3[42] ),
    .C(_08661_),
    .X(_08665_));
 sky130_fd_sc_hd__a21oi_2 _24928_ (.A1(\csr._mcycle_T_3[44] ),
    .A2(_08665_),
    .B1(_06318_),
    .Y(_08666_));
 sky130_fd_sc_hd__o21a_2 _24929_ (.A1(\csr._mcycle_T_3[44] ),
    .A2(_08665_),
    .B1(_08666_),
    .X(_02109_));
 sky130_fd_sc_hd__a21oi_2 _24930_ (.A1(\csr._mcycle_T_3[44] ),
    .A2(_08665_),
    .B1(\csr._mcycle_T_3[45] ),
    .Y(_08667_));
 sky130_fd_sc_hd__and4_2 _24931_ (.A(\csr._mcycle_T_3[45] ),
    .B(\csr._mcycle_T_3[44] ),
    .C(\csr._mcycle_T_3[43] ),
    .D(_08662_),
    .X(_08668_));
 sky130_fd_sc_hd__nor3_2 _24932_ (.A(_07199_),
    .B(_08667_),
    .C(_08668_),
    .Y(_02110_));
 sky130_fd_sc_hd__a21oi_2 _24933_ (.A1(\csr._mcycle_T_3[46] ),
    .A2(_08668_),
    .B1(_06318_),
    .Y(_08669_));
 sky130_fd_sc_hd__o21a_2 _24934_ (.A1(\csr._mcycle_T_3[46] ),
    .A2(_08668_),
    .B1(_08669_),
    .X(_02111_));
 sky130_fd_sc_hd__and4_2 _24935_ (.A(\csr._mcycle_T_3[46] ),
    .B(\csr._mcycle_T_3[45] ),
    .C(\csr._mcycle_T_3[44] ),
    .D(_08665_),
    .X(_08670_));
 sky130_fd_sc_hd__a31o_2 _24936_ (.A1(\csr._mcycle_T_3[47] ),
    .A2(\csr._mcycle_T_3[46] ),
    .A3(_08668_),
    .B1(_06422_),
    .X(_08671_));
 sky130_fd_sc_hd__o21ba_2 _24937_ (.A1(\csr._mcycle_T_3[47] ),
    .A2(_08670_),
    .B1_N(_08671_),
    .X(_02112_));
 sky130_fd_sc_hd__and3_2 _24938_ (.A(\csr._mcycle_T_3[47] ),
    .B(\csr._mcycle_T_3[46] ),
    .C(_08668_),
    .X(_08672_));
 sky130_fd_sc_hd__a41o_2 _24939_ (.A1(\csr._mcycle_T_3[48] ),
    .A2(\csr._mcycle_T_3[47] ),
    .A3(\csr._mcycle_T_3[46] ),
    .A4(_08668_),
    .B1(_03579_),
    .X(_08673_));
 sky130_fd_sc_hd__o21ba_2 _24940_ (.A1(\csr._mcycle_T_3[48] ),
    .A2(_08672_),
    .B1_N(_08673_),
    .X(_02113_));
 sky130_fd_sc_hd__and3_2 _24941_ (.A(\csr._mcycle_T_3[48] ),
    .B(\csr._mcycle_T_3[47] ),
    .C(_08670_),
    .X(_08674_));
 sky130_fd_sc_hd__a31o_2 _24942_ (.A1(\csr._mcycle_T_3[49] ),
    .A2(\csr._mcycle_T_3[48] ),
    .A3(_08672_),
    .B1(_07148_),
    .X(_08675_));
 sky130_fd_sc_hd__o21ba_2 _24943_ (.A1(\csr._mcycle_T_3[49] ),
    .A2(_08674_),
    .B1_N(_08675_),
    .X(_02114_));
 sky130_fd_sc_hd__and3_2 _24944_ (.A(\csr._mcycle_T_3[49] ),
    .B(\csr._mcycle_T_3[48] ),
    .C(_08672_),
    .X(_08676_));
 sky130_fd_sc_hd__a21oi_2 _24945_ (.A1(\csr._mcycle_T_3[50] ),
    .A2(_08676_),
    .B1(_06318_),
    .Y(_08677_));
 sky130_fd_sc_hd__o21a_2 _24946_ (.A1(\csr._mcycle_T_3[50] ),
    .A2(_08676_),
    .B1(_08677_),
    .X(_02115_));
 sky130_fd_sc_hd__and3_2 _24947_ (.A(\csr._mcycle_T_3[50] ),
    .B(\csr._mcycle_T_3[49] ),
    .C(_08674_),
    .X(_08678_));
 sky130_fd_sc_hd__a31o_2 _24948_ (.A1(\csr._mcycle_T_3[51] ),
    .A2(\csr._mcycle_T_3[50] ),
    .A3(_08676_),
    .B1(_07148_),
    .X(_08679_));
 sky130_fd_sc_hd__o21ba_2 _24949_ (.A1(\csr._mcycle_T_3[51] ),
    .A2(_08678_),
    .B1_N(_08679_),
    .X(_02116_));
 sky130_fd_sc_hd__a21oi_2 _24950_ (.A1(\csr._mcycle_T_3[51] ),
    .A2(_08678_),
    .B1(\csr._mcycle_T_3[52] ),
    .Y(_08680_));
 sky130_fd_sc_hd__and4_2 _24951_ (.A(\csr._mcycle_T_3[52] ),
    .B(\csr._mcycle_T_3[51] ),
    .C(\csr._mcycle_T_3[50] ),
    .D(_08676_),
    .X(_08681_));
 sky130_fd_sc_hd__buf_1 _24952_ (.A(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__nor3_2 _24953_ (.A(_07199_),
    .B(_08680_),
    .C(_08682_),
    .Y(_02117_));
 sky130_fd_sc_hd__a21oi_2 _24954_ (.A1(\csr._mcycle_T_3[53] ),
    .A2(_08682_),
    .B1(_06318_),
    .Y(_08683_));
 sky130_fd_sc_hd__o21a_2 _24955_ (.A1(\csr._mcycle_T_3[53] ),
    .A2(_08682_),
    .B1(_08683_),
    .X(_02118_));
 sky130_fd_sc_hd__a21oi_2 _24956_ (.A1(\csr._mcycle_T_3[53] ),
    .A2(_08682_),
    .B1(\csr._mcycle_T_3[54] ),
    .Y(_08684_));
 sky130_fd_sc_hd__and3_2 _24957_ (.A(\csr._mcycle_T_3[54] ),
    .B(\csr._mcycle_T_3[53] ),
    .C(_08682_),
    .X(_08685_));
 sky130_fd_sc_hd__nor3_2 _24958_ (.A(_07199_),
    .B(_08684_),
    .C(_08685_),
    .Y(_02119_));
 sky130_fd_sc_hd__a41o_2 _24959_ (.A1(\csr._mcycle_T_3[55] ),
    .A2(\csr._mcycle_T_3[54] ),
    .A3(\csr._mcycle_T_3[53] ),
    .A4(_08682_),
    .B1(_03579_),
    .X(_08686_));
 sky130_fd_sc_hd__o21ba_2 _24960_ (.A1(\csr._mcycle_T_3[55] ),
    .A2(_08685_),
    .B1_N(_08686_),
    .X(_02120_));
 sky130_fd_sc_hd__and4_2 _24961_ (.A(\csr._mcycle_T_3[55] ),
    .B(\csr._mcycle_T_3[54] ),
    .C(\csr._mcycle_T_3[53] ),
    .D(_08682_),
    .X(_08687_));
 sky130_fd_sc_hd__a31o_2 _24962_ (.A1(\csr._mcycle_T_3[56] ),
    .A2(\csr._mcycle_T_3[55] ),
    .A3(_08685_),
    .B1(_07148_),
    .X(_08688_));
 sky130_fd_sc_hd__o21ba_2 _24963_ (.A1(\csr._mcycle_T_3[56] ),
    .A2(_08687_),
    .B1_N(_08688_),
    .X(_02121_));
 sky130_fd_sc_hd__and3_2 _24964_ (.A(\csr._mcycle_T_3[56] ),
    .B(\csr._mcycle_T_3[55] ),
    .C(_08685_),
    .X(_08689_));
 sky130_fd_sc_hd__a31o_2 _24965_ (.A1(\csr._mcycle_T_3[57] ),
    .A2(\csr._mcycle_T_3[56] ),
    .A3(_08687_),
    .B1(_07148_),
    .X(_08690_));
 sky130_fd_sc_hd__o21ba_2 _24966_ (.A1(\csr._mcycle_T_3[57] ),
    .A2(_08689_),
    .B1_N(_08690_),
    .X(_02122_));
 sky130_fd_sc_hd__a21oi_2 _24967_ (.A1(\csr._mcycle_T_3[57] ),
    .A2(_08689_),
    .B1(\csr._mcycle_T_3[58] ),
    .Y(_08691_));
 sky130_fd_sc_hd__and3_2 _24968_ (.A(\csr._mcycle_T_3[58] ),
    .B(\csr._mcycle_T_3[57] ),
    .C(_08689_),
    .X(_08692_));
 sky130_fd_sc_hd__buf_1 _24969_ (.A(_08692_),
    .X(_08693_));
 sky130_fd_sc_hd__nor3_2 _24970_ (.A(_07199_),
    .B(_08691_),
    .C(_08693_),
    .Y(_02123_));
 sky130_fd_sc_hd__a21oi_2 _24971_ (.A1(\csr._mcycle_T_3[59] ),
    .A2(_08693_),
    .B1(_06318_),
    .Y(_08694_));
 sky130_fd_sc_hd__o21a_2 _24972_ (.A1(\csr._mcycle_T_3[59] ),
    .A2(_08693_),
    .B1(_08694_),
    .X(_02124_));
 sky130_fd_sc_hd__a21oi_2 _24973_ (.A1(\csr._mcycle_T_3[59] ),
    .A2(_08693_),
    .B1(\csr._mcycle_T_3[60] ),
    .Y(_08695_));
 sky130_fd_sc_hd__and3_2 _24974_ (.A(\csr._mcycle_T_3[60] ),
    .B(\csr._mcycle_T_3[59] ),
    .C(_08693_),
    .X(_08696_));
 sky130_fd_sc_hd__nor3_2 _24975_ (.A(_07199_),
    .B(_08695_),
    .C(_08696_),
    .Y(_02125_));
 sky130_fd_sc_hd__a41o_2 _24976_ (.A1(\csr._mcycle_T_3[61] ),
    .A2(\csr._mcycle_T_3[60] ),
    .A3(\csr._mcycle_T_3[59] ),
    .A4(_08693_),
    .B1(_03579_),
    .X(_08697_));
 sky130_fd_sc_hd__o21ba_2 _24977_ (.A1(\csr._mcycle_T_3[61] ),
    .A2(_08696_),
    .B1_N(_08697_),
    .X(_02126_));
 sky130_fd_sc_hd__a21oi_2 _24978_ (.A1(\csr._mcycle_T_3[61] ),
    .A2(_08696_),
    .B1(\csr._mcycle_T_3[62] ),
    .Y(_08698_));
 sky130_fd_sc_hd__and3_2 _24979_ (.A(\csr._mcycle_T_3[62] ),
    .B(\csr._mcycle_T_3[61] ),
    .C(_08696_),
    .X(_08699_));
 sky130_fd_sc_hd__nor3_2 _24980_ (.A(_06331_),
    .B(_08698_),
    .C(_08699_),
    .Y(_02127_));
 sky130_fd_sc_hd__a41o_2 _24981_ (.A1(\csr._mcycle_T_3[63] ),
    .A2(\csr._mcycle_T_3[62] ),
    .A3(\csr._mcycle_T_3[61] ),
    .A4(_08696_),
    .B1(_03579_),
    .X(_08700_));
 sky130_fd_sc_hd__o21ba_2 _24982_ (.A1(\csr._mcycle_T_3[63] ),
    .A2(_08699_),
    .B1_N(_08700_),
    .X(_02128_));
 sky130_fd_sc_hd__buf_1 _24983_ (.A(_08633_),
    .X(_08701_));
 sky130_fd_sc_hd__a21oi_2 _24984_ (.A1(_08701_),
    .A2(\csr.mcycle[0] ),
    .B1(_06318_),
    .Y(_08702_));
 sky130_fd_sc_hd__o31a_2 _24985_ (.A1(\csr._mcycle_T_2[0] ),
    .A2(\csr.mcycle[0] ),
    .A3(_08701_),
    .B1(_08702_),
    .X(_02129_));
 sky130_fd_sc_hd__and4_2 _24986_ (.A(\csr.io_csr_write_address[11] ),
    .B(_06313_),
    .C(_06314_),
    .D(_06459_),
    .X(_08703_));
 sky130_fd_sc_hd__buf_1 _24987_ (.A(_08703_),
    .X(_08704_));
 sky130_fd_sc_hd__a21o_2 _24988_ (.A1(_08633_),
    .A2(\csr.mcycle[0] ),
    .B1(\csr.mcycle[1] ),
    .X(_08705_));
 sky130_fd_sc_hd__a21oi_2 _24989_ (.A1(\csr._mcycle_T_2[1] ),
    .A2(_08704_),
    .B1(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__a311oi_2 _24990_ (.A1(\csr.mcycle[0] ),
    .A2(_08701_),
    .A3(\csr.mcycle[1] ),
    .B1(_06318_),
    .C1(_08706_),
    .Y(_02130_));
 sky130_fd_sc_hd__a31o_2 _24991_ (.A1(_08701_),
    .A2(\csr.mcycle[1] ),
    .A3(\csr.mcycle[0] ),
    .B1(\csr.mcycle[2] ),
    .X(_08707_));
 sky130_fd_sc_hd__a21oi_2 _24992_ (.A1(\csr._mcycle_T_2[2] ),
    .A2(_08704_),
    .B1(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__a211oi_2 _24993_ (.A1(_08701_),
    .A2(_03557_),
    .B1(_06327_),
    .C1(_08708_),
    .Y(_02131_));
 sky130_fd_sc_hd__and4_2 _24994_ (.A(_08633_),
    .B(\csr.mcycle[1] ),
    .C(\csr.mcycle[2] ),
    .D(\csr.mcycle[0] ),
    .X(_08709_));
 sky130_fd_sc_hd__buf_1 _24995_ (.A(_08703_),
    .X(_08710_));
 sky130_fd_sc_hd__a211oi_2 _24996_ (.A1(\csr._mcycle_T_2[3] ),
    .A2(_08710_),
    .B1(_08709_),
    .C1(\csr.mcycle[3] ),
    .Y(_08711_));
 sky130_fd_sc_hd__a211oi_2 _24997_ (.A1(\csr.mcycle[3] ),
    .A2(_08709_),
    .B1(_08711_),
    .C1(_06419_),
    .Y(_02132_));
 sky130_fd_sc_hd__buf_1 _24998_ (.A(_08703_),
    .X(_08712_));
 sky130_fd_sc_hd__a221oi_2 _24999_ (.A1(\csr._mcycle_T_2[4] ),
    .A2(_08712_),
    .B1(_08709_),
    .B2(\csr.mcycle[3] ),
    .C1(\csr.mcycle[4] ),
    .Y(_08713_));
 sky130_fd_sc_hd__a311oi_2 _25000_ (.A1(\csr.mcycle[4] ),
    .A2(\csr.mcycle[3] ),
    .A3(_08709_),
    .B1(_08713_),
    .C1(_06336_),
    .Y(_02133_));
 sky130_fd_sc_hd__a31oi_2 _25001_ (.A1(\csr.mcycle[4] ),
    .A2(\csr.mcycle[3] ),
    .A3(_03557_),
    .B1(\csr.mcycle[5] ),
    .Y(_08714_));
 sky130_fd_sc_hd__o21ai_2 _25002_ (.A1(_03558_),
    .A2(_08714_),
    .B1(_08701_),
    .Y(_08715_));
 sky130_fd_sc_hd__o311a_2 _25003_ (.A1(\csr._mcycle_T_2[5] ),
    .A2(\csr.mcycle[5] ),
    .A3(_08701_),
    .B1(_08715_),
    .C1(_05856_),
    .X(_02134_));
 sky130_fd_sc_hd__nand2_2 _25004_ (.A(\csr.mcycle[6] ),
    .B(_03558_),
    .Y(_08716_));
 sky130_fd_sc_hd__a41o_2 _25005_ (.A1(\csr.mcycle[4] ),
    .A2(\csr.mcycle[3] ),
    .A3(\csr.mcycle[5] ),
    .A4(_03557_),
    .B1(\csr.mcycle[6] ),
    .X(_08717_));
 sky130_fd_sc_hd__a21o_2 _25006_ (.A1(_08716_),
    .A2(_08717_),
    .B1(_08704_),
    .X(_08718_));
 sky130_fd_sc_hd__o311a_2 _25007_ (.A1(\csr._mcycle_T_2[6] ),
    .A2(_08701_),
    .A3(\csr.mcycle[6] ),
    .B1(_05856_),
    .C1(_08718_),
    .X(_02135_));
 sky130_fd_sc_hd__a31o_2 _25008_ (.A1(_08701_),
    .A2(_03558_),
    .A3(\csr.mcycle[6] ),
    .B1(\csr.mcycle[7] ),
    .X(_08719_));
 sky130_fd_sc_hd__a21oi_2 _25009_ (.A1(\csr._mcycle_T_2[7] ),
    .A2(_08704_),
    .B1(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__nor3_2 _25010_ (.A(_06331_),
    .B(_08635_),
    .C(_08720_),
    .Y(_02136_));
 sky130_fd_sc_hd__a211oi_2 _25011_ (.A1(\csr._mcycle_T_2[8] ),
    .A2(_08710_),
    .B1(_08635_),
    .C1(\csr.mcycle[8] ),
    .Y(_08721_));
 sky130_fd_sc_hd__a211oi_2 _25012_ (.A1(\csr.mcycle[8] ),
    .A2(_08635_),
    .B1(_08721_),
    .C1(_06419_),
    .Y(_02137_));
 sky130_fd_sc_hd__and4bb_2 _25013_ (.A_N(_08703_),
    .B_N(_08716_),
    .C(\csr.mcycle[7] ),
    .D(\csr.mcycle[8] ),
    .X(_08722_));
 sky130_fd_sc_hd__a221oi_2 _25014_ (.A1(\csr._mcycle_T_2[9] ),
    .A2(_08712_),
    .B1(_08635_),
    .B2(\csr.mcycle[8] ),
    .C1(\csr.mcycle[9] ),
    .Y(_08723_));
 sky130_fd_sc_hd__a211oi_2 _25015_ (.A1(\csr.mcycle[9] ),
    .A2(_08722_),
    .B1(_08723_),
    .C1(_06419_),
    .Y(_02138_));
 sky130_fd_sc_hd__a221oi_2 _25016_ (.A1(\csr._mcycle_T_2[10] ),
    .A2(_08712_),
    .B1(_08722_),
    .B2(\csr.mcycle[9] ),
    .C1(\csr.mcycle[10] ),
    .Y(_08724_));
 sky130_fd_sc_hd__and4_2 _25017_ (.A(\csr.mcycle[8] ),
    .B(\csr.mcycle[10] ),
    .C(\csr.mcycle[9] ),
    .D(_08635_),
    .X(_08725_));
 sky130_fd_sc_hd__nor3_2 _25018_ (.A(_06331_),
    .B(_08724_),
    .C(_08725_),
    .Y(_02139_));
 sky130_fd_sc_hd__a211o_2 _25019_ (.A1(\csr._mcycle_T_2[11] ),
    .A2(_08712_),
    .B1(_08725_),
    .C1(\csr.mcycle[11] ),
    .X(_08726_));
 sky130_fd_sc_hd__nand2_2 _25020_ (.A(\csr.mcycle[11] ),
    .B(_08725_),
    .Y(_08727_));
 sky130_fd_sc_hd__and3_2 _25021_ (.A(_10019_),
    .B(_08726_),
    .C(_08727_),
    .X(_08728_));
 sky130_fd_sc_hd__buf_1 _25022_ (.A(_08728_),
    .X(_02140_));
 sky130_fd_sc_hd__a21oi_2 _25023_ (.A1(\csr._mcycle_T_2[12] ),
    .A2(_08704_),
    .B1(\csr.mcycle[12] ),
    .Y(_08729_));
 sky130_fd_sc_hd__and3_2 _25024_ (.A(\csr.mcycle[12] ),
    .B(\csr.mcycle[11] ),
    .C(_08725_),
    .X(_08730_));
 sky130_fd_sc_hd__a211oi_2 _25025_ (.A1(_08729_),
    .A2(_08727_),
    .B1(_06327_),
    .C1(_08730_),
    .Y(_02141_));
 sky130_fd_sc_hd__a211oi_2 _25026_ (.A1(\csr._mcycle_T_2[13] ),
    .A2(_08710_),
    .B1(_08730_),
    .C1(\csr.mcycle[13] ),
    .Y(_08731_));
 sky130_fd_sc_hd__a211oi_2 _25027_ (.A1(\csr.mcycle[13] ),
    .A2(_08730_),
    .B1(_08731_),
    .C1(_06419_),
    .Y(_02142_));
 sky130_fd_sc_hd__a221oi_2 _25028_ (.A1(\csr._mcycle_T_2[14] ),
    .A2(_08712_),
    .B1(_08730_),
    .B2(\csr.mcycle[13] ),
    .C1(\csr.mcycle[14] ),
    .Y(_08732_));
 sky130_fd_sc_hd__and3_2 _25029_ (.A(\csr.mcycle[14] ),
    .B(\csr.mcycle[13] ),
    .C(_08730_),
    .X(_08733_));
 sky130_fd_sc_hd__nor3_2 _25030_ (.A(_06331_),
    .B(_08732_),
    .C(_08733_),
    .Y(_02143_));
 sky130_fd_sc_hd__a211o_2 _25031_ (.A1(\csr._mcycle_T_2[15] ),
    .A2(_08712_),
    .B1(_08733_),
    .C1(\csr.mcycle[15] ),
    .X(_08734_));
 sky130_fd_sc_hd__nand2_2 _25032_ (.A(\csr.mcycle[15] ),
    .B(_08733_),
    .Y(_08735_));
 sky130_fd_sc_hd__and3_2 _25033_ (.A(_10019_),
    .B(_08734_),
    .C(_08735_),
    .X(_08736_));
 sky130_fd_sc_hd__buf_1 _25034_ (.A(_08736_),
    .X(_02144_));
 sky130_fd_sc_hd__a21oi_2 _25035_ (.A1(\csr._mcycle_T_2[16] ),
    .A2(_08704_),
    .B1(\csr.mcycle[16] ),
    .Y(_08737_));
 sky130_fd_sc_hd__and3_2 _25036_ (.A(\csr.mcycle[16] ),
    .B(\csr.mcycle[15] ),
    .C(_08733_),
    .X(_08738_));
 sky130_fd_sc_hd__a211oi_2 _25037_ (.A1(_08737_),
    .A2(_08735_),
    .B1(_06327_),
    .C1(_08738_),
    .Y(_02145_));
 sky130_fd_sc_hd__a211oi_2 _25038_ (.A1(\csr._mcycle_T_2[17] ),
    .A2(_08710_),
    .B1(_08738_),
    .C1(\csr.mcycle[17] ),
    .Y(_08739_));
 sky130_fd_sc_hd__a211oi_2 _25039_ (.A1(\csr.mcycle[17] ),
    .A2(_08738_),
    .B1(_08739_),
    .C1(_06419_),
    .Y(_02146_));
 sky130_fd_sc_hd__and3_2 _25040_ (.A(_03556_),
    .B(_03561_),
    .C(_08633_),
    .X(_08740_));
 sky130_fd_sc_hd__a211oi_2 _25041_ (.A1(\csr._mcycle_T_2[18] ),
    .A2(_08704_),
    .B1(_08740_),
    .C1(\csr.mcycle[18] ),
    .Y(_08741_));
 sky130_fd_sc_hd__a211oi_2 _25042_ (.A1(_08701_),
    .A2(_03562_),
    .B1(_06327_),
    .C1(_08741_),
    .Y(_02147_));
 sky130_fd_sc_hd__and3_2 _25043_ (.A(\csr.mcycle[8] ),
    .B(_08628_),
    .C(_08635_),
    .X(_08742_));
 sky130_fd_sc_hd__a211oi_2 _25044_ (.A1(\csr._mcycle_T_2[19] ),
    .A2(_08710_),
    .B1(_08742_),
    .C1(_03554_),
    .Y(_08743_));
 sky130_fd_sc_hd__a211oi_2 _25045_ (.A1(_03554_),
    .A2(_08644_),
    .B1(_08743_),
    .C1(_06419_),
    .Y(_02148_));
 sky130_fd_sc_hd__a221oi_2 _25046_ (.A1(\csr._mcycle_T_2[20] ),
    .A2(_08712_),
    .B1(_08742_),
    .B2(_03554_),
    .C1(\csr.mcycle[20] ),
    .Y(_08744_));
 sky130_fd_sc_hd__and4_2 _25047_ (.A(_08633_),
    .B(_03562_),
    .C(_03554_),
    .D(\csr.mcycle[20] ),
    .X(_08745_));
 sky130_fd_sc_hd__nor3_2 _25048_ (.A(_06331_),
    .B(_08744_),
    .C(_08745_),
    .Y(_02149_));
 sky130_fd_sc_hd__a211oi_2 _25049_ (.A1(\csr._mcycle_T_2[21] ),
    .A2(_08710_),
    .B1(_08645_),
    .C1(\csr.mcycle[21] ),
    .Y(_08746_));
 sky130_fd_sc_hd__a211oi_2 _25050_ (.A1(\csr.mcycle[21] ),
    .A2(_08645_),
    .B1(_08746_),
    .C1(_06419_),
    .Y(_02150_));
 sky130_fd_sc_hd__and4_2 _25051_ (.A(\csr.mcycle[20] ),
    .B(_03554_),
    .C(\csr.mcycle[21] ),
    .D(_08644_),
    .X(_08747_));
 sky130_fd_sc_hd__and4_2 _25052_ (.A(\csr.mcycle[20] ),
    .B(_03554_),
    .C(\csr.mcycle[21] ),
    .D(_08742_),
    .X(_08748_));
 sky130_fd_sc_hd__a211oi_2 _25053_ (.A1(\csr._mcycle_T_2[22] ),
    .A2(_08710_),
    .B1(_08748_),
    .C1(_03555_),
    .Y(_08749_));
 sky130_fd_sc_hd__a211oi_2 _25054_ (.A1(_03555_),
    .A2(_08747_),
    .B1(_08749_),
    .C1(_06419_),
    .Y(_02151_));
 sky130_fd_sc_hd__a21oi_2 _25055_ (.A1(_03555_),
    .A2(_08748_),
    .B1(\csr.mcycle[23] ),
    .Y(_08750_));
 sky130_fd_sc_hd__and3_2 _25056_ (.A(_03555_),
    .B(\csr.mcycle[23] ),
    .C(_08747_),
    .X(_08751_));
 sky130_fd_sc_hd__o2bb2a_2 _25057_ (.A1_N(\csr._mcycle_T_2[23] ),
    .A2_N(_08704_),
    .B1(_08750_),
    .B2(_08751_),
    .X(_08752_));
 sky130_fd_sc_hd__nor2_2 _25058_ (.A(_03580_),
    .B(_08752_),
    .Y(_02152_));
 sky130_fd_sc_hd__a211oi_2 _25059_ (.A1(\csr._mcycle_T_2[24] ),
    .A2(_08710_),
    .B1(_08751_),
    .C1(\csr.mcycle[24] ),
    .Y(_08753_));
 sky130_fd_sc_hd__a211oi_2 _25060_ (.A1(\csr.mcycle[24] ),
    .A2(_08751_),
    .B1(_08753_),
    .C1(_06327_),
    .Y(_02153_));
 sky130_fd_sc_hd__and4_2 _25061_ (.A(_03555_),
    .B(\csr.mcycle[24] ),
    .C(\csr.mcycle[23] ),
    .D(_08748_),
    .X(_08754_));
 sky130_fd_sc_hd__a211oi_2 _25062_ (.A1(\csr._mcycle_T_2[25] ),
    .A2(_08710_),
    .B1(_08754_),
    .C1(\csr.mcycle[25] ),
    .Y(_08755_));
 sky130_fd_sc_hd__a211oi_2 _25063_ (.A1(\csr.mcycle[25] ),
    .A2(_08754_),
    .B1(_08755_),
    .C1(_06327_),
    .Y(_02154_));
 sky130_fd_sc_hd__and3_2 _25064_ (.A(_03555_),
    .B(\csr.mcycle[21] ),
    .C(_08745_),
    .X(_08756_));
 sky130_fd_sc_hd__and3_2 _25065_ (.A(\csr.mcycle[24] ),
    .B(\csr.mcycle[23] ),
    .C(_08756_),
    .X(_08757_));
 sky130_fd_sc_hd__a221oi_2 _25066_ (.A1(\csr._mcycle_T_2[26] ),
    .A2(_08712_),
    .B1(_08757_),
    .B2(\csr.mcycle[25] ),
    .C1(\csr.mcycle[26] ),
    .Y(_08758_));
 sky130_fd_sc_hd__and3_2 _25067_ (.A(\csr.mcycle[26] ),
    .B(\csr.mcycle[25] ),
    .C(_08754_),
    .X(_08759_));
 sky130_fd_sc_hd__nor3_2 _25068_ (.A(_06331_),
    .B(_08758_),
    .C(_08759_),
    .Y(_02155_));
 sky130_fd_sc_hd__a211oi_2 _25069_ (.A1(\csr._mcycle_T_2[27] ),
    .A2(_08712_),
    .B1(_08759_),
    .C1(\csr.mcycle[27] ),
    .Y(_08760_));
 sky130_fd_sc_hd__a211oi_2 _25070_ (.A1(\csr.mcycle[27] ),
    .A2(_08759_),
    .B1(_08760_),
    .C1(_06327_),
    .Y(_02156_));
 sky130_fd_sc_hd__and4_2 _25071_ (.A(\csr.mcycle[26] ),
    .B(\csr.mcycle[25] ),
    .C(\csr.mcycle[27] ),
    .D(_08757_),
    .X(_08761_));
 sky130_fd_sc_hd__a211o_2 _25072_ (.A1(\csr._mcycle_T_2[28] ),
    .A2(_08703_),
    .B1(_08761_),
    .C1(\csr.mcycle[28] ),
    .X(_08762_));
 sky130_fd_sc_hd__nand2_2 _25073_ (.A(\csr.mcycle[28] ),
    .B(_08761_),
    .Y(_08763_));
 sky130_fd_sc_hd__and3_2 _25074_ (.A(_10019_),
    .B(_08762_),
    .C(_08763_),
    .X(_08764_));
 sky130_fd_sc_hd__buf_1 _25075_ (.A(_08764_),
    .X(_02157_));
 sky130_fd_sc_hd__a31oi_2 _25076_ (.A1(\csr.mcycle[28] ),
    .A2(\csr.mcycle[27] ),
    .A3(_08759_),
    .B1(\csr.mcycle[29] ),
    .Y(_08765_));
 sky130_fd_sc_hd__and4_2 _25077_ (.A(\csr.mcycle[28] ),
    .B(\csr.mcycle[27] ),
    .C(\csr.mcycle[29] ),
    .D(_08759_),
    .X(_08766_));
 sky130_fd_sc_hd__o2bb2a_2 _25078_ (.A1_N(\csr._mcycle_T_2[29] ),
    .A2_N(_08710_),
    .B1(_08765_),
    .B2(_08766_),
    .X(_08767_));
 sky130_fd_sc_hd__nor2_2 _25079_ (.A(_03580_),
    .B(_08767_),
    .Y(_02158_));
 sky130_fd_sc_hd__a211o_2 _25080_ (.A1(\csr._mcycle_T_2[30] ),
    .A2(_08704_),
    .B1(_08766_),
    .C1(\csr.mcycle[30] ),
    .X(_08768_));
 sky130_fd_sc_hd__o211a_2 _25081_ (.A1(_08704_),
    .A2(_03567_),
    .B1(_06566_),
    .C1(_08768_),
    .X(_02159_));
 sky130_fd_sc_hd__a211oi_2 _25082_ (.A1(\csr._mcycle_T_2[31] ),
    .A2(_08712_),
    .B1(_08646_),
    .C1(\csr.mcycle[31] ),
    .Y(_08769_));
 sky130_fd_sc_hd__a211oi_2 _25083_ (.A1(\csr.mcycle[31] ),
    .A2(_08646_),
    .B1(_08769_),
    .C1(_06327_),
    .Y(_02160_));
 sky130_fd_sc_hd__mux2_2 _25084_ (.A0(_06101_),
    .A1(\fetch.bht.bhtTable_tag[14][0] ),
    .S(_08596_),
    .X(_08770_));
 sky130_fd_sc_hd__buf_1 _25085_ (.A(_08770_),
    .X(_02161_));
 sky130_fd_sc_hd__mux2_2 _25086_ (.A0(_06103_),
    .A1(\fetch.bht.bhtTable_tag[14][1] ),
    .S(_08596_),
    .X(_08771_));
 sky130_fd_sc_hd__buf_1 _25087_ (.A(_08771_),
    .X(_02162_));
 sky130_fd_sc_hd__mux2_2 _25088_ (.A0(_06105_),
    .A1(\fetch.bht.bhtTable_tag[14][2] ),
    .S(_08596_),
    .X(_08772_));
 sky130_fd_sc_hd__buf_1 _25089_ (.A(_08772_),
    .X(_02163_));
 sky130_fd_sc_hd__mux2_2 _25090_ (.A0(_06107_),
    .A1(\fetch.bht.bhtTable_tag[14][3] ),
    .S(_08596_),
    .X(_08773_));
 sky130_fd_sc_hd__buf_1 _25091_ (.A(_08773_),
    .X(_02164_));
 sky130_fd_sc_hd__mux2_2 _25092_ (.A0(_06109_),
    .A1(\fetch.bht.bhtTable_tag[14][4] ),
    .S(_08596_),
    .X(_08774_));
 sky130_fd_sc_hd__buf_1 _25093_ (.A(_08774_),
    .X(_02165_));
 sky130_fd_sc_hd__mux2_2 _25094_ (.A0(_06111_),
    .A1(\fetch.bht.bhtTable_tag[14][5] ),
    .S(_08596_),
    .X(_08775_));
 sky130_fd_sc_hd__buf_1 _25095_ (.A(_08775_),
    .X(_02166_));
 sky130_fd_sc_hd__mux2_2 _25096_ (.A0(_06113_),
    .A1(\fetch.bht.bhtTable_tag[14][6] ),
    .S(_08596_),
    .X(_08776_));
 sky130_fd_sc_hd__buf_1 _25097_ (.A(_08776_),
    .X(_02167_));
 sky130_fd_sc_hd__mux2_2 _25098_ (.A0(_06115_),
    .A1(\fetch.bht.bhtTable_tag[14][7] ),
    .S(_08596_),
    .X(_08777_));
 sky130_fd_sc_hd__buf_1 _25099_ (.A(_08777_),
    .X(_02168_));
 sky130_fd_sc_hd__buf_1 _25100_ (.A(_08561_),
    .X(_08778_));
 sky130_fd_sc_hd__mux2_2 _25101_ (.A0(_06117_),
    .A1(\fetch.bht.bhtTable_tag[14][8] ),
    .S(_08778_),
    .X(_08779_));
 sky130_fd_sc_hd__buf_1 _25102_ (.A(_08779_),
    .X(_02169_));
 sky130_fd_sc_hd__mux2_2 _25103_ (.A0(_06119_),
    .A1(\fetch.bht.bhtTable_tag[14][9] ),
    .S(_08778_),
    .X(_08780_));
 sky130_fd_sc_hd__buf_1 _25104_ (.A(_08780_),
    .X(_02170_));
 sky130_fd_sc_hd__mux2_2 _25105_ (.A0(_06122_),
    .A1(\fetch.bht.bhtTable_tag[14][10] ),
    .S(_08778_),
    .X(_08781_));
 sky130_fd_sc_hd__buf_1 _25106_ (.A(_08781_),
    .X(_02171_));
 sky130_fd_sc_hd__mux2_2 _25107_ (.A0(_06124_),
    .A1(\fetch.bht.bhtTable_tag[14][11] ),
    .S(_08778_),
    .X(_08782_));
 sky130_fd_sc_hd__buf_1 _25108_ (.A(_08782_),
    .X(_02172_));
 sky130_fd_sc_hd__mux2_2 _25109_ (.A0(_06126_),
    .A1(\fetch.bht.bhtTable_tag[14][12] ),
    .S(_08778_),
    .X(_08783_));
 sky130_fd_sc_hd__buf_1 _25110_ (.A(_08783_),
    .X(_02173_));
 sky130_fd_sc_hd__mux2_2 _25111_ (.A0(_06128_),
    .A1(\fetch.bht.bhtTable_tag[14][13] ),
    .S(_08778_),
    .X(_08784_));
 sky130_fd_sc_hd__buf_1 _25112_ (.A(_08784_),
    .X(_02174_));
 sky130_fd_sc_hd__mux2_2 _25113_ (.A0(_06130_),
    .A1(\fetch.bht.bhtTable_tag[14][14] ),
    .S(_08778_),
    .X(_08785_));
 sky130_fd_sc_hd__buf_1 _25114_ (.A(_08785_),
    .X(_02175_));
 sky130_fd_sc_hd__mux2_2 _25115_ (.A0(_06132_),
    .A1(\fetch.bht.bhtTable_tag[14][15] ),
    .S(_08778_),
    .X(_08786_));
 sky130_fd_sc_hd__buf_1 _25116_ (.A(_08786_),
    .X(_02176_));
 sky130_fd_sc_hd__mux2_2 _25117_ (.A0(_06134_),
    .A1(\fetch.bht.bhtTable_tag[14][16] ),
    .S(_08778_),
    .X(_08787_));
 sky130_fd_sc_hd__buf_1 _25118_ (.A(_08787_),
    .X(_02177_));
 sky130_fd_sc_hd__mux2_2 _25119_ (.A0(_06136_),
    .A1(\fetch.bht.bhtTable_tag[14][17] ),
    .S(_08778_),
    .X(_08788_));
 sky130_fd_sc_hd__buf_1 _25120_ (.A(_08788_),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_2 _25121_ (.A0(_06138_),
    .A1(\fetch.bht.bhtTable_tag[14][18] ),
    .S(_08562_),
    .X(_08789_));
 sky130_fd_sc_hd__buf_1 _25122_ (.A(_08789_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_2 _25123_ (.A0(_06140_),
    .A1(\fetch.bht.bhtTable_tag[14][19] ),
    .S(_08562_),
    .X(_08790_));
 sky130_fd_sc_hd__buf_1 _25124_ (.A(_08790_),
    .X(_02180_));
 sky130_fd_sc_hd__mux2_2 _25125_ (.A0(_06143_),
    .A1(\fetch.bht.bhtTable_tag[14][20] ),
    .S(_08562_),
    .X(_08791_));
 sky130_fd_sc_hd__buf_1 _25126_ (.A(_08791_),
    .X(_02181_));
 sky130_fd_sc_hd__mux2_2 _25127_ (.A0(_06145_),
    .A1(\fetch.bht.bhtTable_tag[14][21] ),
    .S(_08562_),
    .X(_08792_));
 sky130_fd_sc_hd__buf_1 _25128_ (.A(_08792_),
    .X(_02182_));
 sky130_fd_sc_hd__mux2_2 _25129_ (.A0(_06147_),
    .A1(\fetch.bht.bhtTable_tag[14][22] ),
    .S(_08562_),
    .X(_08793_));
 sky130_fd_sc_hd__buf_1 _25130_ (.A(_08793_),
    .X(_02183_));
 sky130_fd_sc_hd__mux2_2 _25131_ (.A0(_06149_),
    .A1(\fetch.bht.bhtTable_tag[14][23] ),
    .S(_08562_),
    .X(_08794_));
 sky130_fd_sc_hd__buf_1 _25132_ (.A(_08794_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_2 _25133_ (.A0(_06151_),
    .A1(\fetch.bht.bhtTable_tag[14][24] ),
    .S(_08562_),
    .X(_08795_));
 sky130_fd_sc_hd__buf_1 _25134_ (.A(_08795_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_2 _25135_ (.A0(_06153_),
    .A1(\fetch.bht.bhtTable_tag[14][25] ),
    .S(_08562_),
    .X(_08796_));
 sky130_fd_sc_hd__buf_1 _25136_ (.A(_08796_),
    .X(_02186_));
 sky130_fd_sc_hd__a211o_2 _25137_ (.A1(_03526_),
    .A2(_03521_),
    .B1(_03524_),
    .C1(_07250_),
    .X(_08797_));
 sky130_fd_sc_hd__and3_2 _25138_ (.A(_08797_),
    .B(_03535_),
    .C(\decode.control.io_funct7[5] ),
    .X(_08798_));
 sky130_fd_sc_hd__o311a_2 _25139_ (.A1(_03528_),
    .A2(_07250_),
    .A3(_08798_),
    .B1(_10998_),
    .C1(_03458_),
    .X(_08799_));
 sky130_fd_sc_hd__a31o_2 _25140_ (.A1(_10946_),
    .A2(_10944_),
    .A3(_00461_),
    .B1(_08799_),
    .X(_02187_));
 sky130_fd_sc_hd__and4b_2 _25141_ (.A_N(_10946_),
    .B(_10944_),
    .C(_10964_),
    .D(_10665_),
    .X(_08800_));
 sky130_fd_sc_hd__o21a_2 _25142_ (.A1(_10949_),
    .A2(_08800_),
    .B1(_10999_),
    .X(_02188_));
 sky130_fd_sc_hd__o311a_2 _25143_ (.A1(io_fetch_address[2]),
    .A2(_06248_),
    .A3(_10916_),
    .B1(_07383_),
    .C1(_05856_),
    .X(_02189_));
 sky130_fd_sc_hd__a211o_2 _25144_ (.A1(io_fetch_address[3]),
    .A2(_07348_),
    .B1(_07399_),
    .C1(_03580_),
    .X(_02190_));
 sky130_fd_sc_hd__o311a_2 _25145_ (.A1(io_fetch_address[4]),
    .A2(_06248_),
    .A3(_10916_),
    .B1(_07415_),
    .C1(_05856_),
    .X(_02191_));
 sky130_fd_sc_hd__o31a_2 _25146_ (.A1(io_fetch_address[5]),
    .A2(_07343_),
    .A3(_07344_),
    .B1(_07432_),
    .X(_02192_));
 sky130_fd_sc_hd__nand2_2 _25147_ (.A(_10568_),
    .B(_09887_),
    .Y(_08801_));
 sky130_fd_sc_hd__or2_2 _25148_ (.A(_06281_),
    .B(_08801_),
    .X(_08802_));
 sky130_fd_sc_hd__xnor2_2 _25149_ (.A(\fetch.btb.btbTable[14][0] ),
    .B(_08802_),
    .Y(_02193_));
 sky130_fd_sc_hd__mux2_2 _25150_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[14][1] ),
    .S(_08802_),
    .X(_08803_));
 sky130_fd_sc_hd__buf_1 _25151_ (.A(_08803_),
    .X(_02194_));
 sky130_fd_sc_hd__or2_2 _25152_ (.A(_06281_),
    .B(_10569_),
    .X(_08804_));
 sky130_fd_sc_hd__xnor2_2 _25153_ (.A(\fetch.btb.btbTable[13][0] ),
    .B(_08804_),
    .Y(_02195_));
 sky130_fd_sc_hd__mux2_2 _25154_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[13][1] ),
    .S(_08804_),
    .X(_08805_));
 sky130_fd_sc_hd__buf_1 _25155_ (.A(_08805_),
    .X(_02196_));
 sky130_fd_sc_hd__or4b_2 _25156_ (.A(_10556_),
    .B(_10557_),
    .C(_06281_),
    .D_N(_10568_),
    .X(_08806_));
 sky130_fd_sc_hd__xnor2_2 _25157_ (.A(\fetch.btb.btbTable[12][0] ),
    .B(_08806_),
    .Y(_02197_));
 sky130_fd_sc_hd__mux2_2 _25158_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[12][1] ),
    .S(_08806_),
    .X(_08807_));
 sky130_fd_sc_hd__buf_1 _25159_ (.A(_08807_),
    .X(_02198_));
 sky130_fd_sc_hd__nand2_2 _25160_ (.A(_10568_),
    .B(_09894_),
    .Y(_08808_));
 sky130_fd_sc_hd__or3b_2 _25161_ (.A(_08808_),
    .B(_09881_),
    .C_N(_09884_),
    .X(_08809_));
 sky130_fd_sc_hd__xnor2_2 _25162_ (.A(\fetch.btb.btbTable[11][0] ),
    .B(_08809_),
    .Y(_02199_));
 sky130_fd_sc_hd__mux2_2 _25163_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[11][1] ),
    .S(_08809_),
    .X(_08810_));
 sky130_fd_sc_hd__buf_1 _25164_ (.A(_08810_),
    .X(_02200_));
 sky130_fd_sc_hd__or3b_2 _25165_ (.A(_08801_),
    .B(_09880_),
    .C_N(_09884_),
    .X(_08811_));
 sky130_fd_sc_hd__xnor2_2 _25166_ (.A(\fetch.btb.btbTable[10][0] ),
    .B(_08811_),
    .Y(_02201_));
 sky130_fd_sc_hd__mux2_2 _25167_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[10][1] ),
    .S(_08811_),
    .X(_08812_));
 sky130_fd_sc_hd__buf_1 _25168_ (.A(_08812_),
    .X(_02202_));
 sky130_fd_sc_hd__or3b_2 _25169_ (.A(_10556_),
    .B(_10557_),
    .C_N(_10568_),
    .X(_08813_));
 sky130_fd_sc_hd__or3_2 _25170_ (.A(_09880_),
    .B(_09883_),
    .C(_08813_),
    .X(_08814_));
 sky130_fd_sc_hd__xnor2_2 _25171_ (.A(\fetch.btb.btbTable[0][0] ),
    .B(_08814_),
    .Y(_02203_));
 sky130_fd_sc_hd__mux2_2 _25172_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[0][1] ),
    .S(_08814_),
    .X(_08815_));
 sky130_fd_sc_hd__buf_1 _25173_ (.A(_08815_),
    .X(_02204_));
 sky130_fd_sc_hd__or3b_2 _25174_ (.A(_08813_),
    .B(_09880_),
    .C_N(_09884_),
    .X(_08816_));
 sky130_fd_sc_hd__xnor2_2 _25175_ (.A(\fetch.btb.btbTable[8][0] ),
    .B(_08816_),
    .Y(_02205_));
 sky130_fd_sc_hd__mux2_2 _25176_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[8][1] ),
    .S(_08816_),
    .X(_08817_));
 sky130_fd_sc_hd__buf_1 _25177_ (.A(_08817_),
    .X(_02206_));
 sky130_fd_sc_hd__or3b_2 _25178_ (.A(_09884_),
    .B(_08808_),
    .C_N(_09881_),
    .X(_08818_));
 sky130_fd_sc_hd__xnor2_2 _25179_ (.A(\fetch.btb.btbTable[7][0] ),
    .B(_08818_),
    .Y(_02207_));
 sky130_fd_sc_hd__mux2_2 _25180_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[7][1] ),
    .S(_08818_),
    .X(_08819_));
 sky130_fd_sc_hd__buf_1 _25181_ (.A(_08819_),
    .X(_02208_));
 sky130_fd_sc_hd__or3b_2 _25182_ (.A(_09883_),
    .B(_08801_),
    .C_N(_09881_),
    .X(_08820_));
 sky130_fd_sc_hd__xnor2_2 _25183_ (.A(\fetch.btb.btbTable[6][0] ),
    .B(_08820_),
    .Y(_02209_));
 sky130_fd_sc_hd__mux2_2 _25184_ (.A0(_10573_),
    .A1(\fetch.btb.btbTable[6][1] ),
    .S(_08820_),
    .X(_08821_));
 sky130_fd_sc_hd__buf_1 _25185_ (.A(_08821_),
    .X(_02210_));
 sky130_fd_sc_hd__or3b_2 _25186_ (.A(_09883_),
    .B(_10569_),
    .C_N(_09881_),
    .X(_08822_));
 sky130_fd_sc_hd__xnor2_2 _25187_ (.A(\fetch.btb.btbTable[5][0] ),
    .B(_08822_),
    .Y(_02211_));
 sky130_fd_sc_hd__mux2_2 _25188_ (.A0(_10572_),
    .A1(\fetch.btb.btbTable[5][1] ),
    .S(_08822_),
    .X(_08823_));
 sky130_fd_sc_hd__buf_1 _25189_ (.A(_08823_),
    .X(_02212_));
 sky130_fd_sc_hd__or3b_2 _25190_ (.A(_09883_),
    .B(_08813_),
    .C_N(_09881_),
    .X(_08824_));
 sky130_fd_sc_hd__xnor2_2 _25191_ (.A(\fetch.btb.btbTable[4][0] ),
    .B(_08824_),
    .Y(_02213_));
 sky130_fd_sc_hd__mux2_2 _25192_ (.A0(_10572_),
    .A1(\fetch.btb.btbTable[4][1] ),
    .S(_08824_),
    .X(_08825_));
 sky130_fd_sc_hd__buf_1 _25193_ (.A(_08825_),
    .X(_02214_));
 sky130_fd_sc_hd__or3_2 _25194_ (.A(_09880_),
    .B(_09883_),
    .C(_08808_),
    .X(_08826_));
 sky130_fd_sc_hd__xnor2_2 _25195_ (.A(\fetch.btb.btbTable[3][0] ),
    .B(_08826_),
    .Y(_02215_));
 sky130_fd_sc_hd__mux2_2 _25196_ (.A0(_10572_),
    .A1(\fetch.btb.btbTable[3][1] ),
    .S(_08826_),
    .X(_08827_));
 sky130_fd_sc_hd__buf_1 _25197_ (.A(_08827_),
    .X(_02216_));
 sky130_fd_sc_hd__or3_2 _25198_ (.A(_09880_),
    .B(_09883_),
    .C(_08801_),
    .X(_08828_));
 sky130_fd_sc_hd__xnor2_2 _25199_ (.A(\fetch.btb.btbTable[2][0] ),
    .B(_08828_),
    .Y(_02217_));
 sky130_fd_sc_hd__mux2_2 _25200_ (.A0(_10572_),
    .A1(\fetch.btb.btbTable[2][1] ),
    .S(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__buf_1 _25201_ (.A(_08829_),
    .X(_02218_));
 sky130_fd_sc_hd__or3_2 _25202_ (.A(_09880_),
    .B(_09883_),
    .C(_10569_),
    .X(_08830_));
 sky130_fd_sc_hd__xnor2_2 _25203_ (.A(\fetch.btb.btbTable[1][0] ),
    .B(_08830_),
    .Y(_02219_));
 sky130_fd_sc_hd__mux2_2 _25204_ (.A0(_10572_),
    .A1(\fetch.btb.btbTable[1][1] ),
    .S(_08830_),
    .X(_08831_));
 sky130_fd_sc_hd__buf_1 _25205_ (.A(_08831_),
    .X(_02220_));
 sky130_fd_sc_hd__nand2_2 _25206_ (.A(_10568_),
    .B(_10815_),
    .Y(_08832_));
 sky130_fd_sc_hd__xnor2_2 _25207_ (.A(\fetch.btb.btbTable[15][0] ),
    .B(_08832_),
    .Y(_02221_));
 sky130_fd_sc_hd__mux2_2 _25208_ (.A0(_10572_),
    .A1(\fetch.btb.btbTable[15][1] ),
    .S(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__buf_1 _25209_ (.A(_08833_),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_2 _25210_ (.A0(_08049_),
    .A1(\fetch.bht.bhtTable_target_pc[9][0] ),
    .S(_08041_),
    .X(_08834_));
 sky130_fd_sc_hd__buf_1 _25211_ (.A(_08834_),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_2 _25212_ (.A0(_08051_),
    .A1(\fetch.bht.bhtTable_target_pc[9][1] ),
    .S(_08041_),
    .X(_08835_));
 sky130_fd_sc_hd__buf_1 _25213_ (.A(_08835_),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_2 _25214_ (.A0(_08053_),
    .A1(\fetch.bht.bhtTable_target_pc[9][2] ),
    .S(_08041_),
    .X(_08836_));
 sky130_fd_sc_hd__buf_1 _25215_ (.A(_08836_),
    .X(_02225_));
 sky130_fd_sc_hd__buf_1 _25216_ (.A(_09905_),
    .X(_08837_));
 sky130_fd_sc_hd__mux2_2 _25217_ (.A0(_08055_),
    .A1(\fetch.bht.bhtTable_target_pc[9][3] ),
    .S(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__buf_1 _25218_ (.A(_08838_),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_2 _25219_ (.A0(_08057_),
    .A1(\fetch.bht.bhtTable_target_pc[9][4] ),
    .S(_08837_),
    .X(_08839_));
 sky130_fd_sc_hd__buf_1 _25220_ (.A(_08839_),
    .X(_02227_));
 sky130_fd_sc_hd__mux2_2 _25221_ (.A0(_08060_),
    .A1(\fetch.bht.bhtTable_target_pc[9][5] ),
    .S(_08837_),
    .X(_08840_));
 sky130_fd_sc_hd__buf_1 _25222_ (.A(_08840_),
    .X(_02228_));
 sky130_fd_sc_hd__mux2_2 _25223_ (.A0(_08062_),
    .A1(\fetch.bht.bhtTable_target_pc[9][6] ),
    .S(_08837_),
    .X(_08841_));
 sky130_fd_sc_hd__buf_1 _25224_ (.A(_08841_),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_2 _25225_ (.A0(_08064_),
    .A1(\fetch.bht.bhtTable_target_pc[9][7] ),
    .S(_08837_),
    .X(_08842_));
 sky130_fd_sc_hd__buf_1 _25226_ (.A(_08842_),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_2 _25227_ (.A0(_08066_),
    .A1(\fetch.bht.bhtTable_target_pc[9][8] ),
    .S(_08837_),
    .X(_08843_));
 sky130_fd_sc_hd__buf_1 _25228_ (.A(_08843_),
    .X(_02231_));
 sky130_fd_sc_hd__mux2_2 _25229_ (.A0(_08068_),
    .A1(\fetch.bht.bhtTable_target_pc[9][9] ),
    .S(_08837_),
    .X(_08844_));
 sky130_fd_sc_hd__buf_1 _25230_ (.A(_08844_),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_2 _25231_ (.A0(_08070_),
    .A1(\fetch.bht.bhtTable_target_pc[9][10] ),
    .S(_08837_),
    .X(_08845_));
 sky130_fd_sc_hd__buf_1 _25232_ (.A(_08845_),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_2 _25233_ (.A0(_08072_),
    .A1(\fetch.bht.bhtTable_target_pc[9][11] ),
    .S(_08837_),
    .X(_08846_));
 sky130_fd_sc_hd__buf_1 _25234_ (.A(_08846_),
    .X(_02234_));
 sky130_fd_sc_hd__mux2_2 _25235_ (.A0(_08074_),
    .A1(\fetch.bht.bhtTable_target_pc[9][12] ),
    .S(_08837_),
    .X(_08847_));
 sky130_fd_sc_hd__buf_1 _25236_ (.A(_08847_),
    .X(_02235_));
 sky130_fd_sc_hd__buf_1 _25237_ (.A(_09905_),
    .X(_08848_));
 sky130_fd_sc_hd__mux2_2 _25238_ (.A0(_08076_),
    .A1(\fetch.bht.bhtTable_target_pc[9][13] ),
    .S(_08848_),
    .X(_08849_));
 sky130_fd_sc_hd__buf_1 _25239_ (.A(_08849_),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_2 _25240_ (.A0(_08078_),
    .A1(\fetch.bht.bhtTable_target_pc[9][14] ),
    .S(_08848_),
    .X(_08850_));
 sky130_fd_sc_hd__buf_1 _25241_ (.A(_08850_),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_2 _25242_ (.A0(_08081_),
    .A1(\fetch.bht.bhtTable_target_pc[9][15] ),
    .S(_08848_),
    .X(_08851_));
 sky130_fd_sc_hd__buf_1 _25243_ (.A(_08851_),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_2 _25244_ (.A0(_08083_),
    .A1(\fetch.bht.bhtTable_target_pc[9][16] ),
    .S(_08848_),
    .X(_08852_));
 sky130_fd_sc_hd__buf_1 _25245_ (.A(_08852_),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_2 _25246_ (.A0(_08085_),
    .A1(\fetch.bht.bhtTable_target_pc[9][17] ),
    .S(_08848_),
    .X(_08853_));
 sky130_fd_sc_hd__buf_1 _25247_ (.A(_08853_),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_2 _25248_ (.A0(_08087_),
    .A1(\fetch.bht.bhtTable_target_pc[9][18] ),
    .S(_08848_),
    .X(_08854_));
 sky130_fd_sc_hd__buf_1 _25249_ (.A(_08854_),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_2 _25250_ (.A0(_08089_),
    .A1(\fetch.bht.bhtTable_target_pc[9][19] ),
    .S(_08848_),
    .X(_08855_));
 sky130_fd_sc_hd__buf_1 _25251_ (.A(_08855_),
    .X(_02242_));
 sky130_fd_sc_hd__mux2_2 _25252_ (.A0(_08091_),
    .A1(\fetch.bht.bhtTable_target_pc[9][20] ),
    .S(_08848_),
    .X(_08856_));
 sky130_fd_sc_hd__buf_1 _25253_ (.A(_08856_),
    .X(_02243_));
 sky130_fd_sc_hd__mux2_2 _25254_ (.A0(_08093_),
    .A1(\fetch.bht.bhtTable_target_pc[9][21] ),
    .S(_08848_),
    .X(_08857_));
 sky130_fd_sc_hd__buf_1 _25255_ (.A(_08857_),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_2 _25256_ (.A0(_08095_),
    .A1(\fetch.bht.bhtTable_target_pc[9][22] ),
    .S(_08848_),
    .X(_08858_));
 sky130_fd_sc_hd__buf_1 _25257_ (.A(_08858_),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_2 _25258_ (.A0(_08097_),
    .A1(\fetch.bht.bhtTable_target_pc[9][23] ),
    .S(_09906_),
    .X(_08859_));
 sky130_fd_sc_hd__buf_1 _25259_ (.A(_08859_),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_2 _25260_ (.A0(_08099_),
    .A1(\fetch.bht.bhtTable_target_pc[9][24] ),
    .S(_09906_),
    .X(_08860_));
 sky130_fd_sc_hd__buf_1 _25261_ (.A(_08860_),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_2 _25262_ (.A0(_08101_),
    .A1(\fetch.bht.bhtTable_target_pc[9][25] ),
    .S(_09906_),
    .X(_08861_));
 sky130_fd_sc_hd__buf_1 _25263_ (.A(_08861_),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_2 _25264_ (.A0(_08103_),
    .A1(\fetch.bht.bhtTable_target_pc[9][26] ),
    .S(_09906_),
    .X(_08862_));
 sky130_fd_sc_hd__buf_1 _25265_ (.A(_08862_),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_2 _25266_ (.A0(_08105_),
    .A1(\fetch.bht.bhtTable_target_pc[9][27] ),
    .S(_09906_),
    .X(_08863_));
 sky130_fd_sc_hd__buf_1 _25267_ (.A(_08863_),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_2 _25268_ (.A0(_08107_),
    .A1(\fetch.bht.bhtTable_target_pc[9][28] ),
    .S(_09906_),
    .X(_08864_));
 sky130_fd_sc_hd__buf_1 _25269_ (.A(_08864_),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_2 _25270_ (.A0(_08109_),
    .A1(\fetch.bht.bhtTable_target_pc[9][29] ),
    .S(_09906_),
    .X(_08865_));
 sky130_fd_sc_hd__buf_1 _25271_ (.A(_08865_),
    .X(_02252_));
 sky130_fd_sc_hd__mux2_2 _25272_ (.A0(_08111_),
    .A1(\fetch.bht.bhtTable_target_pc[9][30] ),
    .S(_09906_),
    .X(_08866_));
 sky130_fd_sc_hd__buf_1 _25273_ (.A(_08866_),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_2 _25274_ (.A0(_08113_),
    .A1(\fetch.bht.bhtTable_target_pc[9][31] ),
    .S(_09906_),
    .X(_08867_));
 sky130_fd_sc_hd__buf_1 _25275_ (.A(_08867_),
    .X(_02254_));
 sky130_fd_sc_hd__and2_2 _25276_ (.A(_05856_),
    .B(\decode.regfile.registers_0[0] ),
    .X(_08868_));
 sky130_fd_sc_hd__buf_1 _25277_ (.A(_08868_),
    .X(_02255_));
 sky130_fd_sc_hd__buf_1 _25278_ (.A(_10018_),
    .X(_08869_));
 sky130_fd_sc_hd__and2_2 _25279_ (.A(_08869_),
    .B(\decode.regfile.registers_0[1] ),
    .X(_08870_));
 sky130_fd_sc_hd__buf_1 _25280_ (.A(_08870_),
    .X(_02256_));
 sky130_fd_sc_hd__and2_2 _25281_ (.A(_08869_),
    .B(\decode.regfile.registers_0[2] ),
    .X(_08871_));
 sky130_fd_sc_hd__buf_1 _25282_ (.A(_08871_),
    .X(_02257_));
 sky130_fd_sc_hd__and2_2 _25283_ (.A(_08869_),
    .B(\decode.regfile.registers_0[3] ),
    .X(_08872_));
 sky130_fd_sc_hd__buf_1 _25284_ (.A(_08872_),
    .X(_02258_));
 sky130_fd_sc_hd__and2_2 _25285_ (.A(_08869_),
    .B(\decode.regfile.registers_0[4] ),
    .X(_08873_));
 sky130_fd_sc_hd__buf_1 _25286_ (.A(_08873_),
    .X(_02259_));
 sky130_fd_sc_hd__and2_2 _25287_ (.A(_08869_),
    .B(\decode.regfile.registers_0[5] ),
    .X(_08874_));
 sky130_fd_sc_hd__buf_1 _25288_ (.A(_08874_),
    .X(_02260_));
 sky130_fd_sc_hd__and2_2 _25289_ (.A(_08869_),
    .B(\decode.regfile.registers_0[6] ),
    .X(_08875_));
 sky130_fd_sc_hd__buf_1 _25290_ (.A(_08875_),
    .X(_02261_));
 sky130_fd_sc_hd__and2_2 _25291_ (.A(_08869_),
    .B(\decode.regfile.registers_0[7] ),
    .X(_08876_));
 sky130_fd_sc_hd__buf_1 _25292_ (.A(_08876_),
    .X(_02262_));
 sky130_fd_sc_hd__and2_2 _25293_ (.A(_08869_),
    .B(\decode.regfile.registers_0[8] ),
    .X(_08877_));
 sky130_fd_sc_hd__buf_1 _25294_ (.A(_08877_),
    .X(_02263_));
 sky130_fd_sc_hd__and2_2 _25295_ (.A(_08869_),
    .B(\decode.regfile.registers_0[9] ),
    .X(_08878_));
 sky130_fd_sc_hd__buf_1 _25296_ (.A(_08878_),
    .X(_02264_));
 sky130_fd_sc_hd__and2_2 _25297_ (.A(_08869_),
    .B(\decode.regfile.registers_0[10] ),
    .X(_08879_));
 sky130_fd_sc_hd__buf_1 _25298_ (.A(_08879_),
    .X(_02265_));
 sky130_fd_sc_hd__buf_1 _25299_ (.A(_10018_),
    .X(_08880_));
 sky130_fd_sc_hd__and2_2 _25300_ (.A(_08880_),
    .B(\decode.regfile.registers_0[11] ),
    .X(_08881_));
 sky130_fd_sc_hd__buf_1 _25301_ (.A(_08881_),
    .X(_02266_));
 sky130_fd_sc_hd__and2_2 _25302_ (.A(_08880_),
    .B(\decode.regfile.registers_0[12] ),
    .X(_08882_));
 sky130_fd_sc_hd__buf_1 _25303_ (.A(_08882_),
    .X(_02267_));
 sky130_fd_sc_hd__and2_2 _25304_ (.A(_08880_),
    .B(\decode.regfile.registers_0[13] ),
    .X(_08883_));
 sky130_fd_sc_hd__buf_1 _25305_ (.A(_08883_),
    .X(_02268_));
 sky130_fd_sc_hd__nor2_2 _25306_ (.A(_03580_),
    .B(_11842_),
    .Y(_02269_));
 sky130_fd_sc_hd__and2_2 _25307_ (.A(_08880_),
    .B(\decode.regfile.registers_0[15] ),
    .X(_08884_));
 sky130_fd_sc_hd__buf_1 _25308_ (.A(_08884_),
    .X(_02270_));
 sky130_fd_sc_hd__and2_2 _25309_ (.A(_08880_),
    .B(\decode.regfile.registers_0[16] ),
    .X(_08885_));
 sky130_fd_sc_hd__buf_1 _25310_ (.A(_08885_),
    .X(_02271_));
 sky130_fd_sc_hd__and2_2 _25311_ (.A(_08880_),
    .B(\decode.regfile.registers_0[17] ),
    .X(_08886_));
 sky130_fd_sc_hd__buf_1 _25312_ (.A(_08886_),
    .X(_02272_));
 sky130_fd_sc_hd__and2_2 _25313_ (.A(_08880_),
    .B(\decode.regfile.registers_0[18] ),
    .X(_08887_));
 sky130_fd_sc_hd__buf_1 _25314_ (.A(_08887_),
    .X(_02273_));
 sky130_fd_sc_hd__and2_2 _25315_ (.A(_08880_),
    .B(\decode.regfile.registers_0[19] ),
    .X(_08888_));
 sky130_fd_sc_hd__buf_1 _25316_ (.A(_08888_),
    .X(_02274_));
 sky130_fd_sc_hd__and2_2 _25317_ (.A(_08880_),
    .B(\decode.regfile.registers_0[20] ),
    .X(_08889_));
 sky130_fd_sc_hd__buf_1 _25318_ (.A(_08889_),
    .X(_02275_));
 sky130_fd_sc_hd__and2_2 _25319_ (.A(_08880_),
    .B(\decode.regfile.registers_0[21] ),
    .X(_08890_));
 sky130_fd_sc_hd__buf_1 _25320_ (.A(_08890_),
    .X(_02276_));
 sky130_fd_sc_hd__buf_1 _25321_ (.A(_10018_),
    .X(_08891_));
 sky130_fd_sc_hd__and2_2 _25322_ (.A(_08891_),
    .B(\decode.regfile.registers_0[22] ),
    .X(_08892_));
 sky130_fd_sc_hd__buf_1 _25323_ (.A(_08892_),
    .X(_02277_));
 sky130_fd_sc_hd__and2_2 _25324_ (.A(_08891_),
    .B(\decode.regfile.registers_0[23] ),
    .X(_08893_));
 sky130_fd_sc_hd__buf_1 _25325_ (.A(_08893_),
    .X(_02278_));
 sky130_fd_sc_hd__and2_2 _25326_ (.A(_08891_),
    .B(\decode.regfile.registers_0[24] ),
    .X(_08894_));
 sky130_fd_sc_hd__buf_1 _25327_ (.A(_08894_),
    .X(_02279_));
 sky130_fd_sc_hd__and2_2 _25328_ (.A(_08891_),
    .B(\decode.regfile.registers_0[25] ),
    .X(_08895_));
 sky130_fd_sc_hd__buf_1 _25329_ (.A(_08895_),
    .X(_02280_));
 sky130_fd_sc_hd__and2_2 _25330_ (.A(_08891_),
    .B(\decode.regfile.registers_0[26] ),
    .X(_08896_));
 sky130_fd_sc_hd__buf_1 _25331_ (.A(_08896_),
    .X(_02281_));
 sky130_fd_sc_hd__and2_2 _25332_ (.A(_08891_),
    .B(\decode.regfile.registers_0[27] ),
    .X(_08897_));
 sky130_fd_sc_hd__buf_1 _25333_ (.A(_08897_),
    .X(_02282_));
 sky130_fd_sc_hd__and2_2 _25334_ (.A(_08891_),
    .B(\decode.regfile.registers_0[28] ),
    .X(_08898_));
 sky130_fd_sc_hd__buf_1 _25335_ (.A(_08898_),
    .X(_02283_));
 sky130_fd_sc_hd__and2_2 _25336_ (.A(_08891_),
    .B(\decode.regfile.registers_0[29] ),
    .X(_08899_));
 sky130_fd_sc_hd__buf_1 _25337_ (.A(_08899_),
    .X(_02284_));
 sky130_fd_sc_hd__and2_2 _25338_ (.A(_08891_),
    .B(\decode.regfile.registers_0[30] ),
    .X(_08900_));
 sky130_fd_sc_hd__buf_1 _25339_ (.A(_08900_),
    .X(_02285_));
 sky130_fd_sc_hd__and2_2 _25340_ (.A(_08891_),
    .B(\decode.regfile.registers_0[31] ),
    .X(_08901_));
 sky130_fd_sc_hd__buf_1 _25341_ (.A(_08901_),
    .X(_02286_));
 sky130_fd_sc_hd__and2b_2 _25342_ (.A_N(\decode.io_wb_rd[4] ),
    .B(\decode.io_wb_regwrite ),
    .X(_08902_));
 sky130_fd_sc_hd__buf_1 _25343_ (.A(_08902_),
    .X(_08903_));
 sky130_fd_sc_hd__and3_2 _25344_ (.A(_10240_),
    .B(_03672_),
    .C(_08903_),
    .X(_08904_));
 sky130_fd_sc_hd__buf_1 _25345_ (.A(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__buf_1 _25346_ (.A(_08905_),
    .X(_08906_));
 sky130_fd_sc_hd__buf_1 _25347_ (.A(_08905_),
    .X(_08907_));
 sky130_fd_sc_hd__nand2_2 _25348_ (.A(_09950_),
    .B(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__o211a_2 _25349_ (.A1(\decode.regfile.registers_1[0] ),
    .A2(_08906_),
    .B1(_08908_),
    .C1(_07247_),
    .X(_02287_));
 sky130_fd_sc_hd__nand2_2 _25350_ (.A(_09964_),
    .B(_08907_),
    .Y(_08909_));
 sky130_fd_sc_hd__o211a_2 _25351_ (.A1(\decode.regfile.registers_1[1] ),
    .A2(_08906_),
    .B1(_08909_),
    .C1(_07247_),
    .X(_02288_));
 sky130_fd_sc_hd__buf_1 _25352_ (.A(_09969_),
    .X(_08910_));
 sky130_fd_sc_hd__nand2_2 _25353_ (.A(_08910_),
    .B(_08907_),
    .Y(_08911_));
 sky130_fd_sc_hd__o211a_2 _25354_ (.A1(\decode.regfile.registers_1[2] ),
    .A2(_08906_),
    .B1(_08911_),
    .C1(_07247_),
    .X(_02289_));
 sky130_fd_sc_hd__buf_1 _25355_ (.A(_09974_),
    .X(_08912_));
 sky130_fd_sc_hd__nand2_2 _25356_ (.A(_08912_),
    .B(_08907_),
    .Y(_08913_));
 sky130_fd_sc_hd__o211a_2 _25357_ (.A1(\decode.regfile.registers_1[3] ),
    .A2(_08906_),
    .B1(_08913_),
    .C1(_07247_),
    .X(_02290_));
 sky130_fd_sc_hd__buf_1 _25358_ (.A(_09983_),
    .X(_08914_));
 sky130_fd_sc_hd__nand2_2 _25359_ (.A(_08914_),
    .B(_08907_),
    .Y(_08915_));
 sky130_fd_sc_hd__o211a_2 _25360_ (.A1(\decode.regfile.registers_1[4] ),
    .A2(_08906_),
    .B1(_08915_),
    .C1(_07247_),
    .X(_02291_));
 sky130_fd_sc_hd__buf_1 _25361_ (.A(_09992_),
    .X(_08916_));
 sky130_fd_sc_hd__nand2_2 _25362_ (.A(_08916_),
    .B(_08907_),
    .Y(_08917_));
 sky130_fd_sc_hd__o211a_2 _25363_ (.A1(\decode.regfile.registers_1[5] ),
    .A2(_08906_),
    .B1(_08917_),
    .C1(_07247_),
    .X(_02292_));
 sky130_fd_sc_hd__buf_1 _25364_ (.A(_09998_),
    .X(_08918_));
 sky130_fd_sc_hd__nand2_2 _25365_ (.A(_08918_),
    .B(_08907_),
    .Y(_08919_));
 sky130_fd_sc_hd__o211a_2 _25366_ (.A1(\decode.regfile.registers_1[6] ),
    .A2(_08906_),
    .B1(_08919_),
    .C1(_07247_),
    .X(_02293_));
 sky130_fd_sc_hd__buf_1 _25367_ (.A(_10007_),
    .X(_08920_));
 sky130_fd_sc_hd__nand2_2 _25368_ (.A(_08920_),
    .B(_08907_),
    .Y(_08921_));
 sky130_fd_sc_hd__o211a_2 _25369_ (.A1(\decode.regfile.registers_1[7] ),
    .A2(_08906_),
    .B1(_08921_),
    .C1(_07247_),
    .X(_02294_));
 sky130_fd_sc_hd__buf_1 _25370_ (.A(_10014_),
    .X(_08922_));
 sky130_fd_sc_hd__buf_1 _25371_ (.A(_08905_),
    .X(_08923_));
 sky130_fd_sc_hd__nand2_2 _25372_ (.A(_08922_),
    .B(_08923_),
    .Y(_08924_));
 sky130_fd_sc_hd__o211a_2 _25373_ (.A1(\decode.regfile.registers_1[8] ),
    .A2(_08906_),
    .B1(_08924_),
    .C1(_07247_),
    .X(_02295_));
 sky130_fd_sc_hd__buf_1 _25374_ (.A(_10024_),
    .X(_08925_));
 sky130_fd_sc_hd__nand2_2 _25375_ (.A(_08925_),
    .B(_08923_),
    .Y(_08926_));
 sky130_fd_sc_hd__buf_1 _25376_ (.A(_06578_),
    .X(_08927_));
 sky130_fd_sc_hd__o211a_2 _25377_ (.A1(\decode.regfile.registers_1[9] ),
    .A2(_08906_),
    .B1(_08926_),
    .C1(_08927_),
    .X(_02296_));
 sky130_fd_sc_hd__buf_1 _25378_ (.A(_08905_),
    .X(_08928_));
 sky130_fd_sc_hd__buf_1 _25379_ (.A(_10030_),
    .X(_08929_));
 sky130_fd_sc_hd__nand2_2 _25380_ (.A(_08929_),
    .B(_08923_),
    .Y(_08930_));
 sky130_fd_sc_hd__o211a_2 _25381_ (.A1(\decode.regfile.registers_1[10] ),
    .A2(_08928_),
    .B1(_08930_),
    .C1(_08927_),
    .X(_02297_));
 sky130_fd_sc_hd__buf_1 _25382_ (.A(_10035_),
    .X(_08931_));
 sky130_fd_sc_hd__nand2_2 _25383_ (.A(_08931_),
    .B(_08923_),
    .Y(_08932_));
 sky130_fd_sc_hd__o211a_2 _25384_ (.A1(\decode.regfile.registers_1[11] ),
    .A2(_08928_),
    .B1(_08932_),
    .C1(_08927_),
    .X(_02298_));
 sky130_fd_sc_hd__buf_1 _25385_ (.A(_10041_),
    .X(_08933_));
 sky130_fd_sc_hd__nand2_2 _25386_ (.A(_08933_),
    .B(_08923_),
    .Y(_08934_));
 sky130_fd_sc_hd__o211a_2 _25387_ (.A1(\decode.regfile.registers_1[12] ),
    .A2(_08928_),
    .B1(_08934_),
    .C1(_08927_),
    .X(_02299_));
 sky130_fd_sc_hd__buf_1 _25388_ (.A(_10047_),
    .X(_08935_));
 sky130_fd_sc_hd__nand2_2 _25389_ (.A(_08935_),
    .B(_08923_),
    .Y(_08936_));
 sky130_fd_sc_hd__o211a_2 _25390_ (.A1(\decode.regfile.registers_1[13] ),
    .A2(_08928_),
    .B1(_08936_),
    .C1(_08927_),
    .X(_02300_));
 sky130_fd_sc_hd__buf_1 _25391_ (.A(_10052_),
    .X(_08937_));
 sky130_fd_sc_hd__nand2_2 _25392_ (.A(_08937_),
    .B(_08923_),
    .Y(_08938_));
 sky130_fd_sc_hd__o211a_2 _25393_ (.A1(\decode.regfile.registers_1[14] ),
    .A2(_08928_),
    .B1(_08938_),
    .C1(_08927_),
    .X(_02301_));
 sky130_fd_sc_hd__buf_1 _25394_ (.A(_10057_),
    .X(_08939_));
 sky130_fd_sc_hd__nand2_2 _25395_ (.A(_08939_),
    .B(_08923_),
    .Y(_08940_));
 sky130_fd_sc_hd__o211a_2 _25396_ (.A1(\decode.regfile.registers_1[15] ),
    .A2(_08928_),
    .B1(_08940_),
    .C1(_08927_),
    .X(_02302_));
 sky130_fd_sc_hd__buf_1 _25397_ (.A(_10063_),
    .X(_08941_));
 sky130_fd_sc_hd__nand2_2 _25398_ (.A(_08941_),
    .B(_08923_),
    .Y(_08942_));
 sky130_fd_sc_hd__o211a_2 _25399_ (.A1(\decode.regfile.registers_1[16] ),
    .A2(_08928_),
    .B1(_08942_),
    .C1(_08927_),
    .X(_02303_));
 sky130_fd_sc_hd__buf_1 _25400_ (.A(_10068_),
    .X(_08943_));
 sky130_fd_sc_hd__nand2_2 _25401_ (.A(_08943_),
    .B(_08923_),
    .Y(_08944_));
 sky130_fd_sc_hd__o211a_2 _25402_ (.A1(\decode.regfile.registers_1[17] ),
    .A2(_08928_),
    .B1(_08944_),
    .C1(_08927_),
    .X(_02304_));
 sky130_fd_sc_hd__buf_1 _25403_ (.A(_10073_),
    .X(_08945_));
 sky130_fd_sc_hd__buf_1 _25404_ (.A(_08905_),
    .X(_08946_));
 sky130_fd_sc_hd__nand2_2 _25405_ (.A(_08945_),
    .B(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__o211a_2 _25406_ (.A1(\decode.regfile.registers_1[18] ),
    .A2(_08928_),
    .B1(_08947_),
    .C1(_08927_),
    .X(_02305_));
 sky130_fd_sc_hd__buf_1 _25407_ (.A(_10080_),
    .X(_08948_));
 sky130_fd_sc_hd__nand2_2 _25408_ (.A(_08948_),
    .B(_08946_),
    .Y(_08949_));
 sky130_fd_sc_hd__buf_1 _25409_ (.A(_06578_),
    .X(_08950_));
 sky130_fd_sc_hd__o211a_2 _25410_ (.A1(\decode.regfile.registers_1[19] ),
    .A2(_08928_),
    .B1(_08949_),
    .C1(_08950_),
    .X(_02306_));
 sky130_fd_sc_hd__buf_1 _25411_ (.A(_08905_),
    .X(_08951_));
 sky130_fd_sc_hd__buf_1 _25412_ (.A(_10086_),
    .X(_08952_));
 sky130_fd_sc_hd__nand2_2 _25413_ (.A(_08952_),
    .B(_08946_),
    .Y(_08953_));
 sky130_fd_sc_hd__o211a_2 _25414_ (.A1(\decode.regfile.registers_1[20] ),
    .A2(_08951_),
    .B1(_08953_),
    .C1(_08950_),
    .X(_02307_));
 sky130_fd_sc_hd__buf_1 _25415_ (.A(_10091_),
    .X(_08954_));
 sky130_fd_sc_hd__nand2_2 _25416_ (.A(_08954_),
    .B(_08946_),
    .Y(_08955_));
 sky130_fd_sc_hd__o211a_2 _25417_ (.A1(\decode.regfile.registers_1[21] ),
    .A2(_08951_),
    .B1(_08955_),
    .C1(_08950_),
    .X(_02308_));
 sky130_fd_sc_hd__buf_1 _25418_ (.A(_10096_),
    .X(_08956_));
 sky130_fd_sc_hd__nand2_2 _25419_ (.A(_08956_),
    .B(_08946_),
    .Y(_08957_));
 sky130_fd_sc_hd__o211a_2 _25420_ (.A1(\decode.regfile.registers_1[22] ),
    .A2(_08951_),
    .B1(_08957_),
    .C1(_08950_),
    .X(_02309_));
 sky130_fd_sc_hd__buf_1 _25421_ (.A(_10101_),
    .X(_08958_));
 sky130_fd_sc_hd__nand2_2 _25422_ (.A(_08958_),
    .B(_08946_),
    .Y(_08959_));
 sky130_fd_sc_hd__o211a_2 _25423_ (.A1(\decode.regfile.registers_1[23] ),
    .A2(_08951_),
    .B1(_08959_),
    .C1(_08950_),
    .X(_02310_));
 sky130_fd_sc_hd__buf_1 _25424_ (.A(_10106_),
    .X(_08960_));
 sky130_fd_sc_hd__nand2_2 _25425_ (.A(_08960_),
    .B(_08946_),
    .Y(_08961_));
 sky130_fd_sc_hd__o211a_2 _25426_ (.A1(\decode.regfile.registers_1[24] ),
    .A2(_08951_),
    .B1(_08961_),
    .C1(_08950_),
    .X(_02311_));
 sky130_fd_sc_hd__buf_1 _25427_ (.A(_10111_),
    .X(_08962_));
 sky130_fd_sc_hd__nand2_2 _25428_ (.A(_08962_),
    .B(_08946_),
    .Y(_08963_));
 sky130_fd_sc_hd__o211a_2 _25429_ (.A1(\decode.regfile.registers_1[25] ),
    .A2(_08951_),
    .B1(_08963_),
    .C1(_08950_),
    .X(_02312_));
 sky130_fd_sc_hd__buf_1 _25430_ (.A(_10116_),
    .X(_08964_));
 sky130_fd_sc_hd__nand2_2 _25431_ (.A(_08964_),
    .B(_08946_),
    .Y(_08965_));
 sky130_fd_sc_hd__o211a_2 _25432_ (.A1(\decode.regfile.registers_1[26] ),
    .A2(_08951_),
    .B1(_08965_),
    .C1(_08950_),
    .X(_02313_));
 sky130_fd_sc_hd__buf_1 _25433_ (.A(_10121_),
    .X(_08966_));
 sky130_fd_sc_hd__nand2_2 _25434_ (.A(_08966_),
    .B(_08946_),
    .Y(_08967_));
 sky130_fd_sc_hd__o211a_2 _25435_ (.A1(\decode.regfile.registers_1[27] ),
    .A2(_08951_),
    .B1(_08967_),
    .C1(_08950_),
    .X(_02314_));
 sky130_fd_sc_hd__buf_1 _25436_ (.A(_10127_),
    .X(_08968_));
 sky130_fd_sc_hd__nand2_2 _25437_ (.A(_08968_),
    .B(_08905_),
    .Y(_08969_));
 sky130_fd_sc_hd__o211a_2 _25438_ (.A1(\decode.regfile.registers_1[28] ),
    .A2(_08951_),
    .B1(_08969_),
    .C1(_08950_),
    .X(_02315_));
 sky130_fd_sc_hd__buf_1 _25439_ (.A(_10135_),
    .X(_08970_));
 sky130_fd_sc_hd__nand2_2 _25440_ (.A(_08970_),
    .B(_08905_),
    .Y(_08971_));
 sky130_fd_sc_hd__buf_1 _25441_ (.A(_06578_),
    .X(_08972_));
 sky130_fd_sc_hd__o211a_2 _25442_ (.A1(\decode.regfile.registers_1[29] ),
    .A2(_08951_),
    .B1(_08971_),
    .C1(_08972_),
    .X(_02316_));
 sky130_fd_sc_hd__buf_1 _25443_ (.A(_10141_),
    .X(_08973_));
 sky130_fd_sc_hd__nand2_2 _25444_ (.A(_08973_),
    .B(_08905_),
    .Y(_08974_));
 sky130_fd_sc_hd__o211a_2 _25445_ (.A1(\decode.regfile.registers_1[30] ),
    .A2(_08907_),
    .B1(_08974_),
    .C1(_08972_),
    .X(_02317_));
 sky130_fd_sc_hd__buf_1 _25446_ (.A(_10146_),
    .X(_08975_));
 sky130_fd_sc_hd__nand2_2 _25447_ (.A(_08975_),
    .B(_08905_),
    .Y(_08976_));
 sky130_fd_sc_hd__o211a_2 _25448_ (.A1(\decode.regfile.registers_1[31] ),
    .A2(_08907_),
    .B1(_08976_),
    .C1(_08972_),
    .X(_02318_));
 sky130_fd_sc_hd__and3_2 _25449_ (.A(_09932_),
    .B(_03672_),
    .C(_08903_),
    .X(_08977_));
 sky130_fd_sc_hd__buf_1 _25450_ (.A(_08977_),
    .X(_08978_));
 sky130_fd_sc_hd__buf_1 _25451_ (.A(_08978_),
    .X(_08979_));
 sky130_fd_sc_hd__buf_1 _25452_ (.A(_08978_),
    .X(_08980_));
 sky130_fd_sc_hd__nand2_2 _25453_ (.A(_09950_),
    .B(_08980_),
    .Y(_08981_));
 sky130_fd_sc_hd__o211a_2 _25454_ (.A1(\decode.regfile.registers_2[0] ),
    .A2(_08979_),
    .B1(_08981_),
    .C1(_08972_),
    .X(_02319_));
 sky130_fd_sc_hd__buf_1 _25455_ (.A(_09963_),
    .X(_08982_));
 sky130_fd_sc_hd__nand2_2 _25456_ (.A(_08982_),
    .B(_08980_),
    .Y(_08983_));
 sky130_fd_sc_hd__o211a_2 _25457_ (.A1(\decode.regfile.registers_2[1] ),
    .A2(_08979_),
    .B1(_08983_),
    .C1(_08972_),
    .X(_02320_));
 sky130_fd_sc_hd__nand2_2 _25458_ (.A(_08910_),
    .B(_08980_),
    .Y(_08984_));
 sky130_fd_sc_hd__o211a_2 _25459_ (.A1(\decode.regfile.registers_2[2] ),
    .A2(_08979_),
    .B1(_08984_),
    .C1(_08972_),
    .X(_02321_));
 sky130_fd_sc_hd__nand2_2 _25460_ (.A(_08912_),
    .B(_08980_),
    .Y(_08985_));
 sky130_fd_sc_hd__o211a_2 _25461_ (.A1(\decode.regfile.registers_2[3] ),
    .A2(_08979_),
    .B1(_08985_),
    .C1(_08972_),
    .X(_02322_));
 sky130_fd_sc_hd__nand2_2 _25462_ (.A(_08914_),
    .B(_08980_),
    .Y(_08986_));
 sky130_fd_sc_hd__o211a_2 _25463_ (.A1(\decode.regfile.registers_2[4] ),
    .A2(_08979_),
    .B1(_08986_),
    .C1(_08972_),
    .X(_02323_));
 sky130_fd_sc_hd__nand2_2 _25464_ (.A(_08916_),
    .B(_08980_),
    .Y(_08987_));
 sky130_fd_sc_hd__o211a_2 _25465_ (.A1(\decode.regfile.registers_2[5] ),
    .A2(_08979_),
    .B1(_08987_),
    .C1(_08972_),
    .X(_02324_));
 sky130_fd_sc_hd__nand2_2 _25466_ (.A(_08918_),
    .B(_08980_),
    .Y(_08988_));
 sky130_fd_sc_hd__o211a_2 _25467_ (.A1(\decode.regfile.registers_2[6] ),
    .A2(_08979_),
    .B1(_08988_),
    .C1(_08972_),
    .X(_02325_));
 sky130_fd_sc_hd__nand2_2 _25468_ (.A(_08920_),
    .B(_08980_),
    .Y(_08989_));
 sky130_fd_sc_hd__buf_1 _25469_ (.A(_10130_),
    .X(_08990_));
 sky130_fd_sc_hd__buf_1 _25470_ (.A(_08990_),
    .X(_08991_));
 sky130_fd_sc_hd__o211a_2 _25471_ (.A1(\decode.regfile.registers_2[7] ),
    .A2(_08979_),
    .B1(_08989_),
    .C1(_08991_),
    .X(_02326_));
 sky130_fd_sc_hd__buf_1 _25472_ (.A(_08978_),
    .X(_08992_));
 sky130_fd_sc_hd__nand2_2 _25473_ (.A(_08922_),
    .B(_08992_),
    .Y(_08993_));
 sky130_fd_sc_hd__o211a_2 _25474_ (.A1(\decode.regfile.registers_2[8] ),
    .A2(_08979_),
    .B1(_08993_),
    .C1(_08991_),
    .X(_02327_));
 sky130_fd_sc_hd__nand2_2 _25475_ (.A(_08925_),
    .B(_08992_),
    .Y(_08994_));
 sky130_fd_sc_hd__o211a_2 _25476_ (.A1(\decode.regfile.registers_2[9] ),
    .A2(_08979_),
    .B1(_08994_),
    .C1(_08991_),
    .X(_02328_));
 sky130_fd_sc_hd__buf_1 _25477_ (.A(_08978_),
    .X(_08995_));
 sky130_fd_sc_hd__nand2_2 _25478_ (.A(_08929_),
    .B(_08992_),
    .Y(_08996_));
 sky130_fd_sc_hd__o211a_2 _25479_ (.A1(\decode.regfile.registers_2[10] ),
    .A2(_08995_),
    .B1(_08996_),
    .C1(_08991_),
    .X(_02329_));
 sky130_fd_sc_hd__nand2_2 _25480_ (.A(_08931_),
    .B(_08992_),
    .Y(_08997_));
 sky130_fd_sc_hd__o211a_2 _25481_ (.A1(\decode.regfile.registers_2[11] ),
    .A2(_08995_),
    .B1(_08997_),
    .C1(_08991_),
    .X(_02330_));
 sky130_fd_sc_hd__nand2_2 _25482_ (.A(_08933_),
    .B(_08992_),
    .Y(_08998_));
 sky130_fd_sc_hd__o211a_2 _25483_ (.A1(\decode.regfile.registers_2[12] ),
    .A2(_08995_),
    .B1(_08998_),
    .C1(_08991_),
    .X(_02331_));
 sky130_fd_sc_hd__nand2_2 _25484_ (.A(_08935_),
    .B(_08992_),
    .Y(_08999_));
 sky130_fd_sc_hd__o211a_2 _25485_ (.A1(\decode.regfile.registers_2[13] ),
    .A2(_08995_),
    .B1(_08999_),
    .C1(_08991_),
    .X(_02332_));
 sky130_fd_sc_hd__nand2_2 _25486_ (.A(_08937_),
    .B(_08992_),
    .Y(_09000_));
 sky130_fd_sc_hd__o211a_2 _25487_ (.A1(\decode.regfile.registers_2[14] ),
    .A2(_08995_),
    .B1(_09000_),
    .C1(_08991_),
    .X(_02333_));
 sky130_fd_sc_hd__nand2_2 _25488_ (.A(_08939_),
    .B(_08992_),
    .Y(_09001_));
 sky130_fd_sc_hd__o211a_2 _25489_ (.A1(\decode.regfile.registers_2[15] ),
    .A2(_08995_),
    .B1(_09001_),
    .C1(_08991_),
    .X(_02334_));
 sky130_fd_sc_hd__nand2_2 _25490_ (.A(_08941_),
    .B(_08992_),
    .Y(_09002_));
 sky130_fd_sc_hd__o211a_2 _25491_ (.A1(\decode.regfile.registers_2[16] ),
    .A2(_08995_),
    .B1(_09002_),
    .C1(_08991_),
    .X(_02335_));
 sky130_fd_sc_hd__nand2_2 _25492_ (.A(_08943_),
    .B(_08992_),
    .Y(_09003_));
 sky130_fd_sc_hd__buf_1 _25493_ (.A(_08990_),
    .X(_09004_));
 sky130_fd_sc_hd__o211a_2 _25494_ (.A1(\decode.regfile.registers_2[17] ),
    .A2(_08995_),
    .B1(_09003_),
    .C1(_09004_),
    .X(_02336_));
 sky130_fd_sc_hd__buf_1 _25495_ (.A(_08978_),
    .X(_09005_));
 sky130_fd_sc_hd__nand2_2 _25496_ (.A(_08945_),
    .B(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__o211a_2 _25497_ (.A1(\decode.regfile.registers_2[18] ),
    .A2(_08995_),
    .B1(_09006_),
    .C1(_09004_),
    .X(_02337_));
 sky130_fd_sc_hd__nand2_2 _25498_ (.A(_08948_),
    .B(_09005_),
    .Y(_09007_));
 sky130_fd_sc_hd__o211a_2 _25499_ (.A1(\decode.regfile.registers_2[19] ),
    .A2(_08995_),
    .B1(_09007_),
    .C1(_09004_),
    .X(_02338_));
 sky130_fd_sc_hd__buf_1 _25500_ (.A(_08978_),
    .X(_09008_));
 sky130_fd_sc_hd__nand2_2 _25501_ (.A(_08952_),
    .B(_09005_),
    .Y(_09009_));
 sky130_fd_sc_hd__o211a_2 _25502_ (.A1(\decode.regfile.registers_2[20] ),
    .A2(_09008_),
    .B1(_09009_),
    .C1(_09004_),
    .X(_02339_));
 sky130_fd_sc_hd__nand2_2 _25503_ (.A(_08954_),
    .B(_09005_),
    .Y(_09010_));
 sky130_fd_sc_hd__o211a_2 _25504_ (.A1(\decode.regfile.registers_2[21] ),
    .A2(_09008_),
    .B1(_09010_),
    .C1(_09004_),
    .X(_02340_));
 sky130_fd_sc_hd__nand2_2 _25505_ (.A(_08956_),
    .B(_09005_),
    .Y(_09011_));
 sky130_fd_sc_hd__o211a_2 _25506_ (.A1(\decode.regfile.registers_2[22] ),
    .A2(_09008_),
    .B1(_09011_),
    .C1(_09004_),
    .X(_02341_));
 sky130_fd_sc_hd__nand2_2 _25507_ (.A(_08958_),
    .B(_09005_),
    .Y(_09012_));
 sky130_fd_sc_hd__o211a_2 _25508_ (.A1(\decode.regfile.registers_2[23] ),
    .A2(_09008_),
    .B1(_09012_),
    .C1(_09004_),
    .X(_02342_));
 sky130_fd_sc_hd__nand2_2 _25509_ (.A(_08960_),
    .B(_09005_),
    .Y(_09013_));
 sky130_fd_sc_hd__o211a_2 _25510_ (.A1(\decode.regfile.registers_2[24] ),
    .A2(_09008_),
    .B1(_09013_),
    .C1(_09004_),
    .X(_02343_));
 sky130_fd_sc_hd__nand2_2 _25511_ (.A(_08962_),
    .B(_09005_),
    .Y(_09014_));
 sky130_fd_sc_hd__o211a_2 _25512_ (.A1(\decode.regfile.registers_2[25] ),
    .A2(_09008_),
    .B1(_09014_),
    .C1(_09004_),
    .X(_02344_));
 sky130_fd_sc_hd__nand2_2 _25513_ (.A(_08964_),
    .B(_09005_),
    .Y(_09015_));
 sky130_fd_sc_hd__o211a_2 _25514_ (.A1(\decode.regfile.registers_2[26] ),
    .A2(_09008_),
    .B1(_09015_),
    .C1(_09004_),
    .X(_02345_));
 sky130_fd_sc_hd__nand2_2 _25515_ (.A(_08966_),
    .B(_09005_),
    .Y(_09016_));
 sky130_fd_sc_hd__buf_1 _25516_ (.A(_08990_),
    .X(_09017_));
 sky130_fd_sc_hd__o211a_2 _25517_ (.A1(\decode.regfile.registers_2[27] ),
    .A2(_09008_),
    .B1(_09016_),
    .C1(_09017_),
    .X(_02346_));
 sky130_fd_sc_hd__nand2_2 _25518_ (.A(_08968_),
    .B(_08978_),
    .Y(_09018_));
 sky130_fd_sc_hd__o211a_2 _25519_ (.A1(\decode.regfile.registers_2[28] ),
    .A2(_09008_),
    .B1(_09018_),
    .C1(_09017_),
    .X(_02347_));
 sky130_fd_sc_hd__nand2_2 _25520_ (.A(_08970_),
    .B(_08978_),
    .Y(_09019_));
 sky130_fd_sc_hd__o211a_2 _25521_ (.A1(\decode.regfile.registers_2[29] ),
    .A2(_09008_),
    .B1(_09019_),
    .C1(_09017_),
    .X(_02348_));
 sky130_fd_sc_hd__nand2_2 _25522_ (.A(_08973_),
    .B(_08978_),
    .Y(_09020_));
 sky130_fd_sc_hd__o211a_2 _25523_ (.A1(\decode.regfile.registers_2[30] ),
    .A2(_08980_),
    .B1(_09020_),
    .C1(_09017_),
    .X(_02349_));
 sky130_fd_sc_hd__nand2_2 _25524_ (.A(_08975_),
    .B(_08978_),
    .Y(_09021_));
 sky130_fd_sc_hd__o211a_2 _25525_ (.A1(\decode.regfile.registers_2[31] ),
    .A2(_08980_),
    .B1(_09021_),
    .C1(_09017_),
    .X(_02350_));
 sky130_fd_sc_hd__and3_2 _25526_ (.A(_10150_),
    .B(_03672_),
    .C(_08903_),
    .X(_09022_));
 sky130_fd_sc_hd__buf_1 _25527_ (.A(_09022_),
    .X(_09023_));
 sky130_fd_sc_hd__buf_1 _25528_ (.A(_09023_),
    .X(_09024_));
 sky130_fd_sc_hd__buf_1 _25529_ (.A(_09949_),
    .X(_09025_));
 sky130_fd_sc_hd__buf_1 _25530_ (.A(_09023_),
    .X(_09026_));
 sky130_fd_sc_hd__nand2_2 _25531_ (.A(_09025_),
    .B(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__o211a_2 _25532_ (.A1(\decode.regfile.registers_3[0] ),
    .A2(_09024_),
    .B1(_09027_),
    .C1(_09017_),
    .X(_02351_));
 sky130_fd_sc_hd__nand2_2 _25533_ (.A(_08982_),
    .B(_09026_),
    .Y(_09028_));
 sky130_fd_sc_hd__o211a_2 _25534_ (.A1(\decode.regfile.registers_3[1] ),
    .A2(_09024_),
    .B1(_09028_),
    .C1(_09017_),
    .X(_02352_));
 sky130_fd_sc_hd__nand2_2 _25535_ (.A(_08910_),
    .B(_09026_),
    .Y(_09029_));
 sky130_fd_sc_hd__o211a_2 _25536_ (.A1(\decode.regfile.registers_3[2] ),
    .A2(_09024_),
    .B1(_09029_),
    .C1(_09017_),
    .X(_02353_));
 sky130_fd_sc_hd__nand2_2 _25537_ (.A(_08912_),
    .B(_09026_),
    .Y(_09030_));
 sky130_fd_sc_hd__o211a_2 _25538_ (.A1(\decode.regfile.registers_3[3] ),
    .A2(_09024_),
    .B1(_09030_),
    .C1(_09017_),
    .X(_02354_));
 sky130_fd_sc_hd__nand2_2 _25539_ (.A(_08914_),
    .B(_09026_),
    .Y(_09031_));
 sky130_fd_sc_hd__o211a_2 _25540_ (.A1(\decode.regfile.registers_3[4] ),
    .A2(_09024_),
    .B1(_09031_),
    .C1(_09017_),
    .X(_02355_));
 sky130_fd_sc_hd__nand2_2 _25541_ (.A(_08916_),
    .B(_09026_),
    .Y(_09032_));
 sky130_fd_sc_hd__buf_1 _25542_ (.A(_08990_),
    .X(_09033_));
 sky130_fd_sc_hd__o211a_2 _25543_ (.A1(\decode.regfile.registers_3[5] ),
    .A2(_09024_),
    .B1(_09032_),
    .C1(_09033_),
    .X(_02356_));
 sky130_fd_sc_hd__nand2_2 _25544_ (.A(_08918_),
    .B(_09026_),
    .Y(_09034_));
 sky130_fd_sc_hd__o211a_2 _25545_ (.A1(\decode.regfile.registers_3[6] ),
    .A2(_09024_),
    .B1(_09034_),
    .C1(_09033_),
    .X(_02357_));
 sky130_fd_sc_hd__nand2_2 _25546_ (.A(_08920_),
    .B(_09026_),
    .Y(_09035_));
 sky130_fd_sc_hd__o211a_2 _25547_ (.A1(\decode.regfile.registers_3[7] ),
    .A2(_09024_),
    .B1(_09035_),
    .C1(_09033_),
    .X(_02358_));
 sky130_fd_sc_hd__buf_1 _25548_ (.A(_09023_),
    .X(_09036_));
 sky130_fd_sc_hd__nand2_2 _25549_ (.A(_08922_),
    .B(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__o211a_2 _25550_ (.A1(\decode.regfile.registers_3[8] ),
    .A2(_09024_),
    .B1(_09037_),
    .C1(_09033_),
    .X(_02359_));
 sky130_fd_sc_hd__nand2_2 _25551_ (.A(_08925_),
    .B(_09036_),
    .Y(_09038_));
 sky130_fd_sc_hd__o211a_2 _25552_ (.A1(\decode.regfile.registers_3[9] ),
    .A2(_09024_),
    .B1(_09038_),
    .C1(_09033_),
    .X(_02360_));
 sky130_fd_sc_hd__buf_1 _25553_ (.A(_09023_),
    .X(_09039_));
 sky130_fd_sc_hd__nand2_2 _25554_ (.A(_08929_),
    .B(_09036_),
    .Y(_09040_));
 sky130_fd_sc_hd__o211a_2 _25555_ (.A1(\decode.regfile.registers_3[10] ),
    .A2(_09039_),
    .B1(_09040_),
    .C1(_09033_),
    .X(_02361_));
 sky130_fd_sc_hd__nand2_2 _25556_ (.A(_08931_),
    .B(_09036_),
    .Y(_09041_));
 sky130_fd_sc_hd__o211a_2 _25557_ (.A1(\decode.regfile.registers_3[11] ),
    .A2(_09039_),
    .B1(_09041_),
    .C1(_09033_),
    .X(_02362_));
 sky130_fd_sc_hd__nand2_2 _25558_ (.A(_08933_),
    .B(_09036_),
    .Y(_09042_));
 sky130_fd_sc_hd__o211a_2 _25559_ (.A1(\decode.regfile.registers_3[12] ),
    .A2(_09039_),
    .B1(_09042_),
    .C1(_09033_),
    .X(_02363_));
 sky130_fd_sc_hd__nand2_2 _25560_ (.A(_08935_),
    .B(_09036_),
    .Y(_09043_));
 sky130_fd_sc_hd__o211a_2 _25561_ (.A1(\decode.regfile.registers_3[13] ),
    .A2(_09039_),
    .B1(_09043_),
    .C1(_09033_),
    .X(_02364_));
 sky130_fd_sc_hd__nand2_2 _25562_ (.A(_08937_),
    .B(_09036_),
    .Y(_09044_));
 sky130_fd_sc_hd__o211a_2 _25563_ (.A1(\decode.regfile.registers_3[14] ),
    .A2(_09039_),
    .B1(_09044_),
    .C1(_09033_),
    .X(_02365_));
 sky130_fd_sc_hd__nand2_2 _25564_ (.A(_08939_),
    .B(_09036_),
    .Y(_09045_));
 sky130_fd_sc_hd__buf_1 _25565_ (.A(_08990_),
    .X(_09046_));
 sky130_fd_sc_hd__o211a_2 _25566_ (.A1(\decode.regfile.registers_3[15] ),
    .A2(_09039_),
    .B1(_09045_),
    .C1(_09046_),
    .X(_02366_));
 sky130_fd_sc_hd__nand2_2 _25567_ (.A(_08941_),
    .B(_09036_),
    .Y(_09047_));
 sky130_fd_sc_hd__o211a_2 _25568_ (.A1(\decode.regfile.registers_3[16] ),
    .A2(_09039_),
    .B1(_09047_),
    .C1(_09046_),
    .X(_02367_));
 sky130_fd_sc_hd__nand2_2 _25569_ (.A(_08943_),
    .B(_09036_),
    .Y(_09048_));
 sky130_fd_sc_hd__o211a_2 _25570_ (.A1(\decode.regfile.registers_3[17] ),
    .A2(_09039_),
    .B1(_09048_),
    .C1(_09046_),
    .X(_02368_));
 sky130_fd_sc_hd__buf_1 _25571_ (.A(_09023_),
    .X(_09049_));
 sky130_fd_sc_hd__nand2_2 _25572_ (.A(_08945_),
    .B(_09049_),
    .Y(_09050_));
 sky130_fd_sc_hd__o211a_2 _25573_ (.A1(\decode.regfile.registers_3[18] ),
    .A2(_09039_),
    .B1(_09050_),
    .C1(_09046_),
    .X(_02369_));
 sky130_fd_sc_hd__nand2_2 _25574_ (.A(_08948_),
    .B(_09049_),
    .Y(_09051_));
 sky130_fd_sc_hd__o211a_2 _25575_ (.A1(\decode.regfile.registers_3[19] ),
    .A2(_09039_),
    .B1(_09051_),
    .C1(_09046_),
    .X(_02370_));
 sky130_fd_sc_hd__buf_1 _25576_ (.A(_09023_),
    .X(_09052_));
 sky130_fd_sc_hd__nand2_2 _25577_ (.A(_08952_),
    .B(_09049_),
    .Y(_09053_));
 sky130_fd_sc_hd__o211a_2 _25578_ (.A1(\decode.regfile.registers_3[20] ),
    .A2(_09052_),
    .B1(_09053_),
    .C1(_09046_),
    .X(_02371_));
 sky130_fd_sc_hd__nand2_2 _25579_ (.A(_08954_),
    .B(_09049_),
    .Y(_09054_));
 sky130_fd_sc_hd__o211a_2 _25580_ (.A1(\decode.regfile.registers_3[21] ),
    .A2(_09052_),
    .B1(_09054_),
    .C1(_09046_),
    .X(_02372_));
 sky130_fd_sc_hd__nand2_2 _25581_ (.A(_08956_),
    .B(_09049_),
    .Y(_09055_));
 sky130_fd_sc_hd__o211a_2 _25582_ (.A1(\decode.regfile.registers_3[22] ),
    .A2(_09052_),
    .B1(_09055_),
    .C1(_09046_),
    .X(_02373_));
 sky130_fd_sc_hd__nand2_2 _25583_ (.A(_08958_),
    .B(_09049_),
    .Y(_09056_));
 sky130_fd_sc_hd__o211a_2 _25584_ (.A1(\decode.regfile.registers_3[23] ),
    .A2(_09052_),
    .B1(_09056_),
    .C1(_09046_),
    .X(_02374_));
 sky130_fd_sc_hd__nand2_2 _25585_ (.A(_08960_),
    .B(_09049_),
    .Y(_09057_));
 sky130_fd_sc_hd__o211a_2 _25586_ (.A1(\decode.regfile.registers_3[24] ),
    .A2(_09052_),
    .B1(_09057_),
    .C1(_09046_),
    .X(_02375_));
 sky130_fd_sc_hd__nand2_2 _25587_ (.A(_08962_),
    .B(_09049_),
    .Y(_09058_));
 sky130_fd_sc_hd__buf_1 _25588_ (.A(_08990_),
    .X(_09059_));
 sky130_fd_sc_hd__o211a_2 _25589_ (.A1(\decode.regfile.registers_3[25] ),
    .A2(_09052_),
    .B1(_09058_),
    .C1(_09059_),
    .X(_02376_));
 sky130_fd_sc_hd__nand2_2 _25590_ (.A(_08964_),
    .B(_09049_),
    .Y(_09060_));
 sky130_fd_sc_hd__o211a_2 _25591_ (.A1(\decode.regfile.registers_3[26] ),
    .A2(_09052_),
    .B1(_09060_),
    .C1(_09059_),
    .X(_02377_));
 sky130_fd_sc_hd__nand2_2 _25592_ (.A(_08966_),
    .B(_09049_),
    .Y(_09061_));
 sky130_fd_sc_hd__o211a_2 _25593_ (.A1(\decode.regfile.registers_3[27] ),
    .A2(_09052_),
    .B1(_09061_),
    .C1(_09059_),
    .X(_02378_));
 sky130_fd_sc_hd__nand2_2 _25594_ (.A(_08968_),
    .B(_09023_),
    .Y(_09062_));
 sky130_fd_sc_hd__o211a_2 _25595_ (.A1(\decode.regfile.registers_3[28] ),
    .A2(_09052_),
    .B1(_09062_),
    .C1(_09059_),
    .X(_02379_));
 sky130_fd_sc_hd__nand2_2 _25596_ (.A(_08970_),
    .B(_09023_),
    .Y(_09063_));
 sky130_fd_sc_hd__o211a_2 _25597_ (.A1(\decode.regfile.registers_3[29] ),
    .A2(_09052_),
    .B1(_09063_),
    .C1(_09059_),
    .X(_02380_));
 sky130_fd_sc_hd__nand2_2 _25598_ (.A(_08973_),
    .B(_09023_),
    .Y(_09064_));
 sky130_fd_sc_hd__o211a_2 _25599_ (.A1(\decode.regfile.registers_3[30] ),
    .A2(_09026_),
    .B1(_09064_),
    .C1(_09059_),
    .X(_02381_));
 sky130_fd_sc_hd__nand2_2 _25600_ (.A(_08975_),
    .B(_09023_),
    .Y(_09065_));
 sky130_fd_sc_hd__o211a_2 _25601_ (.A1(\decode.regfile.registers_3[31] ),
    .A2(_09026_),
    .B1(_09065_),
    .C1(_09059_),
    .X(_02382_));
 sky130_fd_sc_hd__and4_2 _25602_ (.A(_10373_),
    .B(_08903_),
    .C(_09935_),
    .D(_10196_),
    .X(_09066_));
 sky130_fd_sc_hd__buf_1 _25603_ (.A(_09066_),
    .X(_09067_));
 sky130_fd_sc_hd__buf_1 _25604_ (.A(_09067_),
    .X(_09068_));
 sky130_fd_sc_hd__buf_1 _25605_ (.A(_09067_),
    .X(_09069_));
 sky130_fd_sc_hd__nand2_2 _25606_ (.A(_09025_),
    .B(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__o211a_2 _25607_ (.A1(\decode.regfile.registers_4[0] ),
    .A2(_09068_),
    .B1(_09070_),
    .C1(_09059_),
    .X(_02383_));
 sky130_fd_sc_hd__nand2_2 _25608_ (.A(_08982_),
    .B(_09069_),
    .Y(_09071_));
 sky130_fd_sc_hd__o211a_2 _25609_ (.A1(\decode.regfile.registers_4[1] ),
    .A2(_09068_),
    .B1(_09071_),
    .C1(_09059_),
    .X(_02384_));
 sky130_fd_sc_hd__nand2_2 _25610_ (.A(_08910_),
    .B(_09069_),
    .Y(_09072_));
 sky130_fd_sc_hd__o211a_2 _25611_ (.A1(\decode.regfile.registers_4[2] ),
    .A2(_09068_),
    .B1(_09072_),
    .C1(_09059_),
    .X(_02385_));
 sky130_fd_sc_hd__nand2_2 _25612_ (.A(_08912_),
    .B(_09069_),
    .Y(_09073_));
 sky130_fd_sc_hd__buf_1 _25613_ (.A(_08990_),
    .X(_09074_));
 sky130_fd_sc_hd__o211a_2 _25614_ (.A1(\decode.regfile.registers_4[3] ),
    .A2(_09068_),
    .B1(_09073_),
    .C1(_09074_),
    .X(_02386_));
 sky130_fd_sc_hd__nand2_2 _25615_ (.A(_08914_),
    .B(_09069_),
    .Y(_09075_));
 sky130_fd_sc_hd__o211a_2 _25616_ (.A1(\decode.regfile.registers_4[4] ),
    .A2(_09068_),
    .B1(_09075_),
    .C1(_09074_),
    .X(_02387_));
 sky130_fd_sc_hd__nand2_2 _25617_ (.A(_08916_),
    .B(_09069_),
    .Y(_09076_));
 sky130_fd_sc_hd__o211a_2 _25618_ (.A1(\decode.regfile.registers_4[5] ),
    .A2(_09068_),
    .B1(_09076_),
    .C1(_09074_),
    .X(_02388_));
 sky130_fd_sc_hd__nand2_2 _25619_ (.A(_08918_),
    .B(_09069_),
    .Y(_09077_));
 sky130_fd_sc_hd__o211a_2 _25620_ (.A1(\decode.regfile.registers_4[6] ),
    .A2(_09068_),
    .B1(_09077_),
    .C1(_09074_),
    .X(_02389_));
 sky130_fd_sc_hd__nand2_2 _25621_ (.A(_08920_),
    .B(_09069_),
    .Y(_09078_));
 sky130_fd_sc_hd__o211a_2 _25622_ (.A1(\decode.regfile.registers_4[7] ),
    .A2(_09068_),
    .B1(_09078_),
    .C1(_09074_),
    .X(_02390_));
 sky130_fd_sc_hd__buf_1 _25623_ (.A(_09067_),
    .X(_09079_));
 sky130_fd_sc_hd__nand2_2 _25624_ (.A(_08922_),
    .B(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__o211a_2 _25625_ (.A1(\decode.regfile.registers_4[8] ),
    .A2(_09068_),
    .B1(_09080_),
    .C1(_09074_),
    .X(_02391_));
 sky130_fd_sc_hd__nand2_2 _25626_ (.A(_08925_),
    .B(_09079_),
    .Y(_09081_));
 sky130_fd_sc_hd__o211a_2 _25627_ (.A1(\decode.regfile.registers_4[9] ),
    .A2(_09068_),
    .B1(_09081_),
    .C1(_09074_),
    .X(_02392_));
 sky130_fd_sc_hd__buf_1 _25628_ (.A(_09067_),
    .X(_09082_));
 sky130_fd_sc_hd__nand2_2 _25629_ (.A(_08929_),
    .B(_09079_),
    .Y(_09083_));
 sky130_fd_sc_hd__o211a_2 _25630_ (.A1(\decode.regfile.registers_4[10] ),
    .A2(_09082_),
    .B1(_09083_),
    .C1(_09074_),
    .X(_02393_));
 sky130_fd_sc_hd__nand2_2 _25631_ (.A(_08931_),
    .B(_09079_),
    .Y(_09084_));
 sky130_fd_sc_hd__o211a_2 _25632_ (.A1(\decode.regfile.registers_4[11] ),
    .A2(_09082_),
    .B1(_09084_),
    .C1(_09074_),
    .X(_02394_));
 sky130_fd_sc_hd__nand2_2 _25633_ (.A(_08933_),
    .B(_09079_),
    .Y(_09085_));
 sky130_fd_sc_hd__o211a_2 _25634_ (.A1(\decode.regfile.registers_4[12] ),
    .A2(_09082_),
    .B1(_09085_),
    .C1(_09074_),
    .X(_02395_));
 sky130_fd_sc_hd__nand2_2 _25635_ (.A(_08935_),
    .B(_09079_),
    .Y(_09086_));
 sky130_fd_sc_hd__buf_1 _25636_ (.A(_08990_),
    .X(_09087_));
 sky130_fd_sc_hd__o211a_2 _25637_ (.A1(\decode.regfile.registers_4[13] ),
    .A2(_09082_),
    .B1(_09086_),
    .C1(_09087_),
    .X(_02396_));
 sky130_fd_sc_hd__nand2_2 _25638_ (.A(_08937_),
    .B(_09079_),
    .Y(_09088_));
 sky130_fd_sc_hd__o211a_2 _25639_ (.A1(\decode.regfile.registers_4[14] ),
    .A2(_09082_),
    .B1(_09088_),
    .C1(_09087_),
    .X(_02397_));
 sky130_fd_sc_hd__nand2_2 _25640_ (.A(_08939_),
    .B(_09079_),
    .Y(_09089_));
 sky130_fd_sc_hd__o211a_2 _25641_ (.A1(\decode.regfile.registers_4[15] ),
    .A2(_09082_),
    .B1(_09089_),
    .C1(_09087_),
    .X(_02398_));
 sky130_fd_sc_hd__nand2_2 _25642_ (.A(_08941_),
    .B(_09079_),
    .Y(_09090_));
 sky130_fd_sc_hd__o211a_2 _25643_ (.A1(\decode.regfile.registers_4[16] ),
    .A2(_09082_),
    .B1(_09090_),
    .C1(_09087_),
    .X(_02399_));
 sky130_fd_sc_hd__nand2_2 _25644_ (.A(_08943_),
    .B(_09079_),
    .Y(_09091_));
 sky130_fd_sc_hd__o211a_2 _25645_ (.A1(\decode.regfile.registers_4[17] ),
    .A2(_09082_),
    .B1(_09091_),
    .C1(_09087_),
    .X(_02400_));
 sky130_fd_sc_hd__buf_1 _25646_ (.A(_09067_),
    .X(_09092_));
 sky130_fd_sc_hd__nand2_2 _25647_ (.A(_08945_),
    .B(_09092_),
    .Y(_09093_));
 sky130_fd_sc_hd__o211a_2 _25648_ (.A1(\decode.regfile.registers_4[18] ),
    .A2(_09082_),
    .B1(_09093_),
    .C1(_09087_),
    .X(_02401_));
 sky130_fd_sc_hd__nand2_2 _25649_ (.A(_08948_),
    .B(_09092_),
    .Y(_09094_));
 sky130_fd_sc_hd__o211a_2 _25650_ (.A1(\decode.regfile.registers_4[19] ),
    .A2(_09082_),
    .B1(_09094_),
    .C1(_09087_),
    .X(_02402_));
 sky130_fd_sc_hd__buf_1 _25651_ (.A(_09067_),
    .X(_09095_));
 sky130_fd_sc_hd__nand2_2 _25652_ (.A(_08952_),
    .B(_09092_),
    .Y(_09096_));
 sky130_fd_sc_hd__o211a_2 _25653_ (.A1(\decode.regfile.registers_4[20] ),
    .A2(_09095_),
    .B1(_09096_),
    .C1(_09087_),
    .X(_02403_));
 sky130_fd_sc_hd__nand2_2 _25654_ (.A(_08954_),
    .B(_09092_),
    .Y(_09097_));
 sky130_fd_sc_hd__o211a_2 _25655_ (.A1(\decode.regfile.registers_4[21] ),
    .A2(_09095_),
    .B1(_09097_),
    .C1(_09087_),
    .X(_02404_));
 sky130_fd_sc_hd__nand2_2 _25656_ (.A(_08956_),
    .B(_09092_),
    .Y(_09098_));
 sky130_fd_sc_hd__o211a_2 _25657_ (.A1(\decode.regfile.registers_4[22] ),
    .A2(_09095_),
    .B1(_09098_),
    .C1(_09087_),
    .X(_02405_));
 sky130_fd_sc_hd__nand2_2 _25658_ (.A(_08958_),
    .B(_09092_),
    .Y(_09099_));
 sky130_fd_sc_hd__buf_1 _25659_ (.A(_08990_),
    .X(_09100_));
 sky130_fd_sc_hd__o211a_2 _25660_ (.A1(\decode.regfile.registers_4[23] ),
    .A2(_09095_),
    .B1(_09099_),
    .C1(_09100_),
    .X(_02406_));
 sky130_fd_sc_hd__nand2_2 _25661_ (.A(_08960_),
    .B(_09092_),
    .Y(_09101_));
 sky130_fd_sc_hd__o211a_2 _25662_ (.A1(\decode.regfile.registers_4[24] ),
    .A2(_09095_),
    .B1(_09101_),
    .C1(_09100_),
    .X(_02407_));
 sky130_fd_sc_hd__nand2_2 _25663_ (.A(_08962_),
    .B(_09092_),
    .Y(_09102_));
 sky130_fd_sc_hd__o211a_2 _25664_ (.A1(\decode.regfile.registers_4[25] ),
    .A2(_09095_),
    .B1(_09102_),
    .C1(_09100_),
    .X(_02408_));
 sky130_fd_sc_hd__nand2_2 _25665_ (.A(_08964_),
    .B(_09092_),
    .Y(_09103_));
 sky130_fd_sc_hd__o211a_2 _25666_ (.A1(\decode.regfile.registers_4[26] ),
    .A2(_09095_),
    .B1(_09103_),
    .C1(_09100_),
    .X(_02409_));
 sky130_fd_sc_hd__nand2_2 _25667_ (.A(_08966_),
    .B(_09092_),
    .Y(_09104_));
 sky130_fd_sc_hd__o211a_2 _25668_ (.A1(\decode.regfile.registers_4[27] ),
    .A2(_09095_),
    .B1(_09104_),
    .C1(_09100_),
    .X(_02410_));
 sky130_fd_sc_hd__nand2_2 _25669_ (.A(_08968_),
    .B(_09067_),
    .Y(_09105_));
 sky130_fd_sc_hd__o211a_2 _25670_ (.A1(\decode.regfile.registers_4[28] ),
    .A2(_09095_),
    .B1(_09105_),
    .C1(_09100_),
    .X(_02411_));
 sky130_fd_sc_hd__nand2_2 _25671_ (.A(_08970_),
    .B(_09067_),
    .Y(_09106_));
 sky130_fd_sc_hd__o211a_2 _25672_ (.A1(\decode.regfile.registers_4[29] ),
    .A2(_09095_),
    .B1(_09106_),
    .C1(_09100_),
    .X(_02412_));
 sky130_fd_sc_hd__nand2_2 _25673_ (.A(_08973_),
    .B(_09067_),
    .Y(_09107_));
 sky130_fd_sc_hd__o211a_2 _25674_ (.A1(\decode.regfile.registers_4[30] ),
    .A2(_09069_),
    .B1(_09107_),
    .C1(_09100_),
    .X(_02413_));
 sky130_fd_sc_hd__nand2_2 _25675_ (.A(_08975_),
    .B(_09067_),
    .Y(_09108_));
 sky130_fd_sc_hd__o211a_2 _25676_ (.A1(\decode.regfile.registers_4[31] ),
    .A2(_09069_),
    .B1(_09108_),
    .C1(_09100_),
    .X(_02414_));
 sky130_fd_sc_hd__and4_2 _25677_ (.A(_10373_),
    .B(_10240_),
    .C(_08903_),
    .D(_09935_),
    .X(_09109_));
 sky130_fd_sc_hd__buf_1 _25678_ (.A(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__buf_1 _25679_ (.A(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__buf_1 _25680_ (.A(_09110_),
    .X(_09112_));
 sky130_fd_sc_hd__nand2_2 _25681_ (.A(_09025_),
    .B(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__o211a_2 _25682_ (.A1(\decode.regfile.registers_5[0] ),
    .A2(_09111_),
    .B1(_09113_),
    .C1(_09100_),
    .X(_02415_));
 sky130_fd_sc_hd__nand2_2 _25683_ (.A(_08982_),
    .B(_09112_),
    .Y(_09114_));
 sky130_fd_sc_hd__buf_1 _25684_ (.A(_08990_),
    .X(_09115_));
 sky130_fd_sc_hd__o211a_2 _25685_ (.A1(\decode.regfile.registers_5[1] ),
    .A2(_09111_),
    .B1(_09114_),
    .C1(_09115_),
    .X(_02416_));
 sky130_fd_sc_hd__nand2_2 _25686_ (.A(_08910_),
    .B(_09112_),
    .Y(_09116_));
 sky130_fd_sc_hd__o211a_2 _25687_ (.A1(\decode.regfile.registers_5[2] ),
    .A2(_09111_),
    .B1(_09116_),
    .C1(_09115_),
    .X(_02417_));
 sky130_fd_sc_hd__nand2_2 _25688_ (.A(_08912_),
    .B(_09112_),
    .Y(_09117_));
 sky130_fd_sc_hd__o211a_2 _25689_ (.A1(\decode.regfile.registers_5[3] ),
    .A2(_09111_),
    .B1(_09117_),
    .C1(_09115_),
    .X(_02418_));
 sky130_fd_sc_hd__nand2_2 _25690_ (.A(_08914_),
    .B(_09112_),
    .Y(_09118_));
 sky130_fd_sc_hd__o211a_2 _25691_ (.A1(\decode.regfile.registers_5[4] ),
    .A2(_09111_),
    .B1(_09118_),
    .C1(_09115_),
    .X(_02419_));
 sky130_fd_sc_hd__nand2_2 _25692_ (.A(_08916_),
    .B(_09112_),
    .Y(_09119_));
 sky130_fd_sc_hd__o211a_2 _25693_ (.A1(\decode.regfile.registers_5[5] ),
    .A2(_09111_),
    .B1(_09119_),
    .C1(_09115_),
    .X(_02420_));
 sky130_fd_sc_hd__nand2_2 _25694_ (.A(_08918_),
    .B(_09112_),
    .Y(_09120_));
 sky130_fd_sc_hd__o211a_2 _25695_ (.A1(\decode.regfile.registers_5[6] ),
    .A2(_09111_),
    .B1(_09120_),
    .C1(_09115_),
    .X(_02421_));
 sky130_fd_sc_hd__nand2_2 _25696_ (.A(_08920_),
    .B(_09112_),
    .Y(_09121_));
 sky130_fd_sc_hd__o211a_2 _25697_ (.A1(\decode.regfile.registers_5[7] ),
    .A2(_09111_),
    .B1(_09121_),
    .C1(_09115_),
    .X(_02422_));
 sky130_fd_sc_hd__buf_1 _25698_ (.A(_09110_),
    .X(_09122_));
 sky130_fd_sc_hd__nand2_2 _25699_ (.A(_08922_),
    .B(_09122_),
    .Y(_09123_));
 sky130_fd_sc_hd__o211a_2 _25700_ (.A1(\decode.regfile.registers_5[8] ),
    .A2(_09111_),
    .B1(_09123_),
    .C1(_09115_),
    .X(_02423_));
 sky130_fd_sc_hd__nand2_2 _25701_ (.A(_08925_),
    .B(_09122_),
    .Y(_09124_));
 sky130_fd_sc_hd__o211a_2 _25702_ (.A1(\decode.regfile.registers_5[9] ),
    .A2(_09111_),
    .B1(_09124_),
    .C1(_09115_),
    .X(_02424_));
 sky130_fd_sc_hd__buf_1 _25703_ (.A(_09110_),
    .X(_09125_));
 sky130_fd_sc_hd__nand2_2 _25704_ (.A(_08929_),
    .B(_09122_),
    .Y(_09126_));
 sky130_fd_sc_hd__o211a_2 _25705_ (.A1(\decode.regfile.registers_5[10] ),
    .A2(_09125_),
    .B1(_09126_),
    .C1(_09115_),
    .X(_02425_));
 sky130_fd_sc_hd__nand2_2 _25706_ (.A(_08931_),
    .B(_09122_),
    .Y(_09127_));
 sky130_fd_sc_hd__buf_1 _25707_ (.A(_10130_),
    .X(_09128_));
 sky130_fd_sc_hd__buf_1 _25708_ (.A(_09128_),
    .X(_09129_));
 sky130_fd_sc_hd__o211a_2 _25709_ (.A1(\decode.regfile.registers_5[11] ),
    .A2(_09125_),
    .B1(_09127_),
    .C1(_09129_),
    .X(_02426_));
 sky130_fd_sc_hd__nand2_2 _25710_ (.A(_08933_),
    .B(_09122_),
    .Y(_09130_));
 sky130_fd_sc_hd__o211a_2 _25711_ (.A1(\decode.regfile.registers_5[12] ),
    .A2(_09125_),
    .B1(_09130_),
    .C1(_09129_),
    .X(_02427_));
 sky130_fd_sc_hd__nand2_2 _25712_ (.A(_08935_),
    .B(_09122_),
    .Y(_09131_));
 sky130_fd_sc_hd__o211a_2 _25713_ (.A1(\decode.regfile.registers_5[13] ),
    .A2(_09125_),
    .B1(_09131_),
    .C1(_09129_),
    .X(_02428_));
 sky130_fd_sc_hd__nand2_2 _25714_ (.A(_08937_),
    .B(_09122_),
    .Y(_09132_));
 sky130_fd_sc_hd__o211a_2 _25715_ (.A1(\decode.regfile.registers_5[14] ),
    .A2(_09125_),
    .B1(_09132_),
    .C1(_09129_),
    .X(_02429_));
 sky130_fd_sc_hd__nand2_2 _25716_ (.A(_08939_),
    .B(_09122_),
    .Y(_09133_));
 sky130_fd_sc_hd__o211a_2 _25717_ (.A1(\decode.regfile.registers_5[15] ),
    .A2(_09125_),
    .B1(_09133_),
    .C1(_09129_),
    .X(_02430_));
 sky130_fd_sc_hd__nand2_2 _25718_ (.A(_08941_),
    .B(_09122_),
    .Y(_09134_));
 sky130_fd_sc_hd__o211a_2 _25719_ (.A1(\decode.regfile.registers_5[16] ),
    .A2(_09125_),
    .B1(_09134_),
    .C1(_09129_),
    .X(_02431_));
 sky130_fd_sc_hd__nand2_2 _25720_ (.A(_08943_),
    .B(_09122_),
    .Y(_09135_));
 sky130_fd_sc_hd__o211a_2 _25721_ (.A1(\decode.regfile.registers_5[17] ),
    .A2(_09125_),
    .B1(_09135_),
    .C1(_09129_),
    .X(_02432_));
 sky130_fd_sc_hd__buf_1 _25722_ (.A(_09110_),
    .X(_09136_));
 sky130_fd_sc_hd__nand2_2 _25723_ (.A(_08945_),
    .B(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__o211a_2 _25724_ (.A1(\decode.regfile.registers_5[18] ),
    .A2(_09125_),
    .B1(_09137_),
    .C1(_09129_),
    .X(_02433_));
 sky130_fd_sc_hd__nand2_2 _25725_ (.A(_08948_),
    .B(_09136_),
    .Y(_09138_));
 sky130_fd_sc_hd__o211a_2 _25726_ (.A1(\decode.regfile.registers_5[19] ),
    .A2(_09125_),
    .B1(_09138_),
    .C1(_09129_),
    .X(_02434_));
 sky130_fd_sc_hd__buf_1 _25727_ (.A(_09110_),
    .X(_09139_));
 sky130_fd_sc_hd__nand2_2 _25728_ (.A(_08952_),
    .B(_09136_),
    .Y(_09140_));
 sky130_fd_sc_hd__o211a_2 _25729_ (.A1(\decode.regfile.registers_5[20] ),
    .A2(_09139_),
    .B1(_09140_),
    .C1(_09129_),
    .X(_02435_));
 sky130_fd_sc_hd__nand2_2 _25730_ (.A(_08954_),
    .B(_09136_),
    .Y(_09141_));
 sky130_fd_sc_hd__buf_1 _25731_ (.A(_09128_),
    .X(_09142_));
 sky130_fd_sc_hd__o211a_2 _25732_ (.A1(\decode.regfile.registers_5[21] ),
    .A2(_09139_),
    .B1(_09141_),
    .C1(_09142_),
    .X(_02436_));
 sky130_fd_sc_hd__nand2_2 _25733_ (.A(_08956_),
    .B(_09136_),
    .Y(_09143_));
 sky130_fd_sc_hd__o211a_2 _25734_ (.A1(\decode.regfile.registers_5[22] ),
    .A2(_09139_),
    .B1(_09143_),
    .C1(_09142_),
    .X(_02437_));
 sky130_fd_sc_hd__nand2_2 _25735_ (.A(_08958_),
    .B(_09136_),
    .Y(_09144_));
 sky130_fd_sc_hd__o211a_2 _25736_ (.A1(\decode.regfile.registers_5[23] ),
    .A2(_09139_),
    .B1(_09144_),
    .C1(_09142_),
    .X(_02438_));
 sky130_fd_sc_hd__nand2_2 _25737_ (.A(_08960_),
    .B(_09136_),
    .Y(_09145_));
 sky130_fd_sc_hd__o211a_2 _25738_ (.A1(\decode.regfile.registers_5[24] ),
    .A2(_09139_),
    .B1(_09145_),
    .C1(_09142_),
    .X(_02439_));
 sky130_fd_sc_hd__nand2_2 _25739_ (.A(_08962_),
    .B(_09136_),
    .Y(_09146_));
 sky130_fd_sc_hd__o211a_2 _25740_ (.A1(\decode.regfile.registers_5[25] ),
    .A2(_09139_),
    .B1(_09146_),
    .C1(_09142_),
    .X(_02440_));
 sky130_fd_sc_hd__nand2_2 _25741_ (.A(_08964_),
    .B(_09136_),
    .Y(_09147_));
 sky130_fd_sc_hd__o211a_2 _25742_ (.A1(\decode.regfile.registers_5[26] ),
    .A2(_09139_),
    .B1(_09147_),
    .C1(_09142_),
    .X(_02441_));
 sky130_fd_sc_hd__nand2_2 _25743_ (.A(_08966_),
    .B(_09136_),
    .Y(_09148_));
 sky130_fd_sc_hd__o211a_2 _25744_ (.A1(\decode.regfile.registers_5[27] ),
    .A2(_09139_),
    .B1(_09148_),
    .C1(_09142_),
    .X(_02442_));
 sky130_fd_sc_hd__nand2_2 _25745_ (.A(_08968_),
    .B(_09110_),
    .Y(_09149_));
 sky130_fd_sc_hd__o211a_2 _25746_ (.A1(\decode.regfile.registers_5[28] ),
    .A2(_09139_),
    .B1(_09149_),
    .C1(_09142_),
    .X(_02443_));
 sky130_fd_sc_hd__nand2_2 _25747_ (.A(_08970_),
    .B(_09110_),
    .Y(_09150_));
 sky130_fd_sc_hd__o211a_2 _25748_ (.A1(\decode.regfile.registers_5[29] ),
    .A2(_09139_),
    .B1(_09150_),
    .C1(_09142_),
    .X(_02444_));
 sky130_fd_sc_hd__nand2_2 _25749_ (.A(_08973_),
    .B(_09110_),
    .Y(_09151_));
 sky130_fd_sc_hd__o211a_2 _25750_ (.A1(\decode.regfile.registers_5[30] ),
    .A2(_09112_),
    .B1(_09151_),
    .C1(_09142_),
    .X(_02445_));
 sky130_fd_sc_hd__nand2_2 _25751_ (.A(_08975_),
    .B(_09110_),
    .Y(_09152_));
 sky130_fd_sc_hd__buf_1 _25752_ (.A(_09128_),
    .X(_09153_));
 sky130_fd_sc_hd__o211a_2 _25753_ (.A1(\decode.regfile.registers_5[31] ),
    .A2(_09112_),
    .B1(_09152_),
    .C1(_09153_),
    .X(_02446_));
 sky130_fd_sc_hd__and4_2 _25754_ (.A(_10373_),
    .B(_09932_),
    .C(_08903_),
    .D(_09935_),
    .X(_09154_));
 sky130_fd_sc_hd__buf_1 _25755_ (.A(_09154_),
    .X(_09155_));
 sky130_fd_sc_hd__buf_1 _25756_ (.A(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__buf_1 _25757_ (.A(_09155_),
    .X(_09157_));
 sky130_fd_sc_hd__nand2_2 _25758_ (.A(_09025_),
    .B(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__o211a_2 _25759_ (.A1(\decode.regfile.registers_6[0] ),
    .A2(_09156_),
    .B1(_09158_),
    .C1(_09153_),
    .X(_02447_));
 sky130_fd_sc_hd__nand2_2 _25760_ (.A(_08982_),
    .B(_09157_),
    .Y(_09159_));
 sky130_fd_sc_hd__o211a_2 _25761_ (.A1(\decode.regfile.registers_6[1] ),
    .A2(_09156_),
    .B1(_09159_),
    .C1(_09153_),
    .X(_02448_));
 sky130_fd_sc_hd__nand2_2 _25762_ (.A(_08910_),
    .B(_09157_),
    .Y(_09160_));
 sky130_fd_sc_hd__o211a_2 _25763_ (.A1(\decode.regfile.registers_6[2] ),
    .A2(_09156_),
    .B1(_09160_),
    .C1(_09153_),
    .X(_02449_));
 sky130_fd_sc_hd__nand2_2 _25764_ (.A(_08912_),
    .B(_09157_),
    .Y(_09161_));
 sky130_fd_sc_hd__o211a_2 _25765_ (.A1(\decode.regfile.registers_6[3] ),
    .A2(_09156_),
    .B1(_09161_),
    .C1(_09153_),
    .X(_02450_));
 sky130_fd_sc_hd__nand2_2 _25766_ (.A(_08914_),
    .B(_09157_),
    .Y(_09162_));
 sky130_fd_sc_hd__o211a_2 _25767_ (.A1(\decode.regfile.registers_6[4] ),
    .A2(_09156_),
    .B1(_09162_),
    .C1(_09153_),
    .X(_02451_));
 sky130_fd_sc_hd__nand2_2 _25768_ (.A(_08916_),
    .B(_09157_),
    .Y(_09163_));
 sky130_fd_sc_hd__o211a_2 _25769_ (.A1(\decode.regfile.registers_6[5] ),
    .A2(_09156_),
    .B1(_09163_),
    .C1(_09153_),
    .X(_02452_));
 sky130_fd_sc_hd__nand2_2 _25770_ (.A(_08918_),
    .B(_09157_),
    .Y(_09164_));
 sky130_fd_sc_hd__o211a_2 _25771_ (.A1(\decode.regfile.registers_6[6] ),
    .A2(_09156_),
    .B1(_09164_),
    .C1(_09153_),
    .X(_02453_));
 sky130_fd_sc_hd__nand2_2 _25772_ (.A(_08920_),
    .B(_09157_),
    .Y(_09165_));
 sky130_fd_sc_hd__o211a_2 _25773_ (.A1(\decode.regfile.registers_6[7] ),
    .A2(_09156_),
    .B1(_09165_),
    .C1(_09153_),
    .X(_02454_));
 sky130_fd_sc_hd__buf_1 _25774_ (.A(_09155_),
    .X(_09166_));
 sky130_fd_sc_hd__nand2_2 _25775_ (.A(_08922_),
    .B(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__o211a_2 _25776_ (.A1(\decode.regfile.registers_6[8] ),
    .A2(_09156_),
    .B1(_09167_),
    .C1(_09153_),
    .X(_02455_));
 sky130_fd_sc_hd__nand2_2 _25777_ (.A(_08925_),
    .B(_09166_),
    .Y(_09168_));
 sky130_fd_sc_hd__buf_1 _25778_ (.A(_09128_),
    .X(_09169_));
 sky130_fd_sc_hd__o211a_2 _25779_ (.A1(\decode.regfile.registers_6[9] ),
    .A2(_09156_),
    .B1(_09168_),
    .C1(_09169_),
    .X(_02456_));
 sky130_fd_sc_hd__buf_1 _25780_ (.A(_09155_),
    .X(_09170_));
 sky130_fd_sc_hd__nand2_2 _25781_ (.A(_08929_),
    .B(_09166_),
    .Y(_09171_));
 sky130_fd_sc_hd__o211a_2 _25782_ (.A1(\decode.regfile.registers_6[10] ),
    .A2(_09170_),
    .B1(_09171_),
    .C1(_09169_),
    .X(_02457_));
 sky130_fd_sc_hd__nand2_2 _25783_ (.A(_08931_),
    .B(_09166_),
    .Y(_09172_));
 sky130_fd_sc_hd__o211a_2 _25784_ (.A1(\decode.regfile.registers_6[11] ),
    .A2(_09170_),
    .B1(_09172_),
    .C1(_09169_),
    .X(_02458_));
 sky130_fd_sc_hd__nand2_2 _25785_ (.A(_08933_),
    .B(_09166_),
    .Y(_09173_));
 sky130_fd_sc_hd__o211a_2 _25786_ (.A1(\decode.regfile.registers_6[12] ),
    .A2(_09170_),
    .B1(_09173_),
    .C1(_09169_),
    .X(_02459_));
 sky130_fd_sc_hd__nand2_2 _25787_ (.A(_08935_),
    .B(_09166_),
    .Y(_09174_));
 sky130_fd_sc_hd__o211a_2 _25788_ (.A1(\decode.regfile.registers_6[13] ),
    .A2(_09170_),
    .B1(_09174_),
    .C1(_09169_),
    .X(_02460_));
 sky130_fd_sc_hd__nand2_2 _25789_ (.A(_08937_),
    .B(_09166_),
    .Y(_09175_));
 sky130_fd_sc_hd__o211a_2 _25790_ (.A1(\decode.regfile.registers_6[14] ),
    .A2(_09170_),
    .B1(_09175_),
    .C1(_09169_),
    .X(_02461_));
 sky130_fd_sc_hd__nand2_2 _25791_ (.A(_08939_),
    .B(_09166_),
    .Y(_09176_));
 sky130_fd_sc_hd__o211a_2 _25792_ (.A1(\decode.regfile.registers_6[15] ),
    .A2(_09170_),
    .B1(_09176_),
    .C1(_09169_),
    .X(_02462_));
 sky130_fd_sc_hd__nand2_2 _25793_ (.A(_08941_),
    .B(_09166_),
    .Y(_09177_));
 sky130_fd_sc_hd__o211a_2 _25794_ (.A1(\decode.regfile.registers_6[16] ),
    .A2(_09170_),
    .B1(_09177_),
    .C1(_09169_),
    .X(_02463_));
 sky130_fd_sc_hd__nand2_2 _25795_ (.A(_08943_),
    .B(_09166_),
    .Y(_09178_));
 sky130_fd_sc_hd__o211a_2 _25796_ (.A1(\decode.regfile.registers_6[17] ),
    .A2(_09170_),
    .B1(_09178_),
    .C1(_09169_),
    .X(_02464_));
 sky130_fd_sc_hd__buf_1 _25797_ (.A(_09155_),
    .X(_09179_));
 sky130_fd_sc_hd__nand2_2 _25798_ (.A(_08945_),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__o211a_2 _25799_ (.A1(\decode.regfile.registers_6[18] ),
    .A2(_09170_),
    .B1(_09180_),
    .C1(_09169_),
    .X(_02465_));
 sky130_fd_sc_hd__nand2_2 _25800_ (.A(_08948_),
    .B(_09179_),
    .Y(_09181_));
 sky130_fd_sc_hd__buf_1 _25801_ (.A(_09128_),
    .X(_09182_));
 sky130_fd_sc_hd__o211a_2 _25802_ (.A1(\decode.regfile.registers_6[19] ),
    .A2(_09170_),
    .B1(_09181_),
    .C1(_09182_),
    .X(_02466_));
 sky130_fd_sc_hd__buf_1 _25803_ (.A(_09155_),
    .X(_09183_));
 sky130_fd_sc_hd__nand2_2 _25804_ (.A(_08952_),
    .B(_09179_),
    .Y(_09184_));
 sky130_fd_sc_hd__o211a_2 _25805_ (.A1(\decode.regfile.registers_6[20] ),
    .A2(_09183_),
    .B1(_09184_),
    .C1(_09182_),
    .X(_02467_));
 sky130_fd_sc_hd__nand2_2 _25806_ (.A(_08954_),
    .B(_09179_),
    .Y(_09185_));
 sky130_fd_sc_hd__o211a_2 _25807_ (.A1(\decode.regfile.registers_6[21] ),
    .A2(_09183_),
    .B1(_09185_),
    .C1(_09182_),
    .X(_02468_));
 sky130_fd_sc_hd__nand2_2 _25808_ (.A(_08956_),
    .B(_09179_),
    .Y(_09186_));
 sky130_fd_sc_hd__o211a_2 _25809_ (.A1(\decode.regfile.registers_6[22] ),
    .A2(_09183_),
    .B1(_09186_),
    .C1(_09182_),
    .X(_02469_));
 sky130_fd_sc_hd__nand2_2 _25810_ (.A(_08958_),
    .B(_09179_),
    .Y(_09187_));
 sky130_fd_sc_hd__o211a_2 _25811_ (.A1(\decode.regfile.registers_6[23] ),
    .A2(_09183_),
    .B1(_09187_),
    .C1(_09182_),
    .X(_02470_));
 sky130_fd_sc_hd__nand2_2 _25812_ (.A(_08960_),
    .B(_09179_),
    .Y(_09188_));
 sky130_fd_sc_hd__o211a_2 _25813_ (.A1(\decode.regfile.registers_6[24] ),
    .A2(_09183_),
    .B1(_09188_),
    .C1(_09182_),
    .X(_02471_));
 sky130_fd_sc_hd__nand2_2 _25814_ (.A(_08962_),
    .B(_09179_),
    .Y(_09189_));
 sky130_fd_sc_hd__o211a_2 _25815_ (.A1(\decode.regfile.registers_6[25] ),
    .A2(_09183_),
    .B1(_09189_),
    .C1(_09182_),
    .X(_02472_));
 sky130_fd_sc_hd__nand2_2 _25816_ (.A(_08964_),
    .B(_09179_),
    .Y(_09190_));
 sky130_fd_sc_hd__o211a_2 _25817_ (.A1(\decode.regfile.registers_6[26] ),
    .A2(_09183_),
    .B1(_09190_),
    .C1(_09182_),
    .X(_02473_));
 sky130_fd_sc_hd__nand2_2 _25818_ (.A(_08966_),
    .B(_09179_),
    .Y(_09191_));
 sky130_fd_sc_hd__o211a_2 _25819_ (.A1(\decode.regfile.registers_6[27] ),
    .A2(_09183_),
    .B1(_09191_),
    .C1(_09182_),
    .X(_02474_));
 sky130_fd_sc_hd__nand2_2 _25820_ (.A(_08968_),
    .B(_09155_),
    .Y(_09192_));
 sky130_fd_sc_hd__o211a_2 _25821_ (.A1(\decode.regfile.registers_6[28] ),
    .A2(_09183_),
    .B1(_09192_),
    .C1(_09182_),
    .X(_02475_));
 sky130_fd_sc_hd__nand2_2 _25822_ (.A(_08970_),
    .B(_09155_),
    .Y(_09193_));
 sky130_fd_sc_hd__buf_1 _25823_ (.A(_09128_),
    .X(_09194_));
 sky130_fd_sc_hd__o211a_2 _25824_ (.A1(\decode.regfile.registers_6[29] ),
    .A2(_09183_),
    .B1(_09193_),
    .C1(_09194_),
    .X(_02476_));
 sky130_fd_sc_hd__nand2_2 _25825_ (.A(_08973_),
    .B(_09155_),
    .Y(_09195_));
 sky130_fd_sc_hd__o211a_2 _25826_ (.A1(\decode.regfile.registers_6[30] ),
    .A2(_09157_),
    .B1(_09195_),
    .C1(_09194_),
    .X(_02477_));
 sky130_fd_sc_hd__nand2_2 _25827_ (.A(_08975_),
    .B(_09155_),
    .Y(_09196_));
 sky130_fd_sc_hd__o211a_2 _25828_ (.A1(\decode.regfile.registers_6[31] ),
    .A2(_09157_),
    .B1(_09196_),
    .C1(_09194_),
    .X(_02478_));
 sky130_fd_sc_hd__and4_2 _25829_ (.A(_10373_),
    .B(_10150_),
    .C(_08902_),
    .D(_09935_),
    .X(_09197_));
 sky130_fd_sc_hd__buf_1 _25830_ (.A(_09197_),
    .X(_09198_));
 sky130_fd_sc_hd__buf_1 _25831_ (.A(_09198_),
    .X(_09199_));
 sky130_fd_sc_hd__buf_1 _25832_ (.A(_09198_),
    .X(_09200_));
 sky130_fd_sc_hd__nand2_2 _25833_ (.A(_09025_),
    .B(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__o211a_2 _25834_ (.A1(\decode.regfile.registers_7[0] ),
    .A2(_09199_),
    .B1(_09201_),
    .C1(_09194_),
    .X(_02479_));
 sky130_fd_sc_hd__nand2_2 _25835_ (.A(_08982_),
    .B(_09200_),
    .Y(_09202_));
 sky130_fd_sc_hd__o211a_2 _25836_ (.A1(\decode.regfile.registers_7[1] ),
    .A2(_09199_),
    .B1(_09202_),
    .C1(_09194_),
    .X(_02480_));
 sky130_fd_sc_hd__nand2_2 _25837_ (.A(_08910_),
    .B(_09200_),
    .Y(_09203_));
 sky130_fd_sc_hd__o211a_2 _25838_ (.A1(\decode.regfile.registers_7[2] ),
    .A2(_09199_),
    .B1(_09203_),
    .C1(_09194_),
    .X(_02481_));
 sky130_fd_sc_hd__nand2_2 _25839_ (.A(_08912_),
    .B(_09200_),
    .Y(_09204_));
 sky130_fd_sc_hd__o211a_2 _25840_ (.A1(\decode.regfile.registers_7[3] ),
    .A2(_09199_),
    .B1(_09204_),
    .C1(_09194_),
    .X(_02482_));
 sky130_fd_sc_hd__nand2_2 _25841_ (.A(_08914_),
    .B(_09200_),
    .Y(_09205_));
 sky130_fd_sc_hd__o211a_2 _25842_ (.A1(\decode.regfile.registers_7[4] ),
    .A2(_09199_),
    .B1(_09205_),
    .C1(_09194_),
    .X(_02483_));
 sky130_fd_sc_hd__nand2_2 _25843_ (.A(_08916_),
    .B(_09200_),
    .Y(_09206_));
 sky130_fd_sc_hd__o211a_2 _25844_ (.A1(\decode.regfile.registers_7[5] ),
    .A2(_09199_),
    .B1(_09206_),
    .C1(_09194_),
    .X(_02484_));
 sky130_fd_sc_hd__nand2_2 _25845_ (.A(_08918_),
    .B(_09200_),
    .Y(_09207_));
 sky130_fd_sc_hd__o211a_2 _25846_ (.A1(\decode.regfile.registers_7[6] ),
    .A2(_09199_),
    .B1(_09207_),
    .C1(_09194_),
    .X(_02485_));
 sky130_fd_sc_hd__nand2_2 _25847_ (.A(_08920_),
    .B(_09200_),
    .Y(_09208_));
 sky130_fd_sc_hd__buf_1 _25848_ (.A(_09128_),
    .X(_09209_));
 sky130_fd_sc_hd__o211a_2 _25849_ (.A1(\decode.regfile.registers_7[7] ),
    .A2(_09199_),
    .B1(_09208_),
    .C1(_09209_),
    .X(_02486_));
 sky130_fd_sc_hd__buf_1 _25850_ (.A(_09198_),
    .X(_09210_));
 sky130_fd_sc_hd__nand2_2 _25851_ (.A(_08922_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__o211a_2 _25852_ (.A1(\decode.regfile.registers_7[8] ),
    .A2(_09199_),
    .B1(_09211_),
    .C1(_09209_),
    .X(_02487_));
 sky130_fd_sc_hd__nand2_2 _25853_ (.A(_08925_),
    .B(_09210_),
    .Y(_09212_));
 sky130_fd_sc_hd__o211a_2 _25854_ (.A1(\decode.regfile.registers_7[9] ),
    .A2(_09199_),
    .B1(_09212_),
    .C1(_09209_),
    .X(_02488_));
 sky130_fd_sc_hd__buf_1 _25855_ (.A(_09198_),
    .X(_09213_));
 sky130_fd_sc_hd__nand2_2 _25856_ (.A(_08929_),
    .B(_09210_),
    .Y(_09214_));
 sky130_fd_sc_hd__o211a_2 _25857_ (.A1(\decode.regfile.registers_7[10] ),
    .A2(_09213_),
    .B1(_09214_),
    .C1(_09209_),
    .X(_02489_));
 sky130_fd_sc_hd__nand2_2 _25858_ (.A(_08931_),
    .B(_09210_),
    .Y(_09215_));
 sky130_fd_sc_hd__o211a_2 _25859_ (.A1(\decode.regfile.registers_7[11] ),
    .A2(_09213_),
    .B1(_09215_),
    .C1(_09209_),
    .X(_02490_));
 sky130_fd_sc_hd__nand2_2 _25860_ (.A(_08933_),
    .B(_09210_),
    .Y(_09216_));
 sky130_fd_sc_hd__o211a_2 _25861_ (.A1(\decode.regfile.registers_7[12] ),
    .A2(_09213_),
    .B1(_09216_),
    .C1(_09209_),
    .X(_02491_));
 sky130_fd_sc_hd__nand2_2 _25862_ (.A(_08935_),
    .B(_09210_),
    .Y(_09217_));
 sky130_fd_sc_hd__o211a_2 _25863_ (.A1(\decode.regfile.registers_7[13] ),
    .A2(_09213_),
    .B1(_09217_),
    .C1(_09209_),
    .X(_02492_));
 sky130_fd_sc_hd__nand2_2 _25864_ (.A(_08937_),
    .B(_09210_),
    .Y(_09218_));
 sky130_fd_sc_hd__o211a_2 _25865_ (.A1(\decode.regfile.registers_7[14] ),
    .A2(_09213_),
    .B1(_09218_),
    .C1(_09209_),
    .X(_02493_));
 sky130_fd_sc_hd__nand2_2 _25866_ (.A(_08939_),
    .B(_09210_),
    .Y(_09219_));
 sky130_fd_sc_hd__o211a_2 _25867_ (.A1(\decode.regfile.registers_7[15] ),
    .A2(_09213_),
    .B1(_09219_),
    .C1(_09209_),
    .X(_02494_));
 sky130_fd_sc_hd__nand2_2 _25868_ (.A(_08941_),
    .B(_09210_),
    .Y(_09220_));
 sky130_fd_sc_hd__o211a_2 _25869_ (.A1(\decode.regfile.registers_7[16] ),
    .A2(_09213_),
    .B1(_09220_),
    .C1(_09209_),
    .X(_02495_));
 sky130_fd_sc_hd__nand2_2 _25870_ (.A(_08943_),
    .B(_09210_),
    .Y(_09221_));
 sky130_fd_sc_hd__buf_1 _25871_ (.A(_09128_),
    .X(_09222_));
 sky130_fd_sc_hd__o211a_2 _25872_ (.A1(\decode.regfile.registers_7[17] ),
    .A2(_09213_),
    .B1(_09221_),
    .C1(_09222_),
    .X(_02496_));
 sky130_fd_sc_hd__buf_1 _25873_ (.A(_09198_),
    .X(_09223_));
 sky130_fd_sc_hd__nand2_2 _25874_ (.A(_08945_),
    .B(_09223_),
    .Y(_09224_));
 sky130_fd_sc_hd__o211a_2 _25875_ (.A1(\decode.regfile.registers_7[18] ),
    .A2(_09213_),
    .B1(_09224_),
    .C1(_09222_),
    .X(_02497_));
 sky130_fd_sc_hd__nand2_2 _25876_ (.A(_08948_),
    .B(_09223_),
    .Y(_09225_));
 sky130_fd_sc_hd__o211a_2 _25877_ (.A1(\decode.regfile.registers_7[19] ),
    .A2(_09213_),
    .B1(_09225_),
    .C1(_09222_),
    .X(_02498_));
 sky130_fd_sc_hd__buf_1 _25878_ (.A(_09198_),
    .X(_09226_));
 sky130_fd_sc_hd__nand2_2 _25879_ (.A(_08952_),
    .B(_09223_),
    .Y(_09227_));
 sky130_fd_sc_hd__o211a_2 _25880_ (.A1(\decode.regfile.registers_7[20] ),
    .A2(_09226_),
    .B1(_09227_),
    .C1(_09222_),
    .X(_02499_));
 sky130_fd_sc_hd__nand2_2 _25881_ (.A(_08954_),
    .B(_09223_),
    .Y(_09228_));
 sky130_fd_sc_hd__o211a_2 _25882_ (.A1(\decode.regfile.registers_7[21] ),
    .A2(_09226_),
    .B1(_09228_),
    .C1(_09222_),
    .X(_02500_));
 sky130_fd_sc_hd__nand2_2 _25883_ (.A(_08956_),
    .B(_09223_),
    .Y(_09229_));
 sky130_fd_sc_hd__o211a_2 _25884_ (.A1(\decode.regfile.registers_7[22] ),
    .A2(_09226_),
    .B1(_09229_),
    .C1(_09222_),
    .X(_02501_));
 sky130_fd_sc_hd__nand2_2 _25885_ (.A(_08958_),
    .B(_09223_),
    .Y(_09230_));
 sky130_fd_sc_hd__o211a_2 _25886_ (.A1(\decode.regfile.registers_7[23] ),
    .A2(_09226_),
    .B1(_09230_),
    .C1(_09222_),
    .X(_02502_));
 sky130_fd_sc_hd__nand2_2 _25887_ (.A(_08960_),
    .B(_09223_),
    .Y(_09231_));
 sky130_fd_sc_hd__o211a_2 _25888_ (.A1(\decode.regfile.registers_7[24] ),
    .A2(_09226_),
    .B1(_09231_),
    .C1(_09222_),
    .X(_02503_));
 sky130_fd_sc_hd__nand2_2 _25889_ (.A(_08962_),
    .B(_09223_),
    .Y(_09232_));
 sky130_fd_sc_hd__o211a_2 _25890_ (.A1(\decode.regfile.registers_7[25] ),
    .A2(_09226_),
    .B1(_09232_),
    .C1(_09222_),
    .X(_02504_));
 sky130_fd_sc_hd__nand2_2 _25891_ (.A(_08964_),
    .B(_09223_),
    .Y(_09233_));
 sky130_fd_sc_hd__o211a_2 _25892_ (.A1(\decode.regfile.registers_7[26] ),
    .A2(_09226_),
    .B1(_09233_),
    .C1(_09222_),
    .X(_02505_));
 sky130_fd_sc_hd__nand2_2 _25893_ (.A(_08966_),
    .B(_09223_),
    .Y(_09234_));
 sky130_fd_sc_hd__buf_1 _25894_ (.A(_09128_),
    .X(_09235_));
 sky130_fd_sc_hd__o211a_2 _25895_ (.A1(\decode.regfile.registers_7[27] ),
    .A2(_09226_),
    .B1(_09234_),
    .C1(_09235_),
    .X(_02506_));
 sky130_fd_sc_hd__nand2_2 _25896_ (.A(_08968_),
    .B(_09198_),
    .Y(_09236_));
 sky130_fd_sc_hd__o211a_2 _25897_ (.A1(\decode.regfile.registers_7[28] ),
    .A2(_09226_),
    .B1(_09236_),
    .C1(_09235_),
    .X(_02507_));
 sky130_fd_sc_hd__nand2_2 _25898_ (.A(_08970_),
    .B(_09198_),
    .Y(_09237_));
 sky130_fd_sc_hd__o211a_2 _25899_ (.A1(\decode.regfile.registers_7[29] ),
    .A2(_09226_),
    .B1(_09237_),
    .C1(_09235_),
    .X(_02508_));
 sky130_fd_sc_hd__nand2_2 _25900_ (.A(_08973_),
    .B(_09198_),
    .Y(_09238_));
 sky130_fd_sc_hd__o211a_2 _25901_ (.A1(\decode.regfile.registers_7[30] ),
    .A2(_09200_),
    .B1(_09238_),
    .C1(_09235_),
    .X(_02509_));
 sky130_fd_sc_hd__nand2_2 _25902_ (.A(_08975_),
    .B(_09198_),
    .Y(_09239_));
 sky130_fd_sc_hd__o211a_2 _25903_ (.A1(\decode.regfile.registers_7[31] ),
    .A2(_09200_),
    .B1(_09239_),
    .C1(_09235_),
    .X(_02510_));
 sky130_fd_sc_hd__and4b_2 _25904_ (.A_N(_09930_),
    .B(_10194_),
    .C(_10196_),
    .D(_08902_),
    .X(_09240_));
 sky130_fd_sc_hd__buf_1 _25905_ (.A(_09240_),
    .X(_09241_));
 sky130_fd_sc_hd__buf_1 _25906_ (.A(_09241_),
    .X(_09242_));
 sky130_fd_sc_hd__buf_1 _25907_ (.A(_09241_),
    .X(_09243_));
 sky130_fd_sc_hd__nand2_2 _25908_ (.A(_09025_),
    .B(_09243_),
    .Y(_09244_));
 sky130_fd_sc_hd__o211a_2 _25909_ (.A1(\decode.regfile.registers_8[0] ),
    .A2(_09242_),
    .B1(_09244_),
    .C1(_09235_),
    .X(_02511_));
 sky130_fd_sc_hd__nand2_2 _25910_ (.A(_08982_),
    .B(_09243_),
    .Y(_09245_));
 sky130_fd_sc_hd__o211a_2 _25911_ (.A1(\decode.regfile.registers_8[1] ),
    .A2(_09242_),
    .B1(_09245_),
    .C1(_09235_),
    .X(_02512_));
 sky130_fd_sc_hd__nand2_2 _25912_ (.A(_08910_),
    .B(_09243_),
    .Y(_09246_));
 sky130_fd_sc_hd__o211a_2 _25913_ (.A1(\decode.regfile.registers_8[2] ),
    .A2(_09242_),
    .B1(_09246_),
    .C1(_09235_),
    .X(_02513_));
 sky130_fd_sc_hd__nand2_2 _25914_ (.A(_08912_),
    .B(_09243_),
    .Y(_09247_));
 sky130_fd_sc_hd__o211a_2 _25915_ (.A1(\decode.regfile.registers_8[3] ),
    .A2(_09242_),
    .B1(_09247_),
    .C1(_09235_),
    .X(_02514_));
 sky130_fd_sc_hd__nand2_2 _25916_ (.A(_08914_),
    .B(_09243_),
    .Y(_09248_));
 sky130_fd_sc_hd__o211a_2 _25917_ (.A1(\decode.regfile.registers_8[4] ),
    .A2(_09242_),
    .B1(_09248_),
    .C1(_09235_),
    .X(_02515_));
 sky130_fd_sc_hd__nand2_2 _25918_ (.A(_08916_),
    .B(_09243_),
    .Y(_09249_));
 sky130_fd_sc_hd__buf_1 _25919_ (.A(_09128_),
    .X(_09250_));
 sky130_fd_sc_hd__o211a_2 _25920_ (.A1(\decode.regfile.registers_8[5] ),
    .A2(_09242_),
    .B1(_09249_),
    .C1(_09250_),
    .X(_02516_));
 sky130_fd_sc_hd__nand2_2 _25921_ (.A(_08918_),
    .B(_09243_),
    .Y(_09251_));
 sky130_fd_sc_hd__o211a_2 _25922_ (.A1(\decode.regfile.registers_8[6] ),
    .A2(_09242_),
    .B1(_09251_),
    .C1(_09250_),
    .X(_02517_));
 sky130_fd_sc_hd__nand2_2 _25923_ (.A(_08920_),
    .B(_09243_),
    .Y(_09252_));
 sky130_fd_sc_hd__o211a_2 _25924_ (.A1(\decode.regfile.registers_8[7] ),
    .A2(_09242_),
    .B1(_09252_),
    .C1(_09250_),
    .X(_02518_));
 sky130_fd_sc_hd__buf_1 _25925_ (.A(_09241_),
    .X(_09253_));
 sky130_fd_sc_hd__nand2_2 _25926_ (.A(_08922_),
    .B(_09253_),
    .Y(_09254_));
 sky130_fd_sc_hd__o211a_2 _25927_ (.A1(\decode.regfile.registers_8[8] ),
    .A2(_09242_),
    .B1(_09254_),
    .C1(_09250_),
    .X(_02519_));
 sky130_fd_sc_hd__nand2_2 _25928_ (.A(_08925_),
    .B(_09253_),
    .Y(_09255_));
 sky130_fd_sc_hd__o211a_2 _25929_ (.A1(\decode.regfile.registers_8[9] ),
    .A2(_09242_),
    .B1(_09255_),
    .C1(_09250_),
    .X(_02520_));
 sky130_fd_sc_hd__buf_1 _25930_ (.A(_09241_),
    .X(_09256_));
 sky130_fd_sc_hd__nand2_2 _25931_ (.A(_08929_),
    .B(_09253_),
    .Y(_09257_));
 sky130_fd_sc_hd__o211a_2 _25932_ (.A1(\decode.regfile.registers_8[10] ),
    .A2(_09256_),
    .B1(_09257_),
    .C1(_09250_),
    .X(_02521_));
 sky130_fd_sc_hd__nand2_2 _25933_ (.A(_08931_),
    .B(_09253_),
    .Y(_09258_));
 sky130_fd_sc_hd__o211a_2 _25934_ (.A1(\decode.regfile.registers_8[11] ),
    .A2(_09256_),
    .B1(_09258_),
    .C1(_09250_),
    .X(_02522_));
 sky130_fd_sc_hd__nand2_2 _25935_ (.A(_08933_),
    .B(_09253_),
    .Y(_09259_));
 sky130_fd_sc_hd__o211a_2 _25936_ (.A1(\decode.regfile.registers_8[12] ),
    .A2(_09256_),
    .B1(_09259_),
    .C1(_09250_),
    .X(_02523_));
 sky130_fd_sc_hd__nand2_2 _25937_ (.A(_08935_),
    .B(_09253_),
    .Y(_09260_));
 sky130_fd_sc_hd__o211a_2 _25938_ (.A1(\decode.regfile.registers_8[13] ),
    .A2(_09256_),
    .B1(_09260_),
    .C1(_09250_),
    .X(_02524_));
 sky130_fd_sc_hd__nand2_2 _25939_ (.A(_08937_),
    .B(_09253_),
    .Y(_09261_));
 sky130_fd_sc_hd__o211a_2 _25940_ (.A1(\decode.regfile.registers_8[14] ),
    .A2(_09256_),
    .B1(_09261_),
    .C1(_09250_),
    .X(_02525_));
 sky130_fd_sc_hd__nand2_2 _25941_ (.A(_08939_),
    .B(_09253_),
    .Y(_09262_));
 sky130_fd_sc_hd__buf_1 _25942_ (.A(_10130_),
    .X(_09263_));
 sky130_fd_sc_hd__buf_1 _25943_ (.A(_09263_),
    .X(_09264_));
 sky130_fd_sc_hd__o211a_2 _25944_ (.A1(\decode.regfile.registers_8[15] ),
    .A2(_09256_),
    .B1(_09262_),
    .C1(_09264_),
    .X(_02526_));
 sky130_fd_sc_hd__nand2_2 _25945_ (.A(_08941_),
    .B(_09253_),
    .Y(_09265_));
 sky130_fd_sc_hd__o211a_2 _25946_ (.A1(\decode.regfile.registers_8[16] ),
    .A2(_09256_),
    .B1(_09265_),
    .C1(_09264_),
    .X(_02527_));
 sky130_fd_sc_hd__nand2_2 _25947_ (.A(_08943_),
    .B(_09253_),
    .Y(_09266_));
 sky130_fd_sc_hd__o211a_2 _25948_ (.A1(\decode.regfile.registers_8[17] ),
    .A2(_09256_),
    .B1(_09266_),
    .C1(_09264_),
    .X(_02528_));
 sky130_fd_sc_hd__buf_1 _25949_ (.A(_09241_),
    .X(_09267_));
 sky130_fd_sc_hd__nand2_2 _25950_ (.A(_08945_),
    .B(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__o211a_2 _25951_ (.A1(\decode.regfile.registers_8[18] ),
    .A2(_09256_),
    .B1(_09268_),
    .C1(_09264_),
    .X(_02529_));
 sky130_fd_sc_hd__nand2_2 _25952_ (.A(_08948_),
    .B(_09267_),
    .Y(_09269_));
 sky130_fd_sc_hd__o211a_2 _25953_ (.A1(\decode.regfile.registers_8[19] ),
    .A2(_09256_),
    .B1(_09269_),
    .C1(_09264_),
    .X(_02530_));
 sky130_fd_sc_hd__buf_1 _25954_ (.A(_09241_),
    .X(_09270_));
 sky130_fd_sc_hd__nand2_2 _25955_ (.A(_08952_),
    .B(_09267_),
    .Y(_09271_));
 sky130_fd_sc_hd__o211a_2 _25956_ (.A1(\decode.regfile.registers_8[20] ),
    .A2(_09270_),
    .B1(_09271_),
    .C1(_09264_),
    .X(_02531_));
 sky130_fd_sc_hd__nand2_2 _25957_ (.A(_08954_),
    .B(_09267_),
    .Y(_09272_));
 sky130_fd_sc_hd__o211a_2 _25958_ (.A1(\decode.regfile.registers_8[21] ),
    .A2(_09270_),
    .B1(_09272_),
    .C1(_09264_),
    .X(_02532_));
 sky130_fd_sc_hd__nand2_2 _25959_ (.A(_08956_),
    .B(_09267_),
    .Y(_09273_));
 sky130_fd_sc_hd__o211a_2 _25960_ (.A1(\decode.regfile.registers_8[22] ),
    .A2(_09270_),
    .B1(_09273_),
    .C1(_09264_),
    .X(_02533_));
 sky130_fd_sc_hd__nand2_2 _25961_ (.A(_08958_),
    .B(_09267_),
    .Y(_09274_));
 sky130_fd_sc_hd__o211a_2 _25962_ (.A1(\decode.regfile.registers_8[23] ),
    .A2(_09270_),
    .B1(_09274_),
    .C1(_09264_),
    .X(_02534_));
 sky130_fd_sc_hd__nand2_2 _25963_ (.A(_08960_),
    .B(_09267_),
    .Y(_09275_));
 sky130_fd_sc_hd__o211a_2 _25964_ (.A1(\decode.regfile.registers_8[24] ),
    .A2(_09270_),
    .B1(_09275_),
    .C1(_09264_),
    .X(_02535_));
 sky130_fd_sc_hd__nand2_2 _25965_ (.A(_08962_),
    .B(_09267_),
    .Y(_09276_));
 sky130_fd_sc_hd__buf_1 _25966_ (.A(_09263_),
    .X(_09277_));
 sky130_fd_sc_hd__o211a_2 _25967_ (.A1(\decode.regfile.registers_8[25] ),
    .A2(_09270_),
    .B1(_09276_),
    .C1(_09277_),
    .X(_02536_));
 sky130_fd_sc_hd__nand2_2 _25968_ (.A(_08964_),
    .B(_09267_),
    .Y(_09278_));
 sky130_fd_sc_hd__o211a_2 _25969_ (.A1(\decode.regfile.registers_8[26] ),
    .A2(_09270_),
    .B1(_09278_),
    .C1(_09277_),
    .X(_02537_));
 sky130_fd_sc_hd__nand2_2 _25970_ (.A(_08966_),
    .B(_09267_),
    .Y(_09279_));
 sky130_fd_sc_hd__o211a_2 _25971_ (.A1(\decode.regfile.registers_8[27] ),
    .A2(_09270_),
    .B1(_09279_),
    .C1(_09277_),
    .X(_02538_));
 sky130_fd_sc_hd__nand2_2 _25972_ (.A(_08968_),
    .B(_09241_),
    .Y(_09280_));
 sky130_fd_sc_hd__o211a_2 _25973_ (.A1(\decode.regfile.registers_8[28] ),
    .A2(_09270_),
    .B1(_09280_),
    .C1(_09277_),
    .X(_02539_));
 sky130_fd_sc_hd__nand2_2 _25974_ (.A(_08970_),
    .B(_09241_),
    .Y(_09281_));
 sky130_fd_sc_hd__o211a_2 _25975_ (.A1(\decode.regfile.registers_8[29] ),
    .A2(_09270_),
    .B1(_09281_),
    .C1(_09277_),
    .X(_02540_));
 sky130_fd_sc_hd__nand2_2 _25976_ (.A(_08973_),
    .B(_09241_),
    .Y(_09282_));
 sky130_fd_sc_hd__o211a_2 _25977_ (.A1(\decode.regfile.registers_8[30] ),
    .A2(_09243_),
    .B1(_09282_),
    .C1(_09277_),
    .X(_02541_));
 sky130_fd_sc_hd__nand2_2 _25978_ (.A(_08975_),
    .B(_09241_),
    .Y(_09283_));
 sky130_fd_sc_hd__o211a_2 _25979_ (.A1(\decode.regfile.registers_8[31] ),
    .A2(_09243_),
    .B1(_09283_),
    .C1(_09277_),
    .X(_02542_));
 sky130_fd_sc_hd__and4b_2 _25980_ (.A_N(_09930_),
    .B(_10194_),
    .C(_10240_),
    .D(_08902_),
    .X(_09284_));
 sky130_fd_sc_hd__buf_1 _25981_ (.A(_09284_),
    .X(_09285_));
 sky130_fd_sc_hd__buf_1 _25982_ (.A(_09285_),
    .X(_09286_));
 sky130_fd_sc_hd__buf_1 _25983_ (.A(_09285_),
    .X(_09287_));
 sky130_fd_sc_hd__nand2_2 _25984_ (.A(_09287_),
    .B(_09949_),
    .Y(_09288_));
 sky130_fd_sc_hd__o211a_2 _25985_ (.A1(\decode.regfile.registers_9[0] ),
    .A2(_09286_),
    .B1(_09288_),
    .C1(_09277_),
    .X(_02543_));
 sky130_fd_sc_hd__nand2_2 _25986_ (.A(_08982_),
    .B(_09287_),
    .Y(_09289_));
 sky130_fd_sc_hd__o211a_2 _25987_ (.A1(\decode.regfile.registers_9[1] ),
    .A2(_09286_),
    .B1(_09289_),
    .C1(_09277_),
    .X(_02544_));
 sky130_fd_sc_hd__nand2_2 _25988_ (.A(_08910_),
    .B(_09287_),
    .Y(_09290_));
 sky130_fd_sc_hd__o211a_2 _25989_ (.A1(\decode.regfile.registers_9[2] ),
    .A2(_09286_),
    .B1(_09290_),
    .C1(_09277_),
    .X(_02545_));
 sky130_fd_sc_hd__nand2_2 _25990_ (.A(_08912_),
    .B(_09287_),
    .Y(_09291_));
 sky130_fd_sc_hd__buf_1 _25991_ (.A(_09263_),
    .X(_09292_));
 sky130_fd_sc_hd__o211a_2 _25992_ (.A1(\decode.regfile.registers_9[3] ),
    .A2(_09286_),
    .B1(_09291_),
    .C1(_09292_),
    .X(_02546_));
 sky130_fd_sc_hd__nand2_2 _25993_ (.A(_08914_),
    .B(_09287_),
    .Y(_09293_));
 sky130_fd_sc_hd__o211a_2 _25994_ (.A1(\decode.regfile.registers_9[4] ),
    .A2(_09286_),
    .B1(_09293_),
    .C1(_09292_),
    .X(_02547_));
 sky130_fd_sc_hd__nand2_2 _25995_ (.A(_08916_),
    .B(_09287_),
    .Y(_09294_));
 sky130_fd_sc_hd__o211a_2 _25996_ (.A1(\decode.regfile.registers_9[5] ),
    .A2(_09286_),
    .B1(_09294_),
    .C1(_09292_),
    .X(_02548_));
 sky130_fd_sc_hd__nand2_2 _25997_ (.A(_08918_),
    .B(_09287_),
    .Y(_09295_));
 sky130_fd_sc_hd__o211a_2 _25998_ (.A1(\decode.regfile.registers_9[6] ),
    .A2(_09286_),
    .B1(_09295_),
    .C1(_09292_),
    .X(_02549_));
 sky130_fd_sc_hd__nand2_2 _25999_ (.A(_08920_),
    .B(_09287_),
    .Y(_09296_));
 sky130_fd_sc_hd__o211a_2 _26000_ (.A1(\decode.regfile.registers_9[7] ),
    .A2(_09286_),
    .B1(_09296_),
    .C1(_09292_),
    .X(_02550_));
 sky130_fd_sc_hd__buf_1 _26001_ (.A(_09285_),
    .X(_09297_));
 sky130_fd_sc_hd__nand2_2 _26002_ (.A(_08922_),
    .B(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__o211a_2 _26003_ (.A1(\decode.regfile.registers_9[8] ),
    .A2(_09286_),
    .B1(_09298_),
    .C1(_09292_),
    .X(_02551_));
 sky130_fd_sc_hd__nand2_2 _26004_ (.A(_08925_),
    .B(_09297_),
    .Y(_09299_));
 sky130_fd_sc_hd__o211a_2 _26005_ (.A1(\decode.regfile.registers_9[9] ),
    .A2(_09286_),
    .B1(_09299_),
    .C1(_09292_),
    .X(_02552_));
 sky130_fd_sc_hd__buf_1 _26006_ (.A(_09285_),
    .X(_09300_));
 sky130_fd_sc_hd__nand2_2 _26007_ (.A(_08929_),
    .B(_09297_),
    .Y(_09301_));
 sky130_fd_sc_hd__o211a_2 _26008_ (.A1(\decode.regfile.registers_9[10] ),
    .A2(_09300_),
    .B1(_09301_),
    .C1(_09292_),
    .X(_02553_));
 sky130_fd_sc_hd__nand2_2 _26009_ (.A(_08931_),
    .B(_09297_),
    .Y(_09302_));
 sky130_fd_sc_hd__o211a_2 _26010_ (.A1(\decode.regfile.registers_9[11] ),
    .A2(_09300_),
    .B1(_09302_),
    .C1(_09292_),
    .X(_02554_));
 sky130_fd_sc_hd__nand2_2 _26011_ (.A(_08933_),
    .B(_09297_),
    .Y(_09303_));
 sky130_fd_sc_hd__o211a_2 _26012_ (.A1(\decode.regfile.registers_9[12] ),
    .A2(_09300_),
    .B1(_09303_),
    .C1(_09292_),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_2 _26013_ (.A(_08935_),
    .B(_09297_),
    .Y(_09304_));
 sky130_fd_sc_hd__buf_1 _26014_ (.A(_09263_),
    .X(_09305_));
 sky130_fd_sc_hd__o211a_2 _26015_ (.A1(\decode.regfile.registers_9[13] ),
    .A2(_09300_),
    .B1(_09304_),
    .C1(_09305_),
    .X(_02556_));
 sky130_fd_sc_hd__nand2_2 _26016_ (.A(_08937_),
    .B(_09297_),
    .Y(_09306_));
 sky130_fd_sc_hd__o211a_2 _26017_ (.A1(\decode.regfile.registers_9[14] ),
    .A2(_09300_),
    .B1(_09306_),
    .C1(_09305_),
    .X(_02557_));
 sky130_fd_sc_hd__nand2_2 _26018_ (.A(_08939_),
    .B(_09297_),
    .Y(_09307_));
 sky130_fd_sc_hd__o211a_2 _26019_ (.A1(\decode.regfile.registers_9[15] ),
    .A2(_09300_),
    .B1(_09307_),
    .C1(_09305_),
    .X(_02558_));
 sky130_fd_sc_hd__nand2_2 _26020_ (.A(_08941_),
    .B(_09297_),
    .Y(_09308_));
 sky130_fd_sc_hd__o211a_2 _26021_ (.A1(\decode.regfile.registers_9[16] ),
    .A2(_09300_),
    .B1(_09308_),
    .C1(_09305_),
    .X(_02559_));
 sky130_fd_sc_hd__nand2_2 _26022_ (.A(_08943_),
    .B(_09297_),
    .Y(_09309_));
 sky130_fd_sc_hd__o211a_2 _26023_ (.A1(\decode.regfile.registers_9[17] ),
    .A2(_09300_),
    .B1(_09309_),
    .C1(_09305_),
    .X(_02560_));
 sky130_fd_sc_hd__buf_1 _26024_ (.A(_09285_),
    .X(_09310_));
 sky130_fd_sc_hd__nand2_2 _26025_ (.A(_08945_),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__o211a_2 _26026_ (.A1(\decode.regfile.registers_9[18] ),
    .A2(_09300_),
    .B1(_09311_),
    .C1(_09305_),
    .X(_02561_));
 sky130_fd_sc_hd__nand2_2 _26027_ (.A(_08948_),
    .B(_09310_),
    .Y(_09312_));
 sky130_fd_sc_hd__o211a_2 _26028_ (.A1(\decode.regfile.registers_9[19] ),
    .A2(_09300_),
    .B1(_09312_),
    .C1(_09305_),
    .X(_02562_));
 sky130_fd_sc_hd__buf_1 _26029_ (.A(_09285_),
    .X(_09313_));
 sky130_fd_sc_hd__nand2_2 _26030_ (.A(_08952_),
    .B(_09310_),
    .Y(_09314_));
 sky130_fd_sc_hd__o211a_2 _26031_ (.A1(\decode.regfile.registers_9[20] ),
    .A2(_09313_),
    .B1(_09314_),
    .C1(_09305_),
    .X(_02563_));
 sky130_fd_sc_hd__nand2_2 _26032_ (.A(_08954_),
    .B(_09310_),
    .Y(_09315_));
 sky130_fd_sc_hd__o211a_2 _26033_ (.A1(\decode.regfile.registers_9[21] ),
    .A2(_09313_),
    .B1(_09315_),
    .C1(_09305_),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_2 _26034_ (.A(_08956_),
    .B(_09310_),
    .Y(_09316_));
 sky130_fd_sc_hd__o211a_2 _26035_ (.A1(\decode.regfile.registers_9[22] ),
    .A2(_09313_),
    .B1(_09316_),
    .C1(_09305_),
    .X(_02565_));
 sky130_fd_sc_hd__nand2_2 _26036_ (.A(_08958_),
    .B(_09310_),
    .Y(_09317_));
 sky130_fd_sc_hd__buf_1 _26037_ (.A(_09263_),
    .X(_09318_));
 sky130_fd_sc_hd__o211a_2 _26038_ (.A1(\decode.regfile.registers_9[23] ),
    .A2(_09313_),
    .B1(_09317_),
    .C1(_09318_),
    .X(_02566_));
 sky130_fd_sc_hd__nand2_2 _26039_ (.A(_08960_),
    .B(_09310_),
    .Y(_09319_));
 sky130_fd_sc_hd__o211a_2 _26040_ (.A1(\decode.regfile.registers_9[24] ),
    .A2(_09313_),
    .B1(_09319_),
    .C1(_09318_),
    .X(_02567_));
 sky130_fd_sc_hd__nand2_2 _26041_ (.A(_08962_),
    .B(_09310_),
    .Y(_09320_));
 sky130_fd_sc_hd__o211a_2 _26042_ (.A1(\decode.regfile.registers_9[25] ),
    .A2(_09313_),
    .B1(_09320_),
    .C1(_09318_),
    .X(_02568_));
 sky130_fd_sc_hd__nand2_2 _26043_ (.A(_08964_),
    .B(_09310_),
    .Y(_09321_));
 sky130_fd_sc_hd__o211a_2 _26044_ (.A1(\decode.regfile.registers_9[26] ),
    .A2(_09313_),
    .B1(_09321_),
    .C1(_09318_),
    .X(_02569_));
 sky130_fd_sc_hd__nand2_2 _26045_ (.A(_08966_),
    .B(_09310_),
    .Y(_09322_));
 sky130_fd_sc_hd__o211a_2 _26046_ (.A1(\decode.regfile.registers_9[27] ),
    .A2(_09313_),
    .B1(_09322_),
    .C1(_09318_),
    .X(_02570_));
 sky130_fd_sc_hd__nand2_2 _26047_ (.A(_08968_),
    .B(_09285_),
    .Y(_09323_));
 sky130_fd_sc_hd__o211a_2 _26048_ (.A1(\decode.regfile.registers_9[28] ),
    .A2(_09313_),
    .B1(_09323_),
    .C1(_09318_),
    .X(_02571_));
 sky130_fd_sc_hd__nand2_2 _26049_ (.A(_08970_),
    .B(_09285_),
    .Y(_09324_));
 sky130_fd_sc_hd__o211a_2 _26050_ (.A1(\decode.regfile.registers_9[29] ),
    .A2(_09313_),
    .B1(_09324_),
    .C1(_09318_),
    .X(_02572_));
 sky130_fd_sc_hd__nand2_2 _26051_ (.A(_08973_),
    .B(_09285_),
    .Y(_09325_));
 sky130_fd_sc_hd__o211a_2 _26052_ (.A1(\decode.regfile.registers_9[30] ),
    .A2(_09287_),
    .B1(_09325_),
    .C1(_09318_),
    .X(_02573_));
 sky130_fd_sc_hd__nand2_2 _26053_ (.A(_08975_),
    .B(_09285_),
    .Y(_09326_));
 sky130_fd_sc_hd__o211a_2 _26054_ (.A1(\decode.regfile.registers_9[31] ),
    .A2(_09287_),
    .B1(_09326_),
    .C1(_09318_),
    .X(_02574_));
 sky130_fd_sc_hd__and4b_2 _26055_ (.A_N(_09930_),
    .B(_10194_),
    .C(_09932_),
    .D(_08902_),
    .X(_09327_));
 sky130_fd_sc_hd__buf_1 _26056_ (.A(_09327_),
    .X(_09328_));
 sky130_fd_sc_hd__buf_1 _26057_ (.A(_09328_),
    .X(_09329_));
 sky130_fd_sc_hd__buf_1 _26058_ (.A(_09328_),
    .X(_09330_));
 sky130_fd_sc_hd__nand2_2 _26059_ (.A(_09025_),
    .B(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__o211a_2 _26060_ (.A1(\decode.regfile.registers_10[0] ),
    .A2(_09329_),
    .B1(_09331_),
    .C1(_09318_),
    .X(_02575_));
 sky130_fd_sc_hd__nand2_2 _26061_ (.A(_08982_),
    .B(_09330_),
    .Y(_09332_));
 sky130_fd_sc_hd__buf_1 _26062_ (.A(_09263_),
    .X(_09333_));
 sky130_fd_sc_hd__o211a_2 _26063_ (.A1(\decode.regfile.registers_10[1] ),
    .A2(_09329_),
    .B1(_09332_),
    .C1(_09333_),
    .X(_02576_));
 sky130_fd_sc_hd__nand2_2 _26064_ (.A(_08910_),
    .B(_09330_),
    .Y(_09334_));
 sky130_fd_sc_hd__o211a_2 _26065_ (.A1(\decode.regfile.registers_10[2] ),
    .A2(_09329_),
    .B1(_09334_),
    .C1(_09333_),
    .X(_02577_));
 sky130_fd_sc_hd__nand2_2 _26066_ (.A(_08912_),
    .B(_09330_),
    .Y(_09335_));
 sky130_fd_sc_hd__o211a_2 _26067_ (.A1(\decode.regfile.registers_10[3] ),
    .A2(_09329_),
    .B1(_09335_),
    .C1(_09333_),
    .X(_02578_));
 sky130_fd_sc_hd__nand2_2 _26068_ (.A(_08914_),
    .B(_09330_),
    .Y(_09336_));
 sky130_fd_sc_hd__o211a_2 _26069_ (.A1(\decode.regfile.registers_10[4] ),
    .A2(_09329_),
    .B1(_09336_),
    .C1(_09333_),
    .X(_02579_));
 sky130_fd_sc_hd__nand2_2 _26070_ (.A(_08916_),
    .B(_09330_),
    .Y(_09337_));
 sky130_fd_sc_hd__o211a_2 _26071_ (.A1(\decode.regfile.registers_10[5] ),
    .A2(_09329_),
    .B1(_09337_),
    .C1(_09333_),
    .X(_02580_));
 sky130_fd_sc_hd__nand2_2 _26072_ (.A(_08918_),
    .B(_09330_),
    .Y(_09338_));
 sky130_fd_sc_hd__o211a_2 _26073_ (.A1(\decode.regfile.registers_10[6] ),
    .A2(_09329_),
    .B1(_09338_),
    .C1(_09333_),
    .X(_02581_));
 sky130_fd_sc_hd__nand2_2 _26074_ (.A(_08920_),
    .B(_09330_),
    .Y(_09339_));
 sky130_fd_sc_hd__o211a_2 _26075_ (.A1(\decode.regfile.registers_10[7] ),
    .A2(_09329_),
    .B1(_09339_),
    .C1(_09333_),
    .X(_02582_));
 sky130_fd_sc_hd__buf_1 _26076_ (.A(_09328_),
    .X(_09340_));
 sky130_fd_sc_hd__nand2_2 _26077_ (.A(_08922_),
    .B(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__o211a_2 _26078_ (.A1(\decode.regfile.registers_10[8] ),
    .A2(_09329_),
    .B1(_09341_),
    .C1(_09333_),
    .X(_02583_));
 sky130_fd_sc_hd__nand2_2 _26079_ (.A(_08925_),
    .B(_09340_),
    .Y(_09342_));
 sky130_fd_sc_hd__o211a_2 _26080_ (.A1(\decode.regfile.registers_10[9] ),
    .A2(_09329_),
    .B1(_09342_),
    .C1(_09333_),
    .X(_02584_));
 sky130_fd_sc_hd__buf_1 _26081_ (.A(_09328_),
    .X(_09343_));
 sky130_fd_sc_hd__nand2_2 _26082_ (.A(_08929_),
    .B(_09340_),
    .Y(_09344_));
 sky130_fd_sc_hd__o211a_2 _26083_ (.A1(\decode.regfile.registers_10[10] ),
    .A2(_09343_),
    .B1(_09344_),
    .C1(_09333_),
    .X(_02585_));
 sky130_fd_sc_hd__nand2_2 _26084_ (.A(_08931_),
    .B(_09340_),
    .Y(_09345_));
 sky130_fd_sc_hd__buf_1 _26085_ (.A(_09263_),
    .X(_09346_));
 sky130_fd_sc_hd__o211a_2 _26086_ (.A1(\decode.regfile.registers_10[11] ),
    .A2(_09343_),
    .B1(_09345_),
    .C1(_09346_),
    .X(_02586_));
 sky130_fd_sc_hd__nand2_2 _26087_ (.A(_08933_),
    .B(_09340_),
    .Y(_09347_));
 sky130_fd_sc_hd__o211a_2 _26088_ (.A1(\decode.regfile.registers_10[12] ),
    .A2(_09343_),
    .B1(_09347_),
    .C1(_09346_),
    .X(_02587_));
 sky130_fd_sc_hd__nand2_2 _26089_ (.A(_08935_),
    .B(_09340_),
    .Y(_09348_));
 sky130_fd_sc_hd__o211a_2 _26090_ (.A1(\decode.regfile.registers_10[13] ),
    .A2(_09343_),
    .B1(_09348_),
    .C1(_09346_),
    .X(_02588_));
 sky130_fd_sc_hd__nand2_2 _26091_ (.A(_08937_),
    .B(_09340_),
    .Y(_09349_));
 sky130_fd_sc_hd__o211a_2 _26092_ (.A1(\decode.regfile.registers_10[14] ),
    .A2(_09343_),
    .B1(_09349_),
    .C1(_09346_),
    .X(_02589_));
 sky130_fd_sc_hd__nand2_2 _26093_ (.A(_08939_),
    .B(_09340_),
    .Y(_09350_));
 sky130_fd_sc_hd__o211a_2 _26094_ (.A1(\decode.regfile.registers_10[15] ),
    .A2(_09343_),
    .B1(_09350_),
    .C1(_09346_),
    .X(_02590_));
 sky130_fd_sc_hd__nand2_2 _26095_ (.A(_08941_),
    .B(_09340_),
    .Y(_09351_));
 sky130_fd_sc_hd__o211a_2 _26096_ (.A1(\decode.regfile.registers_10[16] ),
    .A2(_09343_),
    .B1(_09351_),
    .C1(_09346_),
    .X(_02591_));
 sky130_fd_sc_hd__nand2_2 _26097_ (.A(_08943_),
    .B(_09340_),
    .Y(_09352_));
 sky130_fd_sc_hd__o211a_2 _26098_ (.A1(\decode.regfile.registers_10[17] ),
    .A2(_09343_),
    .B1(_09352_),
    .C1(_09346_),
    .X(_02592_));
 sky130_fd_sc_hd__buf_1 _26099_ (.A(_09328_),
    .X(_09353_));
 sky130_fd_sc_hd__nand2_2 _26100_ (.A(_08945_),
    .B(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__o211a_2 _26101_ (.A1(\decode.regfile.registers_10[18] ),
    .A2(_09343_),
    .B1(_09354_),
    .C1(_09346_),
    .X(_02593_));
 sky130_fd_sc_hd__nand2_2 _26102_ (.A(_08948_),
    .B(_09353_),
    .Y(_09355_));
 sky130_fd_sc_hd__o211a_2 _26103_ (.A1(\decode.regfile.registers_10[19] ),
    .A2(_09343_),
    .B1(_09355_),
    .C1(_09346_),
    .X(_02594_));
 sky130_fd_sc_hd__buf_1 _26104_ (.A(_09328_),
    .X(_09356_));
 sky130_fd_sc_hd__nand2_2 _26105_ (.A(_08952_),
    .B(_09353_),
    .Y(_09357_));
 sky130_fd_sc_hd__o211a_2 _26106_ (.A1(\decode.regfile.registers_10[20] ),
    .A2(_09356_),
    .B1(_09357_),
    .C1(_09346_),
    .X(_02595_));
 sky130_fd_sc_hd__nand2_2 _26107_ (.A(_08954_),
    .B(_09353_),
    .Y(_09358_));
 sky130_fd_sc_hd__buf_1 _26108_ (.A(_09263_),
    .X(_09359_));
 sky130_fd_sc_hd__o211a_2 _26109_ (.A1(\decode.regfile.registers_10[21] ),
    .A2(_09356_),
    .B1(_09358_),
    .C1(_09359_),
    .X(_02596_));
 sky130_fd_sc_hd__nand2_2 _26110_ (.A(_08956_),
    .B(_09353_),
    .Y(_09360_));
 sky130_fd_sc_hd__o211a_2 _26111_ (.A1(\decode.regfile.registers_10[22] ),
    .A2(_09356_),
    .B1(_09360_),
    .C1(_09359_),
    .X(_02597_));
 sky130_fd_sc_hd__nand2_2 _26112_ (.A(_08958_),
    .B(_09353_),
    .Y(_09361_));
 sky130_fd_sc_hd__o211a_2 _26113_ (.A1(\decode.regfile.registers_10[23] ),
    .A2(_09356_),
    .B1(_09361_),
    .C1(_09359_),
    .X(_02598_));
 sky130_fd_sc_hd__nand2_2 _26114_ (.A(_08960_),
    .B(_09353_),
    .Y(_09362_));
 sky130_fd_sc_hd__o211a_2 _26115_ (.A1(\decode.regfile.registers_10[24] ),
    .A2(_09356_),
    .B1(_09362_),
    .C1(_09359_),
    .X(_02599_));
 sky130_fd_sc_hd__nand2_2 _26116_ (.A(_08962_),
    .B(_09353_),
    .Y(_09363_));
 sky130_fd_sc_hd__o211a_2 _26117_ (.A1(\decode.regfile.registers_10[25] ),
    .A2(_09356_),
    .B1(_09363_),
    .C1(_09359_),
    .X(_02600_));
 sky130_fd_sc_hd__nand2_2 _26118_ (.A(_08964_),
    .B(_09353_),
    .Y(_09364_));
 sky130_fd_sc_hd__o211a_2 _26119_ (.A1(\decode.regfile.registers_10[26] ),
    .A2(_09356_),
    .B1(_09364_),
    .C1(_09359_),
    .X(_02601_));
 sky130_fd_sc_hd__nand2_2 _26120_ (.A(_08966_),
    .B(_09353_),
    .Y(_09365_));
 sky130_fd_sc_hd__o211a_2 _26121_ (.A1(\decode.regfile.registers_10[27] ),
    .A2(_09356_),
    .B1(_09365_),
    .C1(_09359_),
    .X(_02602_));
 sky130_fd_sc_hd__nand2_2 _26122_ (.A(_08968_),
    .B(_09328_),
    .Y(_09366_));
 sky130_fd_sc_hd__o211a_2 _26123_ (.A1(\decode.regfile.registers_10[28] ),
    .A2(_09356_),
    .B1(_09366_),
    .C1(_09359_),
    .X(_02603_));
 sky130_fd_sc_hd__nand2_2 _26124_ (.A(_08970_),
    .B(_09328_),
    .Y(_09367_));
 sky130_fd_sc_hd__o211a_2 _26125_ (.A1(\decode.regfile.registers_10[29] ),
    .A2(_09356_),
    .B1(_09367_),
    .C1(_09359_),
    .X(_02604_));
 sky130_fd_sc_hd__nand2_2 _26126_ (.A(_08973_),
    .B(_09328_),
    .Y(_09368_));
 sky130_fd_sc_hd__o211a_2 _26127_ (.A1(\decode.regfile.registers_10[30] ),
    .A2(_09330_),
    .B1(_09368_),
    .C1(_09359_),
    .X(_02605_));
 sky130_fd_sc_hd__nand2_2 _26128_ (.A(_08975_),
    .B(_09328_),
    .Y(_09369_));
 sky130_fd_sc_hd__buf_1 _26129_ (.A(_09263_),
    .X(_09370_));
 sky130_fd_sc_hd__o211a_2 _26130_ (.A1(\decode.regfile.registers_10[31] ),
    .A2(_09330_),
    .B1(_09369_),
    .C1(_09370_),
    .X(_02606_));
 sky130_fd_sc_hd__and4b_2 _26131_ (.A_N(_09930_),
    .B(_10194_),
    .C(_10150_),
    .D(_08902_),
    .X(_09371_));
 sky130_fd_sc_hd__buf_1 _26132_ (.A(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__buf_1 _26133_ (.A(_09372_),
    .X(_09373_));
 sky130_fd_sc_hd__buf_1 _26134_ (.A(_09372_),
    .X(_09374_));
 sky130_fd_sc_hd__nand2_2 _26135_ (.A(_09025_),
    .B(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__o211a_2 _26136_ (.A1(\decode.regfile.registers_11[0] ),
    .A2(_09373_),
    .B1(_09375_),
    .C1(_09370_),
    .X(_02607_));
 sky130_fd_sc_hd__nand2_2 _26137_ (.A(_08982_),
    .B(_09374_),
    .Y(_09376_));
 sky130_fd_sc_hd__o211a_2 _26138_ (.A1(\decode.regfile.registers_11[1] ),
    .A2(_09373_),
    .B1(_09376_),
    .C1(_09370_),
    .X(_02608_));
 sky130_fd_sc_hd__buf_1 _26139_ (.A(_09969_),
    .X(_09377_));
 sky130_fd_sc_hd__nand2_2 _26140_ (.A(_09377_),
    .B(_09374_),
    .Y(_09378_));
 sky130_fd_sc_hd__o211a_2 _26141_ (.A1(\decode.regfile.registers_11[2] ),
    .A2(_09373_),
    .B1(_09378_),
    .C1(_09370_),
    .X(_02609_));
 sky130_fd_sc_hd__buf_1 _26142_ (.A(_09974_),
    .X(_09379_));
 sky130_fd_sc_hd__nand2_2 _26143_ (.A(_09379_),
    .B(_09374_),
    .Y(_09380_));
 sky130_fd_sc_hd__o211a_2 _26144_ (.A1(\decode.regfile.registers_11[3] ),
    .A2(_09373_),
    .B1(_09380_),
    .C1(_09370_),
    .X(_02610_));
 sky130_fd_sc_hd__buf_1 _26145_ (.A(_09983_),
    .X(_09381_));
 sky130_fd_sc_hd__nand2_2 _26146_ (.A(_09381_),
    .B(_09374_),
    .Y(_09382_));
 sky130_fd_sc_hd__o211a_2 _26147_ (.A1(\decode.regfile.registers_11[4] ),
    .A2(_09373_),
    .B1(_09382_),
    .C1(_09370_),
    .X(_02611_));
 sky130_fd_sc_hd__buf_1 _26148_ (.A(_09992_),
    .X(_09383_));
 sky130_fd_sc_hd__nand2_2 _26149_ (.A(_09383_),
    .B(_09374_),
    .Y(_09384_));
 sky130_fd_sc_hd__o211a_2 _26150_ (.A1(\decode.regfile.registers_11[5] ),
    .A2(_09373_),
    .B1(_09384_),
    .C1(_09370_),
    .X(_02612_));
 sky130_fd_sc_hd__buf_1 _26151_ (.A(_09998_),
    .X(_09385_));
 sky130_fd_sc_hd__nand2_2 _26152_ (.A(_09385_),
    .B(_09374_),
    .Y(_09386_));
 sky130_fd_sc_hd__o211a_2 _26153_ (.A1(\decode.regfile.registers_11[6] ),
    .A2(_09373_),
    .B1(_09386_),
    .C1(_09370_),
    .X(_02613_));
 sky130_fd_sc_hd__buf_1 _26154_ (.A(_10007_),
    .X(_09387_));
 sky130_fd_sc_hd__nand2_2 _26155_ (.A(_09387_),
    .B(_09374_),
    .Y(_09388_));
 sky130_fd_sc_hd__o211a_2 _26156_ (.A1(\decode.regfile.registers_11[7] ),
    .A2(_09373_),
    .B1(_09388_),
    .C1(_09370_),
    .X(_02614_));
 sky130_fd_sc_hd__buf_1 _26157_ (.A(_10014_),
    .X(_09389_));
 sky130_fd_sc_hd__buf_1 _26158_ (.A(_09372_),
    .X(_09390_));
 sky130_fd_sc_hd__nand2_2 _26159_ (.A(_09389_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__o211a_2 _26160_ (.A1(\decode.regfile.registers_11[8] ),
    .A2(_09373_),
    .B1(_09391_),
    .C1(_09370_),
    .X(_02615_));
 sky130_fd_sc_hd__buf_1 _26161_ (.A(_10024_),
    .X(_09392_));
 sky130_fd_sc_hd__nand2_2 _26162_ (.A(_09392_),
    .B(_09390_),
    .Y(_09393_));
 sky130_fd_sc_hd__buf_1 _26163_ (.A(_09263_),
    .X(_09394_));
 sky130_fd_sc_hd__o211a_2 _26164_ (.A1(\decode.regfile.registers_11[9] ),
    .A2(_09373_),
    .B1(_09393_),
    .C1(_09394_),
    .X(_02616_));
 sky130_fd_sc_hd__buf_1 _26165_ (.A(_09372_),
    .X(_09395_));
 sky130_fd_sc_hd__buf_1 _26166_ (.A(_10030_),
    .X(_09396_));
 sky130_fd_sc_hd__nand2_2 _26167_ (.A(_09396_),
    .B(_09390_),
    .Y(_09397_));
 sky130_fd_sc_hd__o211a_2 _26168_ (.A1(\decode.regfile.registers_11[10] ),
    .A2(_09395_),
    .B1(_09397_),
    .C1(_09394_),
    .X(_02617_));
 sky130_fd_sc_hd__buf_1 _26169_ (.A(_10035_),
    .X(_09398_));
 sky130_fd_sc_hd__nand2_2 _26170_ (.A(_09398_),
    .B(_09390_),
    .Y(_09399_));
 sky130_fd_sc_hd__o211a_2 _26171_ (.A1(\decode.regfile.registers_11[11] ),
    .A2(_09395_),
    .B1(_09399_),
    .C1(_09394_),
    .X(_02618_));
 sky130_fd_sc_hd__buf_1 _26172_ (.A(_10041_),
    .X(_09400_));
 sky130_fd_sc_hd__nand2_2 _26173_ (.A(_09400_),
    .B(_09390_),
    .Y(_09401_));
 sky130_fd_sc_hd__o211a_2 _26174_ (.A1(\decode.regfile.registers_11[12] ),
    .A2(_09395_),
    .B1(_09401_),
    .C1(_09394_),
    .X(_02619_));
 sky130_fd_sc_hd__buf_1 _26175_ (.A(_10047_),
    .X(_09402_));
 sky130_fd_sc_hd__nand2_2 _26176_ (.A(_09402_),
    .B(_09390_),
    .Y(_09403_));
 sky130_fd_sc_hd__o211a_2 _26177_ (.A1(\decode.regfile.registers_11[13] ),
    .A2(_09395_),
    .B1(_09403_),
    .C1(_09394_),
    .X(_02620_));
 sky130_fd_sc_hd__buf_1 _26178_ (.A(_10052_),
    .X(_09404_));
 sky130_fd_sc_hd__nand2_2 _26179_ (.A(_09404_),
    .B(_09390_),
    .Y(_09405_));
 sky130_fd_sc_hd__o211a_2 _26180_ (.A1(\decode.regfile.registers_11[14] ),
    .A2(_09395_),
    .B1(_09405_),
    .C1(_09394_),
    .X(_02621_));
 sky130_fd_sc_hd__buf_1 _26181_ (.A(_10057_),
    .X(_09406_));
 sky130_fd_sc_hd__nand2_2 _26182_ (.A(_09406_),
    .B(_09390_),
    .Y(_09407_));
 sky130_fd_sc_hd__o211a_2 _26183_ (.A1(\decode.regfile.registers_11[15] ),
    .A2(_09395_),
    .B1(_09407_),
    .C1(_09394_),
    .X(_02622_));
 sky130_fd_sc_hd__buf_1 _26184_ (.A(_10063_),
    .X(_09408_));
 sky130_fd_sc_hd__nand2_2 _26185_ (.A(_09408_),
    .B(_09390_),
    .Y(_09409_));
 sky130_fd_sc_hd__o211a_2 _26186_ (.A1(\decode.regfile.registers_11[16] ),
    .A2(_09395_),
    .B1(_09409_),
    .C1(_09394_),
    .X(_02623_));
 sky130_fd_sc_hd__buf_1 _26187_ (.A(_10068_),
    .X(_09410_));
 sky130_fd_sc_hd__nand2_2 _26188_ (.A(_09410_),
    .B(_09390_),
    .Y(_09411_));
 sky130_fd_sc_hd__o211a_2 _26189_ (.A1(\decode.regfile.registers_11[17] ),
    .A2(_09395_),
    .B1(_09411_),
    .C1(_09394_),
    .X(_02624_));
 sky130_fd_sc_hd__buf_1 _26190_ (.A(_10073_),
    .X(_09412_));
 sky130_fd_sc_hd__buf_1 _26191_ (.A(_09372_),
    .X(_09413_));
 sky130_fd_sc_hd__nand2_2 _26192_ (.A(_09412_),
    .B(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__o211a_2 _26193_ (.A1(\decode.regfile.registers_11[18] ),
    .A2(_09395_),
    .B1(_09414_),
    .C1(_09394_),
    .X(_02625_));
 sky130_fd_sc_hd__buf_1 _26194_ (.A(_10080_),
    .X(_09415_));
 sky130_fd_sc_hd__nand2_2 _26195_ (.A(_09415_),
    .B(_09413_),
    .Y(_09416_));
 sky130_fd_sc_hd__buf_1 _26196_ (.A(_10130_),
    .X(_09417_));
 sky130_fd_sc_hd__buf_1 _26197_ (.A(_09417_),
    .X(_09418_));
 sky130_fd_sc_hd__o211a_2 _26198_ (.A1(\decode.regfile.registers_11[19] ),
    .A2(_09395_),
    .B1(_09416_),
    .C1(_09418_),
    .X(_02626_));
 sky130_fd_sc_hd__buf_1 _26199_ (.A(_09372_),
    .X(_09419_));
 sky130_fd_sc_hd__buf_1 _26200_ (.A(_10086_),
    .X(_09420_));
 sky130_fd_sc_hd__nand2_2 _26201_ (.A(_09420_),
    .B(_09413_),
    .Y(_09421_));
 sky130_fd_sc_hd__o211a_2 _26202_ (.A1(\decode.regfile.registers_11[20] ),
    .A2(_09419_),
    .B1(_09421_),
    .C1(_09418_),
    .X(_02627_));
 sky130_fd_sc_hd__buf_1 _26203_ (.A(_10091_),
    .X(_09422_));
 sky130_fd_sc_hd__nand2_2 _26204_ (.A(_09422_),
    .B(_09413_),
    .Y(_09423_));
 sky130_fd_sc_hd__o211a_2 _26205_ (.A1(\decode.regfile.registers_11[21] ),
    .A2(_09419_),
    .B1(_09423_),
    .C1(_09418_),
    .X(_02628_));
 sky130_fd_sc_hd__buf_1 _26206_ (.A(_10096_),
    .X(_09424_));
 sky130_fd_sc_hd__nand2_2 _26207_ (.A(_09424_),
    .B(_09413_),
    .Y(_09425_));
 sky130_fd_sc_hd__o211a_2 _26208_ (.A1(\decode.regfile.registers_11[22] ),
    .A2(_09419_),
    .B1(_09425_),
    .C1(_09418_),
    .X(_02629_));
 sky130_fd_sc_hd__buf_1 _26209_ (.A(_10101_),
    .X(_09426_));
 sky130_fd_sc_hd__nand2_2 _26210_ (.A(_09426_),
    .B(_09413_),
    .Y(_09427_));
 sky130_fd_sc_hd__o211a_2 _26211_ (.A1(\decode.regfile.registers_11[23] ),
    .A2(_09419_),
    .B1(_09427_),
    .C1(_09418_),
    .X(_02630_));
 sky130_fd_sc_hd__buf_1 _26212_ (.A(_10106_),
    .X(_09428_));
 sky130_fd_sc_hd__nand2_2 _26213_ (.A(_09428_),
    .B(_09413_),
    .Y(_09429_));
 sky130_fd_sc_hd__o211a_2 _26214_ (.A1(\decode.regfile.registers_11[24] ),
    .A2(_09419_),
    .B1(_09429_),
    .C1(_09418_),
    .X(_02631_));
 sky130_fd_sc_hd__buf_1 _26215_ (.A(_10111_),
    .X(_09430_));
 sky130_fd_sc_hd__nand2_2 _26216_ (.A(_09430_),
    .B(_09413_),
    .Y(_09431_));
 sky130_fd_sc_hd__o211a_2 _26217_ (.A1(\decode.regfile.registers_11[25] ),
    .A2(_09419_),
    .B1(_09431_),
    .C1(_09418_),
    .X(_02632_));
 sky130_fd_sc_hd__buf_1 _26218_ (.A(_10116_),
    .X(_09432_));
 sky130_fd_sc_hd__nand2_2 _26219_ (.A(_09432_),
    .B(_09413_),
    .Y(_09433_));
 sky130_fd_sc_hd__o211a_2 _26220_ (.A1(\decode.regfile.registers_11[26] ),
    .A2(_09419_),
    .B1(_09433_),
    .C1(_09418_),
    .X(_02633_));
 sky130_fd_sc_hd__buf_1 _26221_ (.A(_10121_),
    .X(_09434_));
 sky130_fd_sc_hd__nand2_2 _26222_ (.A(_09434_),
    .B(_09413_),
    .Y(_09435_));
 sky130_fd_sc_hd__o211a_2 _26223_ (.A1(\decode.regfile.registers_11[27] ),
    .A2(_09419_),
    .B1(_09435_),
    .C1(_09418_),
    .X(_02634_));
 sky130_fd_sc_hd__buf_1 _26224_ (.A(_10127_),
    .X(_09436_));
 sky130_fd_sc_hd__nand2_2 _26225_ (.A(_09436_),
    .B(_09372_),
    .Y(_09437_));
 sky130_fd_sc_hd__o211a_2 _26226_ (.A1(\decode.regfile.registers_11[28] ),
    .A2(_09419_),
    .B1(_09437_),
    .C1(_09418_),
    .X(_02635_));
 sky130_fd_sc_hd__buf_1 _26227_ (.A(_10135_),
    .X(_09438_));
 sky130_fd_sc_hd__nand2_2 _26228_ (.A(_09438_),
    .B(_09372_),
    .Y(_09439_));
 sky130_fd_sc_hd__buf_1 _26229_ (.A(_09417_),
    .X(_09440_));
 sky130_fd_sc_hd__o211a_2 _26230_ (.A1(\decode.regfile.registers_11[29] ),
    .A2(_09419_),
    .B1(_09439_),
    .C1(_09440_),
    .X(_02636_));
 sky130_fd_sc_hd__buf_1 _26231_ (.A(_10141_),
    .X(_09441_));
 sky130_fd_sc_hd__nand2_2 _26232_ (.A(_09441_),
    .B(_09372_),
    .Y(_09442_));
 sky130_fd_sc_hd__o211a_2 _26233_ (.A1(\decode.regfile.registers_11[30] ),
    .A2(_09374_),
    .B1(_09442_),
    .C1(_09440_),
    .X(_02637_));
 sky130_fd_sc_hd__buf_1 _26234_ (.A(_10146_),
    .X(_09443_));
 sky130_fd_sc_hd__nand2_2 _26235_ (.A(_09443_),
    .B(_09372_),
    .Y(_09444_));
 sky130_fd_sc_hd__o211a_2 _26236_ (.A1(\decode.regfile.registers_11[31] ),
    .A2(_09374_),
    .B1(_09444_),
    .C1(_09440_),
    .X(_02638_));
 sky130_fd_sc_hd__and4_2 _26237_ (.A(_10373_),
    .B(_10195_),
    .C(_10196_),
    .D(_08903_),
    .X(_09445_));
 sky130_fd_sc_hd__buf_1 _26238_ (.A(_09445_),
    .X(_09446_));
 sky130_fd_sc_hd__buf_1 _26239_ (.A(_09446_),
    .X(_09447_));
 sky130_fd_sc_hd__buf_1 _26240_ (.A(_09446_),
    .X(_09448_));
 sky130_fd_sc_hd__nand2_2 _26241_ (.A(_09025_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__o211a_2 _26242_ (.A1(\decode.regfile.registers_12[0] ),
    .A2(_09447_),
    .B1(_09449_),
    .C1(_09440_),
    .X(_02639_));
 sky130_fd_sc_hd__buf_1 _26243_ (.A(_09963_),
    .X(_09450_));
 sky130_fd_sc_hd__nand2_2 _26244_ (.A(_09450_),
    .B(_09448_),
    .Y(_09451_));
 sky130_fd_sc_hd__o211a_2 _26245_ (.A1(\decode.regfile.registers_12[1] ),
    .A2(_09447_),
    .B1(_09451_),
    .C1(_09440_),
    .X(_02640_));
 sky130_fd_sc_hd__nand2_2 _26246_ (.A(_09377_),
    .B(_09448_),
    .Y(_09452_));
 sky130_fd_sc_hd__o211a_2 _26247_ (.A1(\decode.regfile.registers_12[2] ),
    .A2(_09447_),
    .B1(_09452_),
    .C1(_09440_),
    .X(_02641_));
 sky130_fd_sc_hd__nand2_2 _26248_ (.A(_09379_),
    .B(_09448_),
    .Y(_09453_));
 sky130_fd_sc_hd__o211a_2 _26249_ (.A1(\decode.regfile.registers_12[3] ),
    .A2(_09447_),
    .B1(_09453_),
    .C1(_09440_),
    .X(_02642_));
 sky130_fd_sc_hd__nand2_2 _26250_ (.A(_09381_),
    .B(_09448_),
    .Y(_09454_));
 sky130_fd_sc_hd__o211a_2 _26251_ (.A1(\decode.regfile.registers_12[4] ),
    .A2(_09447_),
    .B1(_09454_),
    .C1(_09440_),
    .X(_02643_));
 sky130_fd_sc_hd__nand2_2 _26252_ (.A(_09383_),
    .B(_09448_),
    .Y(_09455_));
 sky130_fd_sc_hd__o211a_2 _26253_ (.A1(\decode.regfile.registers_12[5] ),
    .A2(_09447_),
    .B1(_09455_),
    .C1(_09440_),
    .X(_02644_));
 sky130_fd_sc_hd__nand2_2 _26254_ (.A(_09385_),
    .B(_09448_),
    .Y(_09456_));
 sky130_fd_sc_hd__o211a_2 _26255_ (.A1(\decode.regfile.registers_12[6] ),
    .A2(_09447_),
    .B1(_09456_),
    .C1(_09440_),
    .X(_02645_));
 sky130_fd_sc_hd__nand2_2 _26256_ (.A(_09387_),
    .B(_09448_),
    .Y(_09457_));
 sky130_fd_sc_hd__buf_1 _26257_ (.A(_09417_),
    .X(_09458_));
 sky130_fd_sc_hd__o211a_2 _26258_ (.A1(\decode.regfile.registers_12[7] ),
    .A2(_09447_),
    .B1(_09457_),
    .C1(_09458_),
    .X(_02646_));
 sky130_fd_sc_hd__buf_1 _26259_ (.A(_09446_),
    .X(_09459_));
 sky130_fd_sc_hd__nand2_2 _26260_ (.A(_09389_),
    .B(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__o211a_2 _26261_ (.A1(\decode.regfile.registers_12[8] ),
    .A2(_09447_),
    .B1(_09460_),
    .C1(_09458_),
    .X(_02647_));
 sky130_fd_sc_hd__nand2_2 _26262_ (.A(_09392_),
    .B(_09459_),
    .Y(_09461_));
 sky130_fd_sc_hd__o211a_2 _26263_ (.A1(\decode.regfile.registers_12[9] ),
    .A2(_09447_),
    .B1(_09461_),
    .C1(_09458_),
    .X(_02648_));
 sky130_fd_sc_hd__buf_1 _26264_ (.A(_09446_),
    .X(_09462_));
 sky130_fd_sc_hd__nand2_2 _26265_ (.A(_09396_),
    .B(_09459_),
    .Y(_09463_));
 sky130_fd_sc_hd__o211a_2 _26266_ (.A1(\decode.regfile.registers_12[10] ),
    .A2(_09462_),
    .B1(_09463_),
    .C1(_09458_),
    .X(_02649_));
 sky130_fd_sc_hd__nand2_2 _26267_ (.A(_09398_),
    .B(_09459_),
    .Y(_09464_));
 sky130_fd_sc_hd__o211a_2 _26268_ (.A1(\decode.regfile.registers_12[11] ),
    .A2(_09462_),
    .B1(_09464_),
    .C1(_09458_),
    .X(_02650_));
 sky130_fd_sc_hd__nand2_2 _26269_ (.A(_09400_),
    .B(_09459_),
    .Y(_09465_));
 sky130_fd_sc_hd__o211a_2 _26270_ (.A1(\decode.regfile.registers_12[12] ),
    .A2(_09462_),
    .B1(_09465_),
    .C1(_09458_),
    .X(_02651_));
 sky130_fd_sc_hd__nand2_2 _26271_ (.A(_09402_),
    .B(_09459_),
    .Y(_09466_));
 sky130_fd_sc_hd__o211a_2 _26272_ (.A1(\decode.regfile.registers_12[13] ),
    .A2(_09462_),
    .B1(_09466_),
    .C1(_09458_),
    .X(_02652_));
 sky130_fd_sc_hd__nand2_2 _26273_ (.A(_09404_),
    .B(_09459_),
    .Y(_09467_));
 sky130_fd_sc_hd__o211a_2 _26274_ (.A1(\decode.regfile.registers_12[14] ),
    .A2(_09462_),
    .B1(_09467_),
    .C1(_09458_),
    .X(_02653_));
 sky130_fd_sc_hd__nand2_2 _26275_ (.A(_09406_),
    .B(_09459_),
    .Y(_09468_));
 sky130_fd_sc_hd__o211a_2 _26276_ (.A1(\decode.regfile.registers_12[15] ),
    .A2(_09462_),
    .B1(_09468_),
    .C1(_09458_),
    .X(_02654_));
 sky130_fd_sc_hd__nand2_2 _26277_ (.A(_09408_),
    .B(_09459_),
    .Y(_09469_));
 sky130_fd_sc_hd__o211a_2 _26278_ (.A1(\decode.regfile.registers_12[16] ),
    .A2(_09462_),
    .B1(_09469_),
    .C1(_09458_),
    .X(_02655_));
 sky130_fd_sc_hd__nand2_2 _26279_ (.A(_09410_),
    .B(_09459_),
    .Y(_09470_));
 sky130_fd_sc_hd__buf_1 _26280_ (.A(_09417_),
    .X(_09471_));
 sky130_fd_sc_hd__o211a_2 _26281_ (.A1(\decode.regfile.registers_12[17] ),
    .A2(_09462_),
    .B1(_09470_),
    .C1(_09471_),
    .X(_02656_));
 sky130_fd_sc_hd__buf_1 _26282_ (.A(_09446_),
    .X(_09472_));
 sky130_fd_sc_hd__nand2_2 _26283_ (.A(_09412_),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__o211a_2 _26284_ (.A1(\decode.regfile.registers_12[18] ),
    .A2(_09462_),
    .B1(_09473_),
    .C1(_09471_),
    .X(_02657_));
 sky130_fd_sc_hd__nand2_2 _26285_ (.A(_09415_),
    .B(_09472_),
    .Y(_09474_));
 sky130_fd_sc_hd__o211a_2 _26286_ (.A1(\decode.regfile.registers_12[19] ),
    .A2(_09462_),
    .B1(_09474_),
    .C1(_09471_),
    .X(_02658_));
 sky130_fd_sc_hd__buf_1 _26287_ (.A(_09446_),
    .X(_09475_));
 sky130_fd_sc_hd__nand2_2 _26288_ (.A(_09420_),
    .B(_09472_),
    .Y(_09476_));
 sky130_fd_sc_hd__o211a_2 _26289_ (.A1(\decode.regfile.registers_12[20] ),
    .A2(_09475_),
    .B1(_09476_),
    .C1(_09471_),
    .X(_02659_));
 sky130_fd_sc_hd__nand2_2 _26290_ (.A(_09422_),
    .B(_09472_),
    .Y(_09477_));
 sky130_fd_sc_hd__o211a_2 _26291_ (.A1(\decode.regfile.registers_12[21] ),
    .A2(_09475_),
    .B1(_09477_),
    .C1(_09471_),
    .X(_02660_));
 sky130_fd_sc_hd__nand2_2 _26292_ (.A(_09424_),
    .B(_09472_),
    .Y(_09478_));
 sky130_fd_sc_hd__o211a_2 _26293_ (.A1(\decode.regfile.registers_12[22] ),
    .A2(_09475_),
    .B1(_09478_),
    .C1(_09471_),
    .X(_02661_));
 sky130_fd_sc_hd__nand2_2 _26294_ (.A(_09426_),
    .B(_09472_),
    .Y(_09479_));
 sky130_fd_sc_hd__o211a_2 _26295_ (.A1(\decode.regfile.registers_12[23] ),
    .A2(_09475_),
    .B1(_09479_),
    .C1(_09471_),
    .X(_02662_));
 sky130_fd_sc_hd__nand2_2 _26296_ (.A(_09428_),
    .B(_09472_),
    .Y(_09480_));
 sky130_fd_sc_hd__o211a_2 _26297_ (.A1(\decode.regfile.registers_12[24] ),
    .A2(_09475_),
    .B1(_09480_),
    .C1(_09471_),
    .X(_02663_));
 sky130_fd_sc_hd__nand2_2 _26298_ (.A(_09430_),
    .B(_09472_),
    .Y(_09481_));
 sky130_fd_sc_hd__o211a_2 _26299_ (.A1(\decode.regfile.registers_12[25] ),
    .A2(_09475_),
    .B1(_09481_),
    .C1(_09471_),
    .X(_02664_));
 sky130_fd_sc_hd__nand2_2 _26300_ (.A(_09432_),
    .B(_09472_),
    .Y(_09482_));
 sky130_fd_sc_hd__o211a_2 _26301_ (.A1(\decode.regfile.registers_12[26] ),
    .A2(_09475_),
    .B1(_09482_),
    .C1(_09471_),
    .X(_02665_));
 sky130_fd_sc_hd__nand2_2 _26302_ (.A(_09434_),
    .B(_09472_),
    .Y(_09483_));
 sky130_fd_sc_hd__buf_1 _26303_ (.A(_09417_),
    .X(_09484_));
 sky130_fd_sc_hd__o211a_2 _26304_ (.A1(\decode.regfile.registers_12[27] ),
    .A2(_09475_),
    .B1(_09483_),
    .C1(_09484_),
    .X(_02666_));
 sky130_fd_sc_hd__nand2_2 _26305_ (.A(_09436_),
    .B(_09446_),
    .Y(_09485_));
 sky130_fd_sc_hd__o211a_2 _26306_ (.A1(\decode.regfile.registers_12[28] ),
    .A2(_09475_),
    .B1(_09485_),
    .C1(_09484_),
    .X(_02667_));
 sky130_fd_sc_hd__nand2_2 _26307_ (.A(_09438_),
    .B(_09446_),
    .Y(_09486_));
 sky130_fd_sc_hd__o211a_2 _26308_ (.A1(\decode.regfile.registers_12[29] ),
    .A2(_09475_),
    .B1(_09486_),
    .C1(_09484_),
    .X(_02668_));
 sky130_fd_sc_hd__nand2_2 _26309_ (.A(_09441_),
    .B(_09446_),
    .Y(_09487_));
 sky130_fd_sc_hd__o211a_2 _26310_ (.A1(\decode.regfile.registers_12[30] ),
    .A2(_09448_),
    .B1(_09487_),
    .C1(_09484_),
    .X(_02669_));
 sky130_fd_sc_hd__nand2_2 _26311_ (.A(_09443_),
    .B(_09446_),
    .Y(_09488_));
 sky130_fd_sc_hd__o211a_2 _26312_ (.A1(\decode.regfile.registers_12[31] ),
    .A2(_09448_),
    .B1(_09488_),
    .C1(_09484_),
    .X(_02670_));
 sky130_fd_sc_hd__and4_2 _26313_ (.A(_10373_),
    .B(_10195_),
    .C(_10240_),
    .D(_08903_),
    .X(_09489_));
 sky130_fd_sc_hd__buf_1 _26314_ (.A(_09489_),
    .X(_09490_));
 sky130_fd_sc_hd__buf_1 _26315_ (.A(_09490_),
    .X(_09491_));
 sky130_fd_sc_hd__buf_1 _26316_ (.A(_09490_),
    .X(_09492_));
 sky130_fd_sc_hd__nand2_2 _26317_ (.A(_09025_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__o211a_2 _26318_ (.A1(\decode.regfile.registers_13[0] ),
    .A2(_09491_),
    .B1(_09493_),
    .C1(_09484_),
    .X(_02671_));
 sky130_fd_sc_hd__nand2_2 _26319_ (.A(_09450_),
    .B(_09492_),
    .Y(_09494_));
 sky130_fd_sc_hd__o211a_2 _26320_ (.A1(\decode.regfile.registers_13[1] ),
    .A2(_09491_),
    .B1(_09494_),
    .C1(_09484_),
    .X(_02672_));
 sky130_fd_sc_hd__nand2_2 _26321_ (.A(_09377_),
    .B(_09492_),
    .Y(_09495_));
 sky130_fd_sc_hd__o211a_2 _26322_ (.A1(\decode.regfile.registers_13[2] ),
    .A2(_09491_),
    .B1(_09495_),
    .C1(_09484_),
    .X(_02673_));
 sky130_fd_sc_hd__nand2_2 _26323_ (.A(_09379_),
    .B(_09492_),
    .Y(_09496_));
 sky130_fd_sc_hd__o211a_2 _26324_ (.A1(\decode.regfile.registers_13[3] ),
    .A2(_09491_),
    .B1(_09496_),
    .C1(_09484_),
    .X(_02674_));
 sky130_fd_sc_hd__nand2_2 _26325_ (.A(_09381_),
    .B(_09492_),
    .Y(_09497_));
 sky130_fd_sc_hd__o211a_2 _26326_ (.A1(\decode.regfile.registers_13[4] ),
    .A2(_09491_),
    .B1(_09497_),
    .C1(_09484_),
    .X(_02675_));
 sky130_fd_sc_hd__nand2_2 _26327_ (.A(_09383_),
    .B(_09492_),
    .Y(_09498_));
 sky130_fd_sc_hd__buf_1 _26328_ (.A(_09417_),
    .X(_09499_));
 sky130_fd_sc_hd__o211a_2 _26329_ (.A1(\decode.regfile.registers_13[5] ),
    .A2(_09491_),
    .B1(_09498_),
    .C1(_09499_),
    .X(_02676_));
 sky130_fd_sc_hd__nand2_2 _26330_ (.A(_09385_),
    .B(_09492_),
    .Y(_09500_));
 sky130_fd_sc_hd__o211a_2 _26331_ (.A1(\decode.regfile.registers_13[6] ),
    .A2(_09491_),
    .B1(_09500_),
    .C1(_09499_),
    .X(_02677_));
 sky130_fd_sc_hd__nand2_2 _26332_ (.A(_09387_),
    .B(_09492_),
    .Y(_09501_));
 sky130_fd_sc_hd__o211a_2 _26333_ (.A1(\decode.regfile.registers_13[7] ),
    .A2(_09491_),
    .B1(_09501_),
    .C1(_09499_),
    .X(_02678_));
 sky130_fd_sc_hd__buf_1 _26334_ (.A(_09490_),
    .X(_09502_));
 sky130_fd_sc_hd__nand2_2 _26335_ (.A(_09389_),
    .B(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__o211a_2 _26336_ (.A1(\decode.regfile.registers_13[8] ),
    .A2(_09491_),
    .B1(_09503_),
    .C1(_09499_),
    .X(_02679_));
 sky130_fd_sc_hd__nand2_2 _26337_ (.A(_09392_),
    .B(_09502_),
    .Y(_09504_));
 sky130_fd_sc_hd__o211a_2 _26338_ (.A1(\decode.regfile.registers_13[9] ),
    .A2(_09491_),
    .B1(_09504_),
    .C1(_09499_),
    .X(_02680_));
 sky130_fd_sc_hd__buf_1 _26339_ (.A(_09490_),
    .X(_09505_));
 sky130_fd_sc_hd__nand2_2 _26340_ (.A(_09396_),
    .B(_09502_),
    .Y(_09506_));
 sky130_fd_sc_hd__o211a_2 _26341_ (.A1(\decode.regfile.registers_13[10] ),
    .A2(_09505_),
    .B1(_09506_),
    .C1(_09499_),
    .X(_02681_));
 sky130_fd_sc_hd__nand2_2 _26342_ (.A(_09398_),
    .B(_09502_),
    .Y(_09507_));
 sky130_fd_sc_hd__o211a_2 _26343_ (.A1(\decode.regfile.registers_13[11] ),
    .A2(_09505_),
    .B1(_09507_),
    .C1(_09499_),
    .X(_02682_));
 sky130_fd_sc_hd__nand2_2 _26344_ (.A(_09400_),
    .B(_09502_),
    .Y(_09508_));
 sky130_fd_sc_hd__o211a_2 _26345_ (.A1(\decode.regfile.registers_13[12] ),
    .A2(_09505_),
    .B1(_09508_),
    .C1(_09499_),
    .X(_02683_));
 sky130_fd_sc_hd__nand2_2 _26346_ (.A(_09402_),
    .B(_09502_),
    .Y(_09509_));
 sky130_fd_sc_hd__o211a_2 _26347_ (.A1(\decode.regfile.registers_13[13] ),
    .A2(_09505_),
    .B1(_09509_),
    .C1(_09499_),
    .X(_02684_));
 sky130_fd_sc_hd__nand2_2 _26348_ (.A(_09404_),
    .B(_09502_),
    .Y(_09510_));
 sky130_fd_sc_hd__o211a_2 _26349_ (.A1(\decode.regfile.registers_13[14] ),
    .A2(_09505_),
    .B1(_09510_),
    .C1(_09499_),
    .X(_02685_));
 sky130_fd_sc_hd__nand2_2 _26350_ (.A(_09406_),
    .B(_09502_),
    .Y(_09511_));
 sky130_fd_sc_hd__buf_1 _26351_ (.A(_09417_),
    .X(_09512_));
 sky130_fd_sc_hd__o211a_2 _26352_ (.A1(\decode.regfile.registers_13[15] ),
    .A2(_09505_),
    .B1(_09511_),
    .C1(_09512_),
    .X(_02686_));
 sky130_fd_sc_hd__nand2_2 _26353_ (.A(_09408_),
    .B(_09502_),
    .Y(_09513_));
 sky130_fd_sc_hd__o211a_2 _26354_ (.A1(\decode.regfile.registers_13[16] ),
    .A2(_09505_),
    .B1(_09513_),
    .C1(_09512_),
    .X(_02687_));
 sky130_fd_sc_hd__nand2_2 _26355_ (.A(_09410_),
    .B(_09502_),
    .Y(_09514_));
 sky130_fd_sc_hd__o211a_2 _26356_ (.A1(\decode.regfile.registers_13[17] ),
    .A2(_09505_),
    .B1(_09514_),
    .C1(_09512_),
    .X(_02688_));
 sky130_fd_sc_hd__buf_1 _26357_ (.A(_09490_),
    .X(_09515_));
 sky130_fd_sc_hd__nand2_2 _26358_ (.A(_09412_),
    .B(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__o211a_2 _26359_ (.A1(\decode.regfile.registers_13[18] ),
    .A2(_09505_),
    .B1(_09516_),
    .C1(_09512_),
    .X(_02689_));
 sky130_fd_sc_hd__nand2_2 _26360_ (.A(_09415_),
    .B(_09515_),
    .Y(_09517_));
 sky130_fd_sc_hd__o211a_2 _26361_ (.A1(\decode.regfile.registers_13[19] ),
    .A2(_09505_),
    .B1(_09517_),
    .C1(_09512_),
    .X(_02690_));
 sky130_fd_sc_hd__buf_1 _26362_ (.A(_09490_),
    .X(_09518_));
 sky130_fd_sc_hd__nand2_2 _26363_ (.A(_09420_),
    .B(_09515_),
    .Y(_09519_));
 sky130_fd_sc_hd__o211a_2 _26364_ (.A1(\decode.regfile.registers_13[20] ),
    .A2(_09518_),
    .B1(_09519_),
    .C1(_09512_),
    .X(_02691_));
 sky130_fd_sc_hd__nand2_2 _26365_ (.A(_09422_),
    .B(_09515_),
    .Y(_09520_));
 sky130_fd_sc_hd__o211a_2 _26366_ (.A1(\decode.regfile.registers_13[21] ),
    .A2(_09518_),
    .B1(_09520_),
    .C1(_09512_),
    .X(_02692_));
 sky130_fd_sc_hd__nand2_2 _26367_ (.A(_09424_),
    .B(_09515_),
    .Y(_09521_));
 sky130_fd_sc_hd__o211a_2 _26368_ (.A1(\decode.regfile.registers_13[22] ),
    .A2(_09518_),
    .B1(_09521_),
    .C1(_09512_),
    .X(_02693_));
 sky130_fd_sc_hd__nand2_2 _26369_ (.A(_09426_),
    .B(_09515_),
    .Y(_09522_));
 sky130_fd_sc_hd__o211a_2 _26370_ (.A1(\decode.regfile.registers_13[23] ),
    .A2(_09518_),
    .B1(_09522_),
    .C1(_09512_),
    .X(_02694_));
 sky130_fd_sc_hd__nand2_2 _26371_ (.A(_09428_),
    .B(_09515_),
    .Y(_09523_));
 sky130_fd_sc_hd__o211a_2 _26372_ (.A1(\decode.regfile.registers_13[24] ),
    .A2(_09518_),
    .B1(_09523_),
    .C1(_09512_),
    .X(_02695_));
 sky130_fd_sc_hd__nand2_2 _26373_ (.A(_09430_),
    .B(_09515_),
    .Y(_09524_));
 sky130_fd_sc_hd__buf_1 _26374_ (.A(_09417_),
    .X(_09525_));
 sky130_fd_sc_hd__o211a_2 _26375_ (.A1(\decode.regfile.registers_13[25] ),
    .A2(_09518_),
    .B1(_09524_),
    .C1(_09525_),
    .X(_02696_));
 sky130_fd_sc_hd__nand2_2 _26376_ (.A(_09432_),
    .B(_09515_),
    .Y(_09526_));
 sky130_fd_sc_hd__o211a_2 _26377_ (.A1(\decode.regfile.registers_13[26] ),
    .A2(_09518_),
    .B1(_09526_),
    .C1(_09525_),
    .X(_02697_));
 sky130_fd_sc_hd__nand2_2 _26378_ (.A(_09434_),
    .B(_09515_),
    .Y(_09527_));
 sky130_fd_sc_hd__o211a_2 _26379_ (.A1(\decode.regfile.registers_13[27] ),
    .A2(_09518_),
    .B1(_09527_),
    .C1(_09525_),
    .X(_02698_));
 sky130_fd_sc_hd__nand2_2 _26380_ (.A(_09436_),
    .B(_09490_),
    .Y(_09528_));
 sky130_fd_sc_hd__o211a_2 _26381_ (.A1(\decode.regfile.registers_13[28] ),
    .A2(_09518_),
    .B1(_09528_),
    .C1(_09525_),
    .X(_02699_));
 sky130_fd_sc_hd__nand2_2 _26382_ (.A(_09438_),
    .B(_09490_),
    .Y(_09529_));
 sky130_fd_sc_hd__o211a_2 _26383_ (.A1(\decode.regfile.registers_13[29] ),
    .A2(_09518_),
    .B1(_09529_),
    .C1(_09525_),
    .X(_02700_));
 sky130_fd_sc_hd__nand2_2 _26384_ (.A(_09441_),
    .B(_09490_),
    .Y(_09530_));
 sky130_fd_sc_hd__o211a_2 _26385_ (.A1(\decode.regfile.registers_13[30] ),
    .A2(_09492_),
    .B1(_09530_),
    .C1(_09525_),
    .X(_02701_));
 sky130_fd_sc_hd__nand2_2 _26386_ (.A(_09443_),
    .B(_09490_),
    .Y(_09531_));
 sky130_fd_sc_hd__o211a_2 _26387_ (.A1(\decode.regfile.registers_13[31] ),
    .A2(_09492_),
    .B1(_09531_),
    .C1(_09525_),
    .X(_02702_));
 sky130_fd_sc_hd__and4_2 _26388_ (.A(_10373_),
    .B(_10195_),
    .C(_09932_),
    .D(_08903_),
    .X(_09532_));
 sky130_fd_sc_hd__buf_1 _26389_ (.A(_09532_),
    .X(_09533_));
 sky130_fd_sc_hd__buf_1 _26390_ (.A(_09533_),
    .X(_09534_));
 sky130_fd_sc_hd__buf_1 _26391_ (.A(_09533_),
    .X(_09535_));
 sky130_fd_sc_hd__nand2_2 _26392_ (.A(_10245_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__o211a_2 _26393_ (.A1(\decode.regfile.registers_14[0] ),
    .A2(_09534_),
    .B1(_09536_),
    .C1(_09525_),
    .X(_02703_));
 sky130_fd_sc_hd__nand2_2 _26394_ (.A(_09450_),
    .B(_09535_),
    .Y(_09537_));
 sky130_fd_sc_hd__o211a_2 _26395_ (.A1(\decode.regfile.registers_14[1] ),
    .A2(_09534_),
    .B1(_09537_),
    .C1(_09525_),
    .X(_02704_));
 sky130_fd_sc_hd__nand2_2 _26396_ (.A(_09377_),
    .B(_09535_),
    .Y(_09538_));
 sky130_fd_sc_hd__o211a_2 _26397_ (.A1(\decode.regfile.registers_14[2] ),
    .A2(_09534_),
    .B1(_09538_),
    .C1(_09525_),
    .X(_02705_));
 sky130_fd_sc_hd__nand2_2 _26398_ (.A(_09379_),
    .B(_09535_),
    .Y(_09539_));
 sky130_fd_sc_hd__buf_1 _26399_ (.A(_09417_),
    .X(_09540_));
 sky130_fd_sc_hd__o211a_2 _26400_ (.A1(\decode.regfile.registers_14[3] ),
    .A2(_09534_),
    .B1(_09539_),
    .C1(_09540_),
    .X(_02706_));
 sky130_fd_sc_hd__nand2_2 _26401_ (.A(_09381_),
    .B(_09535_),
    .Y(_09541_));
 sky130_fd_sc_hd__o211a_2 _26402_ (.A1(\decode.regfile.registers_14[4] ),
    .A2(_09534_),
    .B1(_09541_),
    .C1(_09540_),
    .X(_02707_));
 sky130_fd_sc_hd__nand2_2 _26403_ (.A(_09383_),
    .B(_09535_),
    .Y(_09542_));
 sky130_fd_sc_hd__o211a_2 _26404_ (.A1(\decode.regfile.registers_14[5] ),
    .A2(_09534_),
    .B1(_09542_),
    .C1(_09540_),
    .X(_02708_));
 sky130_fd_sc_hd__nand2_2 _26405_ (.A(_09385_),
    .B(_09535_),
    .Y(_09543_));
 sky130_fd_sc_hd__o211a_2 _26406_ (.A1(\decode.regfile.registers_14[6] ),
    .A2(_09534_),
    .B1(_09543_),
    .C1(_09540_),
    .X(_02709_));
 sky130_fd_sc_hd__nand2_2 _26407_ (.A(_09387_),
    .B(_09535_),
    .Y(_09544_));
 sky130_fd_sc_hd__o211a_2 _26408_ (.A1(\decode.regfile.registers_14[7] ),
    .A2(_09534_),
    .B1(_09544_),
    .C1(_09540_),
    .X(_02710_));
 sky130_fd_sc_hd__buf_1 _26409_ (.A(_09533_),
    .X(_09545_));
 sky130_fd_sc_hd__nand2_2 _26410_ (.A(_09389_),
    .B(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__o211a_2 _26411_ (.A1(\decode.regfile.registers_14[8] ),
    .A2(_09534_),
    .B1(_09546_),
    .C1(_09540_),
    .X(_02711_));
 sky130_fd_sc_hd__nand2_2 _26412_ (.A(_09392_),
    .B(_09545_),
    .Y(_09547_));
 sky130_fd_sc_hd__o211a_2 _26413_ (.A1(\decode.regfile.registers_14[9] ),
    .A2(_09534_),
    .B1(_09547_),
    .C1(_09540_),
    .X(_02712_));
 sky130_fd_sc_hd__buf_1 _26414_ (.A(_09533_),
    .X(_09548_));
 sky130_fd_sc_hd__nand2_2 _26415_ (.A(_09396_),
    .B(_09545_),
    .Y(_09549_));
 sky130_fd_sc_hd__o211a_2 _26416_ (.A1(\decode.regfile.registers_14[10] ),
    .A2(_09548_),
    .B1(_09549_),
    .C1(_09540_),
    .X(_02713_));
 sky130_fd_sc_hd__nand2_2 _26417_ (.A(_09398_),
    .B(_09545_),
    .Y(_09550_));
 sky130_fd_sc_hd__o211a_2 _26418_ (.A1(\decode.regfile.registers_14[11] ),
    .A2(_09548_),
    .B1(_09550_),
    .C1(_09540_),
    .X(_02714_));
 sky130_fd_sc_hd__nand2_2 _26419_ (.A(_09400_),
    .B(_09545_),
    .Y(_09551_));
 sky130_fd_sc_hd__o211a_2 _26420_ (.A1(\decode.regfile.registers_14[12] ),
    .A2(_09548_),
    .B1(_09551_),
    .C1(_09540_),
    .X(_02715_));
 sky130_fd_sc_hd__nand2_2 _26421_ (.A(_09402_),
    .B(_09545_),
    .Y(_09552_));
 sky130_fd_sc_hd__buf_1 _26422_ (.A(_09417_),
    .X(_09553_));
 sky130_fd_sc_hd__o211a_2 _26423_ (.A1(\decode.regfile.registers_14[13] ),
    .A2(_09548_),
    .B1(_09552_),
    .C1(_09553_),
    .X(_02716_));
 sky130_fd_sc_hd__nand2_2 _26424_ (.A(_09404_),
    .B(_09545_),
    .Y(_09554_));
 sky130_fd_sc_hd__o211a_2 _26425_ (.A1(\decode.regfile.registers_14[14] ),
    .A2(_09548_),
    .B1(_09554_),
    .C1(_09553_),
    .X(_02717_));
 sky130_fd_sc_hd__nand2_2 _26426_ (.A(_09406_),
    .B(_09545_),
    .Y(_09555_));
 sky130_fd_sc_hd__o211a_2 _26427_ (.A1(\decode.regfile.registers_14[15] ),
    .A2(_09548_),
    .B1(_09555_),
    .C1(_09553_),
    .X(_02718_));
 sky130_fd_sc_hd__nand2_2 _26428_ (.A(_09408_),
    .B(_09545_),
    .Y(_09556_));
 sky130_fd_sc_hd__o211a_2 _26429_ (.A1(\decode.regfile.registers_14[16] ),
    .A2(_09548_),
    .B1(_09556_),
    .C1(_09553_),
    .X(_02719_));
 sky130_fd_sc_hd__nand2_2 _26430_ (.A(_09410_),
    .B(_09545_),
    .Y(_09557_));
 sky130_fd_sc_hd__o211a_2 _26431_ (.A1(\decode.regfile.registers_14[17] ),
    .A2(_09548_),
    .B1(_09557_),
    .C1(_09553_),
    .X(_02720_));
 sky130_fd_sc_hd__buf_1 _26432_ (.A(_09533_),
    .X(_09558_));
 sky130_fd_sc_hd__nand2_2 _26433_ (.A(_09412_),
    .B(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__o211a_2 _26434_ (.A1(\decode.regfile.registers_14[18] ),
    .A2(_09548_),
    .B1(_09559_),
    .C1(_09553_),
    .X(_02721_));
 sky130_fd_sc_hd__nand2_2 _26435_ (.A(_09415_),
    .B(_09558_),
    .Y(_09560_));
 sky130_fd_sc_hd__o211a_2 _26436_ (.A1(\decode.regfile.registers_14[19] ),
    .A2(_09548_),
    .B1(_09560_),
    .C1(_09553_),
    .X(_02722_));
 sky130_fd_sc_hd__buf_1 _26437_ (.A(_09533_),
    .X(_09561_));
 sky130_fd_sc_hd__nand2_2 _26438_ (.A(_09420_),
    .B(_09558_),
    .Y(_09562_));
 sky130_fd_sc_hd__o211a_2 _26439_ (.A1(\decode.regfile.registers_14[20] ),
    .A2(_09561_),
    .B1(_09562_),
    .C1(_09553_),
    .X(_02723_));
 sky130_fd_sc_hd__nand2_2 _26440_ (.A(_09422_),
    .B(_09558_),
    .Y(_09563_));
 sky130_fd_sc_hd__o211a_2 _26441_ (.A1(\decode.regfile.registers_14[21] ),
    .A2(_09561_),
    .B1(_09563_),
    .C1(_09553_),
    .X(_02724_));
 sky130_fd_sc_hd__nand2_2 _26442_ (.A(_09424_),
    .B(_09558_),
    .Y(_09564_));
 sky130_fd_sc_hd__o211a_2 _26443_ (.A1(\decode.regfile.registers_14[22] ),
    .A2(_09561_),
    .B1(_09564_),
    .C1(_09553_),
    .X(_02725_));
 sky130_fd_sc_hd__nand2_2 _26444_ (.A(_09426_),
    .B(_09558_),
    .Y(_09565_));
 sky130_fd_sc_hd__buf_1 _26445_ (.A(_10130_),
    .X(_09566_));
 sky130_fd_sc_hd__buf_1 _26446_ (.A(_09566_),
    .X(_09567_));
 sky130_fd_sc_hd__o211a_2 _26447_ (.A1(\decode.regfile.registers_14[23] ),
    .A2(_09561_),
    .B1(_09565_),
    .C1(_09567_),
    .X(_02726_));
 sky130_fd_sc_hd__nand2_2 _26448_ (.A(_09428_),
    .B(_09558_),
    .Y(_09568_));
 sky130_fd_sc_hd__o211a_2 _26449_ (.A1(\decode.regfile.registers_14[24] ),
    .A2(_09561_),
    .B1(_09568_),
    .C1(_09567_),
    .X(_02727_));
 sky130_fd_sc_hd__nand2_2 _26450_ (.A(_09430_),
    .B(_09558_),
    .Y(_09569_));
 sky130_fd_sc_hd__o211a_2 _26451_ (.A1(\decode.regfile.registers_14[25] ),
    .A2(_09561_),
    .B1(_09569_),
    .C1(_09567_),
    .X(_02728_));
 sky130_fd_sc_hd__nand2_2 _26452_ (.A(_09432_),
    .B(_09558_),
    .Y(_09570_));
 sky130_fd_sc_hd__o211a_2 _26453_ (.A1(\decode.regfile.registers_14[26] ),
    .A2(_09561_),
    .B1(_09570_),
    .C1(_09567_),
    .X(_02729_));
 sky130_fd_sc_hd__nand2_2 _26454_ (.A(_09434_),
    .B(_09558_),
    .Y(_09571_));
 sky130_fd_sc_hd__o211a_2 _26455_ (.A1(\decode.regfile.registers_14[27] ),
    .A2(_09561_),
    .B1(_09571_),
    .C1(_09567_),
    .X(_02730_));
 sky130_fd_sc_hd__nand2_2 _26456_ (.A(_09436_),
    .B(_09533_),
    .Y(_09572_));
 sky130_fd_sc_hd__o211a_2 _26457_ (.A1(\decode.regfile.registers_14[28] ),
    .A2(_09561_),
    .B1(_09572_),
    .C1(_09567_),
    .X(_02731_));
 sky130_fd_sc_hd__nand2_2 _26458_ (.A(_09438_),
    .B(_09533_),
    .Y(_09573_));
 sky130_fd_sc_hd__o211a_2 _26459_ (.A1(\decode.regfile.registers_14[29] ),
    .A2(_09561_),
    .B1(_09573_),
    .C1(_09567_),
    .X(_02732_));
 sky130_fd_sc_hd__nand2_2 _26460_ (.A(_09441_),
    .B(_09533_),
    .Y(_09574_));
 sky130_fd_sc_hd__o211a_2 _26461_ (.A1(\decode.regfile.registers_14[30] ),
    .A2(_09535_),
    .B1(_09574_),
    .C1(_09567_),
    .X(_02733_));
 sky130_fd_sc_hd__nand2_2 _26462_ (.A(_09443_),
    .B(_09533_),
    .Y(_09575_));
 sky130_fd_sc_hd__o211a_2 _26463_ (.A1(\decode.regfile.registers_14[31] ),
    .A2(_09535_),
    .B1(_09575_),
    .C1(_09567_),
    .X(_02734_));
 sky130_fd_sc_hd__and4_2 _26464_ (.A(_09929_),
    .B(_10195_),
    .C(_10150_),
    .D(_08903_),
    .X(_09576_));
 sky130_fd_sc_hd__buf_1 _26465_ (.A(_09576_),
    .X(_09577_));
 sky130_fd_sc_hd__buf_1 _26466_ (.A(_09577_),
    .X(_09578_));
 sky130_fd_sc_hd__buf_1 _26467_ (.A(_09577_),
    .X(_09579_));
 sky130_fd_sc_hd__nand2_2 _26468_ (.A(_10245_),
    .B(_09579_),
    .Y(_09580_));
 sky130_fd_sc_hd__o211a_2 _26469_ (.A1(\decode.regfile.registers_15[0] ),
    .A2(_09578_),
    .B1(_09580_),
    .C1(_09567_),
    .X(_02735_));
 sky130_fd_sc_hd__nand2_2 _26470_ (.A(_09450_),
    .B(_09579_),
    .Y(_09581_));
 sky130_fd_sc_hd__buf_1 _26471_ (.A(_09566_),
    .X(_09582_));
 sky130_fd_sc_hd__o211a_2 _26472_ (.A1(\decode.regfile.registers_15[1] ),
    .A2(_09578_),
    .B1(_09581_),
    .C1(_09582_),
    .X(_02736_));
 sky130_fd_sc_hd__nand2_2 _26473_ (.A(_09377_),
    .B(_09579_),
    .Y(_09583_));
 sky130_fd_sc_hd__o211a_2 _26474_ (.A1(\decode.regfile.registers_15[2] ),
    .A2(_09578_),
    .B1(_09583_),
    .C1(_09582_),
    .X(_02737_));
 sky130_fd_sc_hd__nand2_2 _26475_ (.A(_09379_),
    .B(_09579_),
    .Y(_09584_));
 sky130_fd_sc_hd__o211a_2 _26476_ (.A1(\decode.regfile.registers_15[3] ),
    .A2(_09578_),
    .B1(_09584_),
    .C1(_09582_),
    .X(_02738_));
 sky130_fd_sc_hd__nand2_2 _26477_ (.A(_09381_),
    .B(_09579_),
    .Y(_09585_));
 sky130_fd_sc_hd__o211a_2 _26478_ (.A1(\decode.regfile.registers_15[4] ),
    .A2(_09578_),
    .B1(_09585_),
    .C1(_09582_),
    .X(_02739_));
 sky130_fd_sc_hd__nand2_2 _26479_ (.A(_09383_),
    .B(_09579_),
    .Y(_09586_));
 sky130_fd_sc_hd__o211a_2 _26480_ (.A1(\decode.regfile.registers_15[5] ),
    .A2(_09578_),
    .B1(_09586_),
    .C1(_09582_),
    .X(_02740_));
 sky130_fd_sc_hd__nand2_2 _26481_ (.A(_09385_),
    .B(_09579_),
    .Y(_09587_));
 sky130_fd_sc_hd__o211a_2 _26482_ (.A1(\decode.regfile.registers_15[6] ),
    .A2(_09578_),
    .B1(_09587_),
    .C1(_09582_),
    .X(_02741_));
 sky130_fd_sc_hd__nand2_2 _26483_ (.A(_09387_),
    .B(_09579_),
    .Y(_09588_));
 sky130_fd_sc_hd__o211a_2 _26484_ (.A1(\decode.regfile.registers_15[7] ),
    .A2(_09578_),
    .B1(_09588_),
    .C1(_09582_),
    .X(_02742_));
 sky130_fd_sc_hd__buf_1 _26485_ (.A(_09577_),
    .X(_09589_));
 sky130_fd_sc_hd__nand2_2 _26486_ (.A(_09389_),
    .B(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__o211a_2 _26487_ (.A1(\decode.regfile.registers_15[8] ),
    .A2(_09578_),
    .B1(_09590_),
    .C1(_09582_),
    .X(_02743_));
 sky130_fd_sc_hd__nand2_2 _26488_ (.A(_09392_),
    .B(_09589_),
    .Y(_09591_));
 sky130_fd_sc_hd__o211a_2 _26489_ (.A1(\decode.regfile.registers_15[9] ),
    .A2(_09578_),
    .B1(_09591_),
    .C1(_09582_),
    .X(_02744_));
 sky130_fd_sc_hd__buf_1 _26490_ (.A(_09577_),
    .X(_09592_));
 sky130_fd_sc_hd__nand2_2 _26491_ (.A(_09396_),
    .B(_09589_),
    .Y(_09593_));
 sky130_fd_sc_hd__o211a_2 _26492_ (.A1(\decode.regfile.registers_15[10] ),
    .A2(_09592_),
    .B1(_09593_),
    .C1(_09582_),
    .X(_02745_));
 sky130_fd_sc_hd__nand2_2 _26493_ (.A(_09398_),
    .B(_09589_),
    .Y(_09594_));
 sky130_fd_sc_hd__buf_1 _26494_ (.A(_09566_),
    .X(_09595_));
 sky130_fd_sc_hd__o211a_2 _26495_ (.A1(\decode.regfile.registers_15[11] ),
    .A2(_09592_),
    .B1(_09594_),
    .C1(_09595_),
    .X(_02746_));
 sky130_fd_sc_hd__nand2_2 _26496_ (.A(_09400_),
    .B(_09589_),
    .Y(_09596_));
 sky130_fd_sc_hd__o211a_2 _26497_ (.A1(\decode.regfile.registers_15[12] ),
    .A2(_09592_),
    .B1(_09596_),
    .C1(_09595_),
    .X(_02747_));
 sky130_fd_sc_hd__nand2_2 _26498_ (.A(_09402_),
    .B(_09589_),
    .Y(_09597_));
 sky130_fd_sc_hd__o211a_2 _26499_ (.A1(\decode.regfile.registers_15[13] ),
    .A2(_09592_),
    .B1(_09597_),
    .C1(_09595_),
    .X(_02748_));
 sky130_fd_sc_hd__nand2_2 _26500_ (.A(_09404_),
    .B(_09589_),
    .Y(_09598_));
 sky130_fd_sc_hd__o211a_2 _26501_ (.A1(\decode.regfile.registers_15[14] ),
    .A2(_09592_),
    .B1(_09598_),
    .C1(_09595_),
    .X(_02749_));
 sky130_fd_sc_hd__nand2_2 _26502_ (.A(_09406_),
    .B(_09589_),
    .Y(_09599_));
 sky130_fd_sc_hd__o211a_2 _26503_ (.A1(\decode.regfile.registers_15[15] ),
    .A2(_09592_),
    .B1(_09599_),
    .C1(_09595_),
    .X(_02750_));
 sky130_fd_sc_hd__nand2_2 _26504_ (.A(_09408_),
    .B(_09589_),
    .Y(_09600_));
 sky130_fd_sc_hd__o211a_2 _26505_ (.A1(\decode.regfile.registers_15[16] ),
    .A2(_09592_),
    .B1(_09600_),
    .C1(_09595_),
    .X(_02751_));
 sky130_fd_sc_hd__nand2_2 _26506_ (.A(_09410_),
    .B(_09589_),
    .Y(_09601_));
 sky130_fd_sc_hd__o211a_2 _26507_ (.A1(\decode.regfile.registers_15[17] ),
    .A2(_09592_),
    .B1(_09601_),
    .C1(_09595_),
    .X(_02752_));
 sky130_fd_sc_hd__buf_1 _26508_ (.A(_09577_),
    .X(_09602_));
 sky130_fd_sc_hd__nand2_2 _26509_ (.A(_09412_),
    .B(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__o211a_2 _26510_ (.A1(\decode.regfile.registers_15[18] ),
    .A2(_09592_),
    .B1(_09603_),
    .C1(_09595_),
    .X(_02753_));
 sky130_fd_sc_hd__nand2_2 _26511_ (.A(_09415_),
    .B(_09602_),
    .Y(_09604_));
 sky130_fd_sc_hd__o211a_2 _26512_ (.A1(\decode.regfile.registers_15[19] ),
    .A2(_09592_),
    .B1(_09604_),
    .C1(_09595_),
    .X(_02754_));
 sky130_fd_sc_hd__buf_1 _26513_ (.A(_09577_),
    .X(_09605_));
 sky130_fd_sc_hd__nand2_2 _26514_ (.A(_09420_),
    .B(_09602_),
    .Y(_09606_));
 sky130_fd_sc_hd__o211a_2 _26515_ (.A1(\decode.regfile.registers_15[20] ),
    .A2(_09605_),
    .B1(_09606_),
    .C1(_09595_),
    .X(_02755_));
 sky130_fd_sc_hd__nand2_2 _26516_ (.A(_09422_),
    .B(_09602_),
    .Y(_09607_));
 sky130_fd_sc_hd__buf_1 _26517_ (.A(_09566_),
    .X(_09608_));
 sky130_fd_sc_hd__o211a_2 _26518_ (.A1(\decode.regfile.registers_15[21] ),
    .A2(_09605_),
    .B1(_09607_),
    .C1(_09608_),
    .X(_02756_));
 sky130_fd_sc_hd__nand2_2 _26519_ (.A(_09424_),
    .B(_09602_),
    .Y(_09609_));
 sky130_fd_sc_hd__o211a_2 _26520_ (.A1(\decode.regfile.registers_15[22] ),
    .A2(_09605_),
    .B1(_09609_),
    .C1(_09608_),
    .X(_02757_));
 sky130_fd_sc_hd__nand2_2 _26521_ (.A(_09426_),
    .B(_09602_),
    .Y(_09610_));
 sky130_fd_sc_hd__o211a_2 _26522_ (.A1(\decode.regfile.registers_15[23] ),
    .A2(_09605_),
    .B1(_09610_),
    .C1(_09608_),
    .X(_02758_));
 sky130_fd_sc_hd__nand2_2 _26523_ (.A(_09428_),
    .B(_09602_),
    .Y(_09611_));
 sky130_fd_sc_hd__o211a_2 _26524_ (.A1(\decode.regfile.registers_15[24] ),
    .A2(_09605_),
    .B1(_09611_),
    .C1(_09608_),
    .X(_02759_));
 sky130_fd_sc_hd__nand2_2 _26525_ (.A(_09430_),
    .B(_09602_),
    .Y(_09612_));
 sky130_fd_sc_hd__o211a_2 _26526_ (.A1(\decode.regfile.registers_15[25] ),
    .A2(_09605_),
    .B1(_09612_),
    .C1(_09608_),
    .X(_02760_));
 sky130_fd_sc_hd__nand2_2 _26527_ (.A(_09432_),
    .B(_09602_),
    .Y(_09613_));
 sky130_fd_sc_hd__o211a_2 _26528_ (.A1(\decode.regfile.registers_15[26] ),
    .A2(_09605_),
    .B1(_09613_),
    .C1(_09608_),
    .X(_02761_));
 sky130_fd_sc_hd__nand2_2 _26529_ (.A(_09434_),
    .B(_09602_),
    .Y(_09614_));
 sky130_fd_sc_hd__o211a_2 _26530_ (.A1(\decode.regfile.registers_15[27] ),
    .A2(_09605_),
    .B1(_09614_),
    .C1(_09608_),
    .X(_02762_));
 sky130_fd_sc_hd__nand2_2 _26531_ (.A(_09436_),
    .B(_09577_),
    .Y(_09615_));
 sky130_fd_sc_hd__o211a_2 _26532_ (.A1(\decode.regfile.registers_15[28] ),
    .A2(_09605_),
    .B1(_09615_),
    .C1(_09608_),
    .X(_02763_));
 sky130_fd_sc_hd__nand2_2 _26533_ (.A(_09438_),
    .B(_09577_),
    .Y(_09616_));
 sky130_fd_sc_hd__o211a_2 _26534_ (.A1(\decode.regfile.registers_15[29] ),
    .A2(_09605_),
    .B1(_09616_),
    .C1(_09608_),
    .X(_02764_));
 sky130_fd_sc_hd__nand2_2 _26535_ (.A(_09441_),
    .B(_09577_),
    .Y(_09617_));
 sky130_fd_sc_hd__o211a_2 _26536_ (.A1(\decode.regfile.registers_15[30] ),
    .A2(_09579_),
    .B1(_09617_),
    .C1(_09608_),
    .X(_02765_));
 sky130_fd_sc_hd__nand2_2 _26537_ (.A(_09443_),
    .B(_09577_),
    .Y(_09618_));
 sky130_fd_sc_hd__buf_1 _26538_ (.A(_09566_),
    .X(_09619_));
 sky130_fd_sc_hd__o211a_2 _26539_ (.A1(\decode.regfile.registers_15[31] ),
    .A2(_09579_),
    .B1(_09618_),
    .C1(_09619_),
    .X(_02766_));
 sky130_fd_sc_hd__and3_2 _26540_ (.A(_10149_),
    .B(_10196_),
    .C(_03672_),
    .X(_09620_));
 sky130_fd_sc_hd__buf_1 _26541_ (.A(_09620_),
    .X(_09621_));
 sky130_fd_sc_hd__buf_1 _26542_ (.A(_09621_),
    .X(_09622_));
 sky130_fd_sc_hd__buf_1 _26543_ (.A(_09621_),
    .X(_09623_));
 sky130_fd_sc_hd__nand2_2 _26544_ (.A(_10245_),
    .B(_09623_),
    .Y(_09624_));
 sky130_fd_sc_hd__o211a_2 _26545_ (.A1(\decode.regfile.registers_16[0] ),
    .A2(_09622_),
    .B1(_09624_),
    .C1(_09619_),
    .X(_02767_));
 sky130_fd_sc_hd__nand2_2 _26546_ (.A(_09450_),
    .B(_09623_),
    .Y(_09625_));
 sky130_fd_sc_hd__o211a_2 _26547_ (.A1(\decode.regfile.registers_16[1] ),
    .A2(_09622_),
    .B1(_09625_),
    .C1(_09619_),
    .X(_02768_));
 sky130_fd_sc_hd__nand2_2 _26548_ (.A(_09377_),
    .B(_09623_),
    .Y(_09626_));
 sky130_fd_sc_hd__o211a_2 _26549_ (.A1(\decode.regfile.registers_16[2] ),
    .A2(_09622_),
    .B1(_09626_),
    .C1(_09619_),
    .X(_02769_));
 sky130_fd_sc_hd__nand2_2 _26550_ (.A(_09379_),
    .B(_09623_),
    .Y(_09627_));
 sky130_fd_sc_hd__o211a_2 _26551_ (.A1(\decode.regfile.registers_16[3] ),
    .A2(_09622_),
    .B1(_09627_),
    .C1(_09619_),
    .X(_02770_));
 sky130_fd_sc_hd__nand2_2 _26552_ (.A(_09381_),
    .B(_09623_),
    .Y(_09628_));
 sky130_fd_sc_hd__o211a_2 _26553_ (.A1(\decode.regfile.registers_16[4] ),
    .A2(_09622_),
    .B1(_09628_),
    .C1(_09619_),
    .X(_02771_));
 sky130_fd_sc_hd__nand2_2 _26554_ (.A(_09383_),
    .B(_09623_),
    .Y(_09629_));
 sky130_fd_sc_hd__o211a_2 _26555_ (.A1(\decode.regfile.registers_16[5] ),
    .A2(_09622_),
    .B1(_09629_),
    .C1(_09619_),
    .X(_02772_));
 sky130_fd_sc_hd__nand2_2 _26556_ (.A(_09385_),
    .B(_09623_),
    .Y(_09630_));
 sky130_fd_sc_hd__o211a_2 _26557_ (.A1(\decode.regfile.registers_16[6] ),
    .A2(_09622_),
    .B1(_09630_),
    .C1(_09619_),
    .X(_02773_));
 sky130_fd_sc_hd__nand2_2 _26558_ (.A(_09387_),
    .B(_09623_),
    .Y(_09631_));
 sky130_fd_sc_hd__o211a_2 _26559_ (.A1(\decode.regfile.registers_16[7] ),
    .A2(_09622_),
    .B1(_09631_),
    .C1(_09619_),
    .X(_02774_));
 sky130_fd_sc_hd__buf_1 _26560_ (.A(_09621_),
    .X(_09632_));
 sky130_fd_sc_hd__nand2_2 _26561_ (.A(_09389_),
    .B(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__o211a_2 _26562_ (.A1(\decode.regfile.registers_16[8] ),
    .A2(_09622_),
    .B1(_09633_),
    .C1(_09619_),
    .X(_02775_));
 sky130_fd_sc_hd__nand2_2 _26563_ (.A(_09392_),
    .B(_09632_),
    .Y(_09634_));
 sky130_fd_sc_hd__buf_1 _26564_ (.A(_09566_),
    .X(_09635_));
 sky130_fd_sc_hd__o211a_2 _26565_ (.A1(\decode.regfile.registers_16[9] ),
    .A2(_09622_),
    .B1(_09634_),
    .C1(_09635_),
    .X(_02776_));
 sky130_fd_sc_hd__buf_1 _26566_ (.A(_09621_),
    .X(_09636_));
 sky130_fd_sc_hd__nand2_2 _26567_ (.A(_09396_),
    .B(_09632_),
    .Y(_09637_));
 sky130_fd_sc_hd__o211a_2 _26568_ (.A1(\decode.regfile.registers_16[10] ),
    .A2(_09636_),
    .B1(_09637_),
    .C1(_09635_),
    .X(_02777_));
 sky130_fd_sc_hd__nand2_2 _26569_ (.A(_09398_),
    .B(_09632_),
    .Y(_09638_));
 sky130_fd_sc_hd__o211a_2 _26570_ (.A1(\decode.regfile.registers_16[11] ),
    .A2(_09636_),
    .B1(_09638_),
    .C1(_09635_),
    .X(_02778_));
 sky130_fd_sc_hd__nand2_2 _26571_ (.A(_09400_),
    .B(_09632_),
    .Y(_09639_));
 sky130_fd_sc_hd__o211a_2 _26572_ (.A1(\decode.regfile.registers_16[12] ),
    .A2(_09636_),
    .B1(_09639_),
    .C1(_09635_),
    .X(_02779_));
 sky130_fd_sc_hd__nand2_2 _26573_ (.A(_09402_),
    .B(_09632_),
    .Y(_09640_));
 sky130_fd_sc_hd__o211a_2 _26574_ (.A1(\decode.regfile.registers_16[13] ),
    .A2(_09636_),
    .B1(_09640_),
    .C1(_09635_),
    .X(_02780_));
 sky130_fd_sc_hd__nand2_2 _26575_ (.A(_09404_),
    .B(_09632_),
    .Y(_09641_));
 sky130_fd_sc_hd__o211a_2 _26576_ (.A1(\decode.regfile.registers_16[14] ),
    .A2(_09636_),
    .B1(_09641_),
    .C1(_09635_),
    .X(_02781_));
 sky130_fd_sc_hd__nand2_2 _26577_ (.A(_09406_),
    .B(_09632_),
    .Y(_09642_));
 sky130_fd_sc_hd__o211a_2 _26578_ (.A1(\decode.regfile.registers_16[15] ),
    .A2(_09636_),
    .B1(_09642_),
    .C1(_09635_),
    .X(_02782_));
 sky130_fd_sc_hd__nand2_2 _26579_ (.A(_09408_),
    .B(_09632_),
    .Y(_09643_));
 sky130_fd_sc_hd__o211a_2 _26580_ (.A1(\decode.regfile.registers_16[16] ),
    .A2(_09636_),
    .B1(_09643_),
    .C1(_09635_),
    .X(_02783_));
 sky130_fd_sc_hd__nand2_2 _26581_ (.A(_09410_),
    .B(_09632_),
    .Y(_09644_));
 sky130_fd_sc_hd__o211a_2 _26582_ (.A1(\decode.regfile.registers_16[17] ),
    .A2(_09636_),
    .B1(_09644_),
    .C1(_09635_),
    .X(_02784_));
 sky130_fd_sc_hd__buf_1 _26583_ (.A(_09621_),
    .X(_09645_));
 sky130_fd_sc_hd__nand2_2 _26584_ (.A(_09412_),
    .B(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__o211a_2 _26585_ (.A1(\decode.regfile.registers_16[18] ),
    .A2(_09636_),
    .B1(_09646_),
    .C1(_09635_),
    .X(_02785_));
 sky130_fd_sc_hd__nand2_2 _26586_ (.A(_09415_),
    .B(_09645_),
    .Y(_09647_));
 sky130_fd_sc_hd__buf_1 _26587_ (.A(_09566_),
    .X(_09648_));
 sky130_fd_sc_hd__o211a_2 _26588_ (.A1(\decode.regfile.registers_16[19] ),
    .A2(_09636_),
    .B1(_09647_),
    .C1(_09648_),
    .X(_02786_));
 sky130_fd_sc_hd__buf_1 _26589_ (.A(_09621_),
    .X(_09649_));
 sky130_fd_sc_hd__nand2_2 _26590_ (.A(_09420_),
    .B(_09645_),
    .Y(_09650_));
 sky130_fd_sc_hd__o211a_2 _26591_ (.A1(\decode.regfile.registers_16[20] ),
    .A2(_09649_),
    .B1(_09650_),
    .C1(_09648_),
    .X(_02787_));
 sky130_fd_sc_hd__nand2_2 _26592_ (.A(_09422_),
    .B(_09645_),
    .Y(_09651_));
 sky130_fd_sc_hd__o211a_2 _26593_ (.A1(\decode.regfile.registers_16[21] ),
    .A2(_09649_),
    .B1(_09651_),
    .C1(_09648_),
    .X(_02788_));
 sky130_fd_sc_hd__nand2_2 _26594_ (.A(_09424_),
    .B(_09645_),
    .Y(_09652_));
 sky130_fd_sc_hd__o211a_2 _26595_ (.A1(\decode.regfile.registers_16[22] ),
    .A2(_09649_),
    .B1(_09652_),
    .C1(_09648_),
    .X(_02789_));
 sky130_fd_sc_hd__nand2_2 _26596_ (.A(_09426_),
    .B(_09645_),
    .Y(_09653_));
 sky130_fd_sc_hd__o211a_2 _26597_ (.A1(\decode.regfile.registers_16[23] ),
    .A2(_09649_),
    .B1(_09653_),
    .C1(_09648_),
    .X(_02790_));
 sky130_fd_sc_hd__nand2_2 _26598_ (.A(_09428_),
    .B(_09645_),
    .Y(_09654_));
 sky130_fd_sc_hd__o211a_2 _26599_ (.A1(\decode.regfile.registers_16[24] ),
    .A2(_09649_),
    .B1(_09654_),
    .C1(_09648_),
    .X(_02791_));
 sky130_fd_sc_hd__nand2_2 _26600_ (.A(_09430_),
    .B(_09645_),
    .Y(_09655_));
 sky130_fd_sc_hd__o211a_2 _26601_ (.A1(\decode.regfile.registers_16[25] ),
    .A2(_09649_),
    .B1(_09655_),
    .C1(_09648_),
    .X(_02792_));
 sky130_fd_sc_hd__nand2_2 _26602_ (.A(_09432_),
    .B(_09645_),
    .Y(_09656_));
 sky130_fd_sc_hd__o211a_2 _26603_ (.A1(\decode.regfile.registers_16[26] ),
    .A2(_09649_),
    .B1(_09656_),
    .C1(_09648_),
    .X(_02793_));
 sky130_fd_sc_hd__nand2_2 _26604_ (.A(_09434_),
    .B(_09645_),
    .Y(_09657_));
 sky130_fd_sc_hd__o211a_2 _26605_ (.A1(\decode.regfile.registers_16[27] ),
    .A2(_09649_),
    .B1(_09657_),
    .C1(_09648_),
    .X(_02794_));
 sky130_fd_sc_hd__nand2_2 _26606_ (.A(_09436_),
    .B(_09621_),
    .Y(_09658_));
 sky130_fd_sc_hd__o211a_2 _26607_ (.A1(\decode.regfile.registers_16[28] ),
    .A2(_09649_),
    .B1(_09658_),
    .C1(_09648_),
    .X(_02795_));
 sky130_fd_sc_hd__nand2_2 _26608_ (.A(_09438_),
    .B(_09621_),
    .Y(_09659_));
 sky130_fd_sc_hd__buf_1 _26609_ (.A(_09566_),
    .X(_09660_));
 sky130_fd_sc_hd__o211a_2 _26610_ (.A1(\decode.regfile.registers_16[29] ),
    .A2(_09649_),
    .B1(_09659_),
    .C1(_09660_),
    .X(_02796_));
 sky130_fd_sc_hd__nand2_2 _26611_ (.A(_09441_),
    .B(_09621_),
    .Y(_09661_));
 sky130_fd_sc_hd__o211a_2 _26612_ (.A1(\decode.regfile.registers_16[30] ),
    .A2(_09623_),
    .B1(_09661_),
    .C1(_09660_),
    .X(_02797_));
 sky130_fd_sc_hd__nand2_2 _26613_ (.A(_09443_),
    .B(_09621_),
    .Y(_09662_));
 sky130_fd_sc_hd__o211a_2 _26614_ (.A1(\decode.regfile.registers_16[31] ),
    .A2(_09623_),
    .B1(_09662_),
    .C1(_09660_),
    .X(_02798_));
 sky130_fd_sc_hd__and3_2 _26615_ (.A(_10149_),
    .B(_10240_),
    .C(_03672_),
    .X(_09663_));
 sky130_fd_sc_hd__buf_1 _26616_ (.A(_09663_),
    .X(_09664_));
 sky130_fd_sc_hd__buf_1 _26617_ (.A(_09664_),
    .X(_09665_));
 sky130_fd_sc_hd__buf_1 _26618_ (.A(_09664_),
    .X(_09666_));
 sky130_fd_sc_hd__nand2_2 _26619_ (.A(_10245_),
    .B(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__o211a_2 _26620_ (.A1(\decode.regfile.registers_17[0] ),
    .A2(_09665_),
    .B1(_09667_),
    .C1(_09660_),
    .X(_02799_));
 sky130_fd_sc_hd__nand2_2 _26621_ (.A(_09450_),
    .B(_09666_),
    .Y(_09668_));
 sky130_fd_sc_hd__o211a_2 _26622_ (.A1(\decode.regfile.registers_17[1] ),
    .A2(_09665_),
    .B1(_09668_),
    .C1(_09660_),
    .X(_02800_));
 sky130_fd_sc_hd__nand2_2 _26623_ (.A(_09377_),
    .B(_09666_),
    .Y(_09669_));
 sky130_fd_sc_hd__o211a_2 _26624_ (.A1(\decode.regfile.registers_17[2] ),
    .A2(_09665_),
    .B1(_09669_),
    .C1(_09660_),
    .X(_02801_));
 sky130_fd_sc_hd__nand2_2 _26625_ (.A(_09379_),
    .B(_09666_),
    .Y(_09670_));
 sky130_fd_sc_hd__o211a_2 _26626_ (.A1(\decode.regfile.registers_17[3] ),
    .A2(_09665_),
    .B1(_09670_),
    .C1(_09660_),
    .X(_02802_));
 sky130_fd_sc_hd__nand2_2 _26627_ (.A(_09381_),
    .B(_09666_),
    .Y(_09671_));
 sky130_fd_sc_hd__o211a_2 _26628_ (.A1(\decode.regfile.registers_17[4] ),
    .A2(_09665_),
    .B1(_09671_),
    .C1(_09660_),
    .X(_02803_));
 sky130_fd_sc_hd__nand2_2 _26629_ (.A(_09383_),
    .B(_09666_),
    .Y(_09672_));
 sky130_fd_sc_hd__o211a_2 _26630_ (.A1(\decode.regfile.registers_17[5] ),
    .A2(_09665_),
    .B1(_09672_),
    .C1(_09660_),
    .X(_02804_));
 sky130_fd_sc_hd__nand2_2 _26631_ (.A(_09385_),
    .B(_09666_),
    .Y(_09673_));
 sky130_fd_sc_hd__o211a_2 _26632_ (.A1(\decode.regfile.registers_17[6] ),
    .A2(_09665_),
    .B1(_09673_),
    .C1(_09660_),
    .X(_02805_));
 sky130_fd_sc_hd__nand2_2 _26633_ (.A(_09387_),
    .B(_09666_),
    .Y(_09674_));
 sky130_fd_sc_hd__buf_1 _26634_ (.A(_09566_),
    .X(_09675_));
 sky130_fd_sc_hd__o211a_2 _26635_ (.A1(\decode.regfile.registers_17[7] ),
    .A2(_09665_),
    .B1(_09674_),
    .C1(_09675_),
    .X(_02806_));
 sky130_fd_sc_hd__buf_1 _26636_ (.A(_09664_),
    .X(_09676_));
 sky130_fd_sc_hd__nand2_2 _26637_ (.A(_09389_),
    .B(_09676_),
    .Y(_09677_));
 sky130_fd_sc_hd__o211a_2 _26638_ (.A1(\decode.regfile.registers_17[8] ),
    .A2(_09665_),
    .B1(_09677_),
    .C1(_09675_),
    .X(_02807_));
 sky130_fd_sc_hd__nand2_2 _26639_ (.A(_09392_),
    .B(_09676_),
    .Y(_09678_));
 sky130_fd_sc_hd__o211a_2 _26640_ (.A1(\decode.regfile.registers_17[9] ),
    .A2(_09665_),
    .B1(_09678_),
    .C1(_09675_),
    .X(_02808_));
 sky130_fd_sc_hd__buf_1 _26641_ (.A(_09664_),
    .X(_09679_));
 sky130_fd_sc_hd__nand2_2 _26642_ (.A(_09396_),
    .B(_09676_),
    .Y(_09680_));
 sky130_fd_sc_hd__o211a_2 _26643_ (.A1(\decode.regfile.registers_17[10] ),
    .A2(_09679_),
    .B1(_09680_),
    .C1(_09675_),
    .X(_02809_));
 sky130_fd_sc_hd__nand2_2 _26644_ (.A(_09398_),
    .B(_09676_),
    .Y(_09681_));
 sky130_fd_sc_hd__o211a_2 _26645_ (.A1(\decode.regfile.registers_17[11] ),
    .A2(_09679_),
    .B1(_09681_),
    .C1(_09675_),
    .X(_02810_));
 sky130_fd_sc_hd__nand2_2 _26646_ (.A(_09400_),
    .B(_09676_),
    .Y(_09682_));
 sky130_fd_sc_hd__o211a_2 _26647_ (.A1(\decode.regfile.registers_17[12] ),
    .A2(_09679_),
    .B1(_09682_),
    .C1(_09675_),
    .X(_02811_));
 sky130_fd_sc_hd__nand2_2 _26648_ (.A(_09402_),
    .B(_09676_),
    .Y(_09683_));
 sky130_fd_sc_hd__o211a_2 _26649_ (.A1(\decode.regfile.registers_17[13] ),
    .A2(_09679_),
    .B1(_09683_),
    .C1(_09675_),
    .X(_02812_));
 sky130_fd_sc_hd__nand2_2 _26650_ (.A(_09404_),
    .B(_09676_),
    .Y(_09684_));
 sky130_fd_sc_hd__o211a_2 _26651_ (.A1(\decode.regfile.registers_17[14] ),
    .A2(_09679_),
    .B1(_09684_),
    .C1(_09675_),
    .X(_02813_));
 sky130_fd_sc_hd__nand2_2 _26652_ (.A(_09406_),
    .B(_09676_),
    .Y(_09685_));
 sky130_fd_sc_hd__o211a_2 _26653_ (.A1(\decode.regfile.registers_17[15] ),
    .A2(_09679_),
    .B1(_09685_),
    .C1(_09675_),
    .X(_02814_));
 sky130_fd_sc_hd__nand2_2 _26654_ (.A(_09408_),
    .B(_09676_),
    .Y(_09686_));
 sky130_fd_sc_hd__o211a_2 _26655_ (.A1(\decode.regfile.registers_17[16] ),
    .A2(_09679_),
    .B1(_09686_),
    .C1(_09675_),
    .X(_02815_));
 sky130_fd_sc_hd__nand2_2 _26656_ (.A(_09410_),
    .B(_09676_),
    .Y(_09687_));
 sky130_fd_sc_hd__buf_1 _26657_ (.A(_09566_),
    .X(_09688_));
 sky130_fd_sc_hd__o211a_2 _26658_ (.A1(\decode.regfile.registers_17[17] ),
    .A2(_09679_),
    .B1(_09687_),
    .C1(_09688_),
    .X(_02816_));
 sky130_fd_sc_hd__buf_1 _26659_ (.A(_09664_),
    .X(_09689_));
 sky130_fd_sc_hd__nand2_2 _26660_ (.A(_09412_),
    .B(_09689_),
    .Y(_09690_));
 sky130_fd_sc_hd__o211a_2 _26661_ (.A1(\decode.regfile.registers_17[18] ),
    .A2(_09679_),
    .B1(_09690_),
    .C1(_09688_),
    .X(_02817_));
 sky130_fd_sc_hd__nand2_2 _26662_ (.A(_09415_),
    .B(_09689_),
    .Y(_09691_));
 sky130_fd_sc_hd__o211a_2 _26663_ (.A1(\decode.regfile.registers_17[19] ),
    .A2(_09679_),
    .B1(_09691_),
    .C1(_09688_),
    .X(_02818_));
 sky130_fd_sc_hd__buf_1 _26664_ (.A(_09664_),
    .X(_09692_));
 sky130_fd_sc_hd__nand2_2 _26665_ (.A(_09420_),
    .B(_09689_),
    .Y(_09693_));
 sky130_fd_sc_hd__o211a_2 _26666_ (.A1(\decode.regfile.registers_17[20] ),
    .A2(_09692_),
    .B1(_09693_),
    .C1(_09688_),
    .X(_02819_));
 sky130_fd_sc_hd__nand2_2 _26667_ (.A(_09422_),
    .B(_09689_),
    .Y(_09694_));
 sky130_fd_sc_hd__o211a_2 _26668_ (.A1(\decode.regfile.registers_17[21] ),
    .A2(_09692_),
    .B1(_09694_),
    .C1(_09688_),
    .X(_02820_));
 sky130_fd_sc_hd__nand2_2 _26669_ (.A(_09424_),
    .B(_09689_),
    .Y(_09695_));
 sky130_fd_sc_hd__o211a_2 _26670_ (.A1(\decode.regfile.registers_17[22] ),
    .A2(_09692_),
    .B1(_09695_),
    .C1(_09688_),
    .X(_02821_));
 sky130_fd_sc_hd__nand2_2 _26671_ (.A(_09426_),
    .B(_09689_),
    .Y(_09696_));
 sky130_fd_sc_hd__o211a_2 _26672_ (.A1(\decode.regfile.registers_17[23] ),
    .A2(_09692_),
    .B1(_09696_),
    .C1(_09688_),
    .X(_02822_));
 sky130_fd_sc_hd__nand2_2 _26673_ (.A(_09428_),
    .B(_09689_),
    .Y(_09697_));
 sky130_fd_sc_hd__o211a_2 _26674_ (.A1(\decode.regfile.registers_17[24] ),
    .A2(_09692_),
    .B1(_09697_),
    .C1(_09688_),
    .X(_02823_));
 sky130_fd_sc_hd__nand2_2 _26675_ (.A(_09430_),
    .B(_09689_),
    .Y(_09698_));
 sky130_fd_sc_hd__o211a_2 _26676_ (.A1(\decode.regfile.registers_17[25] ),
    .A2(_09692_),
    .B1(_09698_),
    .C1(_09688_),
    .X(_02824_));
 sky130_fd_sc_hd__nand2_2 _26677_ (.A(_09432_),
    .B(_09689_),
    .Y(_09699_));
 sky130_fd_sc_hd__o211a_2 _26678_ (.A1(\decode.regfile.registers_17[26] ),
    .A2(_09692_),
    .B1(_09699_),
    .C1(_09688_),
    .X(_02825_));
 sky130_fd_sc_hd__nand2_2 _26679_ (.A(_09434_),
    .B(_09689_),
    .Y(_09700_));
 sky130_fd_sc_hd__buf_1 _26680_ (.A(_10130_),
    .X(_09701_));
 sky130_fd_sc_hd__buf_1 _26681_ (.A(_09701_),
    .X(_09702_));
 sky130_fd_sc_hd__o211a_2 _26682_ (.A1(\decode.regfile.registers_17[27] ),
    .A2(_09692_),
    .B1(_09700_),
    .C1(_09702_),
    .X(_02826_));
 sky130_fd_sc_hd__nand2_2 _26683_ (.A(_09436_),
    .B(_09664_),
    .Y(_09703_));
 sky130_fd_sc_hd__o211a_2 _26684_ (.A1(\decode.regfile.registers_17[28] ),
    .A2(_09692_),
    .B1(_09703_),
    .C1(_09702_),
    .X(_02827_));
 sky130_fd_sc_hd__nand2_2 _26685_ (.A(_09438_),
    .B(_09664_),
    .Y(_09704_));
 sky130_fd_sc_hd__o211a_2 _26686_ (.A1(\decode.regfile.registers_17[29] ),
    .A2(_09692_),
    .B1(_09704_),
    .C1(_09702_),
    .X(_02828_));
 sky130_fd_sc_hd__nand2_2 _26687_ (.A(_09441_),
    .B(_09664_),
    .Y(_09705_));
 sky130_fd_sc_hd__o211a_2 _26688_ (.A1(\decode.regfile.registers_17[30] ),
    .A2(_09666_),
    .B1(_09705_),
    .C1(_09702_),
    .X(_02829_));
 sky130_fd_sc_hd__nand2_2 _26689_ (.A(_09443_),
    .B(_09664_),
    .Y(_09706_));
 sky130_fd_sc_hd__o211a_2 _26690_ (.A1(\decode.regfile.registers_17[31] ),
    .A2(_09666_),
    .B1(_09706_),
    .C1(_09702_),
    .X(_02830_));
 sky130_fd_sc_hd__and3_2 _26691_ (.A(_09932_),
    .B(_10149_),
    .C(_03672_),
    .X(_09707_));
 sky130_fd_sc_hd__buf_1 _26692_ (.A(_09707_),
    .X(_09708_));
 sky130_fd_sc_hd__buf_1 _26693_ (.A(_09708_),
    .X(_09709_));
 sky130_fd_sc_hd__buf_1 _26694_ (.A(_09708_),
    .X(_09710_));
 sky130_fd_sc_hd__nand2_2 _26695_ (.A(_10245_),
    .B(_09710_),
    .Y(_09711_));
 sky130_fd_sc_hd__o211a_2 _26696_ (.A1(\decode.regfile.registers_18[0] ),
    .A2(_09709_),
    .B1(_09711_),
    .C1(_09702_),
    .X(_02831_));
 sky130_fd_sc_hd__nand2_2 _26697_ (.A(_09450_),
    .B(_09710_),
    .Y(_09712_));
 sky130_fd_sc_hd__o211a_2 _26698_ (.A1(\decode.regfile.registers_18[1] ),
    .A2(_09709_),
    .B1(_09712_),
    .C1(_09702_),
    .X(_02832_));
 sky130_fd_sc_hd__nand2_2 _26699_ (.A(_09377_),
    .B(_09710_),
    .Y(_09713_));
 sky130_fd_sc_hd__o211a_2 _26700_ (.A1(\decode.regfile.registers_18[2] ),
    .A2(_09709_),
    .B1(_09713_),
    .C1(_09702_),
    .X(_02833_));
 sky130_fd_sc_hd__nand2_2 _26701_ (.A(_09379_),
    .B(_09710_),
    .Y(_09714_));
 sky130_fd_sc_hd__o211a_2 _26702_ (.A1(\decode.regfile.registers_18[3] ),
    .A2(_09709_),
    .B1(_09714_),
    .C1(_09702_),
    .X(_02834_));
 sky130_fd_sc_hd__nand2_2 _26703_ (.A(_09381_),
    .B(_09710_),
    .Y(_09715_));
 sky130_fd_sc_hd__o211a_2 _26704_ (.A1(\decode.regfile.registers_18[4] ),
    .A2(_09709_),
    .B1(_09715_),
    .C1(_09702_),
    .X(_02835_));
 sky130_fd_sc_hd__nand2_2 _26705_ (.A(_09383_),
    .B(_09710_),
    .Y(_09716_));
 sky130_fd_sc_hd__buf_1 _26706_ (.A(_09701_),
    .X(_09717_));
 sky130_fd_sc_hd__o211a_2 _26707_ (.A1(\decode.regfile.registers_18[5] ),
    .A2(_09709_),
    .B1(_09716_),
    .C1(_09717_),
    .X(_02836_));
 sky130_fd_sc_hd__nand2_2 _26708_ (.A(_09385_),
    .B(_09710_),
    .Y(_09718_));
 sky130_fd_sc_hd__o211a_2 _26709_ (.A1(\decode.regfile.registers_18[6] ),
    .A2(_09709_),
    .B1(_09718_),
    .C1(_09717_),
    .X(_02837_));
 sky130_fd_sc_hd__nand2_2 _26710_ (.A(_09387_),
    .B(_09710_),
    .Y(_09719_));
 sky130_fd_sc_hd__o211a_2 _26711_ (.A1(\decode.regfile.registers_18[7] ),
    .A2(_09709_),
    .B1(_09719_),
    .C1(_09717_),
    .X(_02838_));
 sky130_fd_sc_hd__buf_1 _26712_ (.A(_09708_),
    .X(_09720_));
 sky130_fd_sc_hd__nand2_2 _26713_ (.A(_09389_),
    .B(_09720_),
    .Y(_09721_));
 sky130_fd_sc_hd__o211a_2 _26714_ (.A1(\decode.regfile.registers_18[8] ),
    .A2(_09709_),
    .B1(_09721_),
    .C1(_09717_),
    .X(_02839_));
 sky130_fd_sc_hd__nand2_2 _26715_ (.A(_09392_),
    .B(_09720_),
    .Y(_09722_));
 sky130_fd_sc_hd__o211a_2 _26716_ (.A1(\decode.regfile.registers_18[9] ),
    .A2(_09709_),
    .B1(_09722_),
    .C1(_09717_),
    .X(_02840_));
 sky130_fd_sc_hd__buf_1 _26717_ (.A(_09708_),
    .X(_09723_));
 sky130_fd_sc_hd__nand2_2 _26718_ (.A(_09396_),
    .B(_09720_),
    .Y(_09724_));
 sky130_fd_sc_hd__o211a_2 _26719_ (.A1(\decode.regfile.registers_18[10] ),
    .A2(_09723_),
    .B1(_09724_),
    .C1(_09717_),
    .X(_02841_));
 sky130_fd_sc_hd__nand2_2 _26720_ (.A(_09398_),
    .B(_09720_),
    .Y(_09725_));
 sky130_fd_sc_hd__o211a_2 _26721_ (.A1(\decode.regfile.registers_18[11] ),
    .A2(_09723_),
    .B1(_09725_),
    .C1(_09717_),
    .X(_02842_));
 sky130_fd_sc_hd__nand2_2 _26722_ (.A(_09400_),
    .B(_09720_),
    .Y(_09726_));
 sky130_fd_sc_hd__o211a_2 _26723_ (.A1(\decode.regfile.registers_18[12] ),
    .A2(_09723_),
    .B1(_09726_),
    .C1(_09717_),
    .X(_02843_));
 sky130_fd_sc_hd__nand2_2 _26724_ (.A(_09402_),
    .B(_09720_),
    .Y(_09727_));
 sky130_fd_sc_hd__o211a_2 _26725_ (.A1(\decode.regfile.registers_18[13] ),
    .A2(_09723_),
    .B1(_09727_),
    .C1(_09717_),
    .X(_02844_));
 sky130_fd_sc_hd__nand2_2 _26726_ (.A(_09404_),
    .B(_09720_),
    .Y(_09728_));
 sky130_fd_sc_hd__o211a_2 _26727_ (.A1(\decode.regfile.registers_18[14] ),
    .A2(_09723_),
    .B1(_09728_),
    .C1(_09717_),
    .X(_02845_));
 sky130_fd_sc_hd__nand2_2 _26728_ (.A(_09406_),
    .B(_09720_),
    .Y(_09729_));
 sky130_fd_sc_hd__buf_1 _26729_ (.A(_09701_),
    .X(_09730_));
 sky130_fd_sc_hd__o211a_2 _26730_ (.A1(\decode.regfile.registers_18[15] ),
    .A2(_09723_),
    .B1(_09729_),
    .C1(_09730_),
    .X(_02846_));
 sky130_fd_sc_hd__nand2_2 _26731_ (.A(_09408_),
    .B(_09720_),
    .Y(_09731_));
 sky130_fd_sc_hd__o211a_2 _26732_ (.A1(\decode.regfile.registers_18[16] ),
    .A2(_09723_),
    .B1(_09731_),
    .C1(_09730_),
    .X(_02847_));
 sky130_fd_sc_hd__nand2_2 _26733_ (.A(_09410_),
    .B(_09720_),
    .Y(_09732_));
 sky130_fd_sc_hd__o211a_2 _26734_ (.A1(\decode.regfile.registers_18[17] ),
    .A2(_09723_),
    .B1(_09732_),
    .C1(_09730_),
    .X(_02848_));
 sky130_fd_sc_hd__buf_1 _26735_ (.A(_09708_),
    .X(_09733_));
 sky130_fd_sc_hd__nand2_2 _26736_ (.A(_09412_),
    .B(_09733_),
    .Y(_09734_));
 sky130_fd_sc_hd__o211a_2 _26737_ (.A1(\decode.regfile.registers_18[18] ),
    .A2(_09723_),
    .B1(_09734_),
    .C1(_09730_),
    .X(_02849_));
 sky130_fd_sc_hd__nand2_2 _26738_ (.A(_09415_),
    .B(_09733_),
    .Y(_09735_));
 sky130_fd_sc_hd__o211a_2 _26739_ (.A1(\decode.regfile.registers_18[19] ),
    .A2(_09723_),
    .B1(_09735_),
    .C1(_09730_),
    .X(_02850_));
 sky130_fd_sc_hd__buf_1 _26740_ (.A(_09708_),
    .X(_09736_));
 sky130_fd_sc_hd__nand2_2 _26741_ (.A(_09420_),
    .B(_09733_),
    .Y(_09737_));
 sky130_fd_sc_hd__o211a_2 _26742_ (.A1(\decode.regfile.registers_18[20] ),
    .A2(_09736_),
    .B1(_09737_),
    .C1(_09730_),
    .X(_02851_));
 sky130_fd_sc_hd__nand2_2 _26743_ (.A(_09422_),
    .B(_09733_),
    .Y(_09738_));
 sky130_fd_sc_hd__o211a_2 _26744_ (.A1(\decode.regfile.registers_18[21] ),
    .A2(_09736_),
    .B1(_09738_),
    .C1(_09730_),
    .X(_02852_));
 sky130_fd_sc_hd__nand2_2 _26745_ (.A(_09424_),
    .B(_09733_),
    .Y(_09739_));
 sky130_fd_sc_hd__o211a_2 _26746_ (.A1(\decode.regfile.registers_18[22] ),
    .A2(_09736_),
    .B1(_09739_),
    .C1(_09730_),
    .X(_02853_));
 sky130_fd_sc_hd__nand2_2 _26747_ (.A(_09426_),
    .B(_09733_),
    .Y(_09740_));
 sky130_fd_sc_hd__o211a_2 _26748_ (.A1(\decode.regfile.registers_18[23] ),
    .A2(_09736_),
    .B1(_09740_),
    .C1(_09730_),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_2 _26749_ (.A(_09428_),
    .B(_09733_),
    .Y(_09741_));
 sky130_fd_sc_hd__o211a_2 _26750_ (.A1(\decode.regfile.registers_18[24] ),
    .A2(_09736_),
    .B1(_09741_),
    .C1(_09730_),
    .X(_02855_));
 sky130_fd_sc_hd__nand2_2 _26751_ (.A(_09430_),
    .B(_09733_),
    .Y(_09742_));
 sky130_fd_sc_hd__buf_1 _26752_ (.A(_09701_),
    .X(_09743_));
 sky130_fd_sc_hd__o211a_2 _26753_ (.A1(\decode.regfile.registers_18[25] ),
    .A2(_09736_),
    .B1(_09742_),
    .C1(_09743_),
    .X(_02856_));
 sky130_fd_sc_hd__nand2_2 _26754_ (.A(_09432_),
    .B(_09733_),
    .Y(_09744_));
 sky130_fd_sc_hd__o211a_2 _26755_ (.A1(\decode.regfile.registers_18[26] ),
    .A2(_09736_),
    .B1(_09744_),
    .C1(_09743_),
    .X(_02857_));
 sky130_fd_sc_hd__nand2_2 _26756_ (.A(_09434_),
    .B(_09733_),
    .Y(_09745_));
 sky130_fd_sc_hd__o211a_2 _26757_ (.A1(\decode.regfile.registers_18[27] ),
    .A2(_09736_),
    .B1(_09745_),
    .C1(_09743_),
    .X(_02858_));
 sky130_fd_sc_hd__nand2_2 _26758_ (.A(_09436_),
    .B(_09708_),
    .Y(_09746_));
 sky130_fd_sc_hd__o211a_2 _26759_ (.A1(\decode.regfile.registers_18[28] ),
    .A2(_09736_),
    .B1(_09746_),
    .C1(_09743_),
    .X(_02859_));
 sky130_fd_sc_hd__nand2_2 _26760_ (.A(_09438_),
    .B(_09708_),
    .Y(_09747_));
 sky130_fd_sc_hd__o211a_2 _26761_ (.A1(\decode.regfile.registers_18[29] ),
    .A2(_09736_),
    .B1(_09747_),
    .C1(_09743_),
    .X(_02860_));
 sky130_fd_sc_hd__nand2_2 _26762_ (.A(_09441_),
    .B(_09708_),
    .Y(_09748_));
 sky130_fd_sc_hd__o211a_2 _26763_ (.A1(\decode.regfile.registers_18[30] ),
    .A2(_09710_),
    .B1(_09748_),
    .C1(_09743_),
    .X(_02861_));
 sky130_fd_sc_hd__nand2_2 _26764_ (.A(_09443_),
    .B(_09708_),
    .Y(_09749_));
 sky130_fd_sc_hd__o211a_2 _26765_ (.A1(\decode.regfile.registers_18[31] ),
    .A2(_09710_),
    .B1(_09749_),
    .C1(_09743_),
    .X(_02862_));
 sky130_fd_sc_hd__and3_2 _26766_ (.A(_10149_),
    .B(_10150_),
    .C(_03672_),
    .X(_09750_));
 sky130_fd_sc_hd__buf_1 _26767_ (.A(_09750_),
    .X(_09751_));
 sky130_fd_sc_hd__buf_1 _26768_ (.A(_09751_),
    .X(_09752_));
 sky130_fd_sc_hd__buf_1 _26769_ (.A(_09751_),
    .X(_09753_));
 sky130_fd_sc_hd__nand2_2 _26770_ (.A(_10245_),
    .B(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__o211a_2 _26771_ (.A1(\decode.regfile.registers_19[0] ),
    .A2(_09752_),
    .B1(_09754_),
    .C1(_09743_),
    .X(_02863_));
 sky130_fd_sc_hd__nand2_2 _26772_ (.A(_09450_),
    .B(_09753_),
    .Y(_09755_));
 sky130_fd_sc_hd__o211a_2 _26773_ (.A1(\decode.regfile.registers_19[1] ),
    .A2(_09752_),
    .B1(_09755_),
    .C1(_09743_),
    .X(_02864_));
 sky130_fd_sc_hd__nand2_2 _26774_ (.A(_09377_),
    .B(_09753_),
    .Y(_09756_));
 sky130_fd_sc_hd__o211a_2 _26775_ (.A1(\decode.regfile.registers_19[2] ),
    .A2(_09752_),
    .B1(_09756_),
    .C1(_09743_),
    .X(_02865_));
 sky130_fd_sc_hd__nand2_2 _26776_ (.A(_09379_),
    .B(_09753_),
    .Y(_09757_));
 sky130_fd_sc_hd__buf_1 _26777_ (.A(_09701_),
    .X(_09758_));
 sky130_fd_sc_hd__o211a_2 _26778_ (.A1(\decode.regfile.registers_19[3] ),
    .A2(_09752_),
    .B1(_09757_),
    .C1(_09758_),
    .X(_02866_));
 sky130_fd_sc_hd__nand2_2 _26779_ (.A(_09381_),
    .B(_09753_),
    .Y(_09759_));
 sky130_fd_sc_hd__o211a_2 _26780_ (.A1(\decode.regfile.registers_19[4] ),
    .A2(_09752_),
    .B1(_09759_),
    .C1(_09758_),
    .X(_02867_));
 sky130_fd_sc_hd__nand2_2 _26781_ (.A(_09383_),
    .B(_09753_),
    .Y(_09760_));
 sky130_fd_sc_hd__o211a_2 _26782_ (.A1(\decode.regfile.registers_19[5] ),
    .A2(_09752_),
    .B1(_09760_),
    .C1(_09758_),
    .X(_02868_));
 sky130_fd_sc_hd__nand2_2 _26783_ (.A(_09385_),
    .B(_09753_),
    .Y(_09761_));
 sky130_fd_sc_hd__o211a_2 _26784_ (.A1(\decode.regfile.registers_19[6] ),
    .A2(_09752_),
    .B1(_09761_),
    .C1(_09758_),
    .X(_02869_));
 sky130_fd_sc_hd__nand2_2 _26785_ (.A(_09387_),
    .B(_09753_),
    .Y(_09762_));
 sky130_fd_sc_hd__o211a_2 _26786_ (.A1(\decode.regfile.registers_19[7] ),
    .A2(_09752_),
    .B1(_09762_),
    .C1(_09758_),
    .X(_02870_));
 sky130_fd_sc_hd__buf_1 _26787_ (.A(_09751_),
    .X(_09763_));
 sky130_fd_sc_hd__nand2_2 _26788_ (.A(_09389_),
    .B(_09763_),
    .Y(_09764_));
 sky130_fd_sc_hd__o211a_2 _26789_ (.A1(\decode.regfile.registers_19[8] ),
    .A2(_09752_),
    .B1(_09764_),
    .C1(_09758_),
    .X(_02871_));
 sky130_fd_sc_hd__nand2_2 _26790_ (.A(_09392_),
    .B(_09763_),
    .Y(_09765_));
 sky130_fd_sc_hd__o211a_2 _26791_ (.A1(\decode.regfile.registers_19[9] ),
    .A2(_09752_),
    .B1(_09765_),
    .C1(_09758_),
    .X(_02872_));
 sky130_fd_sc_hd__buf_1 _26792_ (.A(_09751_),
    .X(_09766_));
 sky130_fd_sc_hd__nand2_2 _26793_ (.A(_09396_),
    .B(_09763_),
    .Y(_09767_));
 sky130_fd_sc_hd__o211a_2 _26794_ (.A1(\decode.regfile.registers_19[10] ),
    .A2(_09766_),
    .B1(_09767_),
    .C1(_09758_),
    .X(_02873_));
 sky130_fd_sc_hd__nand2_2 _26795_ (.A(_09398_),
    .B(_09763_),
    .Y(_09768_));
 sky130_fd_sc_hd__o211a_2 _26796_ (.A1(\decode.regfile.registers_19[11] ),
    .A2(_09766_),
    .B1(_09768_),
    .C1(_09758_),
    .X(_02874_));
 sky130_fd_sc_hd__nand2_2 _26797_ (.A(_09400_),
    .B(_09763_),
    .Y(_09769_));
 sky130_fd_sc_hd__o211a_2 _26798_ (.A1(\decode.regfile.registers_19[12] ),
    .A2(_09766_),
    .B1(_09769_),
    .C1(_09758_),
    .X(_02875_));
 sky130_fd_sc_hd__nand2_2 _26799_ (.A(_09402_),
    .B(_09763_),
    .Y(_09770_));
 sky130_fd_sc_hd__buf_1 _26800_ (.A(_09701_),
    .X(_09771_));
 sky130_fd_sc_hd__o211a_2 _26801_ (.A1(\decode.regfile.registers_19[13] ),
    .A2(_09766_),
    .B1(_09770_),
    .C1(_09771_),
    .X(_02876_));
 sky130_fd_sc_hd__nand2_2 _26802_ (.A(_09404_),
    .B(_09763_),
    .Y(_09772_));
 sky130_fd_sc_hd__o211a_2 _26803_ (.A1(\decode.regfile.registers_19[14] ),
    .A2(_09766_),
    .B1(_09772_),
    .C1(_09771_),
    .X(_02877_));
 sky130_fd_sc_hd__nand2_2 _26804_ (.A(_09406_),
    .B(_09763_),
    .Y(_09773_));
 sky130_fd_sc_hd__o211a_2 _26805_ (.A1(\decode.regfile.registers_19[15] ),
    .A2(_09766_),
    .B1(_09773_),
    .C1(_09771_),
    .X(_02878_));
 sky130_fd_sc_hd__nand2_2 _26806_ (.A(_09408_),
    .B(_09763_),
    .Y(_09774_));
 sky130_fd_sc_hd__o211a_2 _26807_ (.A1(\decode.regfile.registers_19[16] ),
    .A2(_09766_),
    .B1(_09774_),
    .C1(_09771_),
    .X(_02879_));
 sky130_fd_sc_hd__nand2_2 _26808_ (.A(_09410_),
    .B(_09763_),
    .Y(_09775_));
 sky130_fd_sc_hd__o211a_2 _26809_ (.A1(\decode.regfile.registers_19[17] ),
    .A2(_09766_),
    .B1(_09775_),
    .C1(_09771_),
    .X(_02880_));
 sky130_fd_sc_hd__buf_1 _26810_ (.A(_09751_),
    .X(_09776_));
 sky130_fd_sc_hd__nand2_2 _26811_ (.A(_09412_),
    .B(_09776_),
    .Y(_09777_));
 sky130_fd_sc_hd__o211a_2 _26812_ (.A1(\decode.regfile.registers_19[18] ),
    .A2(_09766_),
    .B1(_09777_),
    .C1(_09771_),
    .X(_02881_));
 sky130_fd_sc_hd__nand2_2 _26813_ (.A(_09415_),
    .B(_09776_),
    .Y(_09778_));
 sky130_fd_sc_hd__o211a_2 _26814_ (.A1(\decode.regfile.registers_19[19] ),
    .A2(_09766_),
    .B1(_09778_),
    .C1(_09771_),
    .X(_02882_));
 sky130_fd_sc_hd__buf_1 _26815_ (.A(_09751_),
    .X(_09779_));
 sky130_fd_sc_hd__nand2_2 _26816_ (.A(_09420_),
    .B(_09776_),
    .Y(_09780_));
 sky130_fd_sc_hd__o211a_2 _26817_ (.A1(\decode.regfile.registers_19[20] ),
    .A2(_09779_),
    .B1(_09780_),
    .C1(_09771_),
    .X(_02883_));
 sky130_fd_sc_hd__nand2_2 _26818_ (.A(_09422_),
    .B(_09776_),
    .Y(_09781_));
 sky130_fd_sc_hd__o211a_2 _26819_ (.A1(\decode.regfile.registers_19[21] ),
    .A2(_09779_),
    .B1(_09781_),
    .C1(_09771_),
    .X(_02884_));
 sky130_fd_sc_hd__nand2_2 _26820_ (.A(_09424_),
    .B(_09776_),
    .Y(_09782_));
 sky130_fd_sc_hd__o211a_2 _26821_ (.A1(\decode.regfile.registers_19[22] ),
    .A2(_09779_),
    .B1(_09782_),
    .C1(_09771_),
    .X(_02885_));
 sky130_fd_sc_hd__nand2_2 _26822_ (.A(_09426_),
    .B(_09776_),
    .Y(_09783_));
 sky130_fd_sc_hd__buf_1 _26823_ (.A(_09701_),
    .X(_09784_));
 sky130_fd_sc_hd__o211a_2 _26824_ (.A1(\decode.regfile.registers_19[23] ),
    .A2(_09779_),
    .B1(_09783_),
    .C1(_09784_),
    .X(_02886_));
 sky130_fd_sc_hd__nand2_2 _26825_ (.A(_09428_),
    .B(_09776_),
    .Y(_09785_));
 sky130_fd_sc_hd__o211a_2 _26826_ (.A1(\decode.regfile.registers_19[24] ),
    .A2(_09779_),
    .B1(_09785_),
    .C1(_09784_),
    .X(_02887_));
 sky130_fd_sc_hd__nand2_2 _26827_ (.A(_09430_),
    .B(_09776_),
    .Y(_09786_));
 sky130_fd_sc_hd__o211a_2 _26828_ (.A1(\decode.regfile.registers_19[25] ),
    .A2(_09779_),
    .B1(_09786_),
    .C1(_09784_),
    .X(_02888_));
 sky130_fd_sc_hd__nand2_2 _26829_ (.A(_09432_),
    .B(_09776_),
    .Y(_09787_));
 sky130_fd_sc_hd__o211a_2 _26830_ (.A1(\decode.regfile.registers_19[26] ),
    .A2(_09779_),
    .B1(_09787_),
    .C1(_09784_),
    .X(_02889_));
 sky130_fd_sc_hd__nand2_2 _26831_ (.A(_09434_),
    .B(_09776_),
    .Y(_09788_));
 sky130_fd_sc_hd__o211a_2 _26832_ (.A1(\decode.regfile.registers_19[27] ),
    .A2(_09779_),
    .B1(_09788_),
    .C1(_09784_),
    .X(_02890_));
 sky130_fd_sc_hd__nand2_2 _26833_ (.A(_09436_),
    .B(_09751_),
    .Y(_09789_));
 sky130_fd_sc_hd__o211a_2 _26834_ (.A1(\decode.regfile.registers_19[28] ),
    .A2(_09779_),
    .B1(_09789_),
    .C1(_09784_),
    .X(_02891_));
 sky130_fd_sc_hd__nand2_2 _26835_ (.A(_09438_),
    .B(_09751_),
    .Y(_09790_));
 sky130_fd_sc_hd__o211a_2 _26836_ (.A1(\decode.regfile.registers_19[29] ),
    .A2(_09779_),
    .B1(_09790_),
    .C1(_09784_),
    .X(_02892_));
 sky130_fd_sc_hd__nand2_2 _26837_ (.A(_09441_),
    .B(_09751_),
    .Y(_09791_));
 sky130_fd_sc_hd__o211a_2 _26838_ (.A1(\decode.regfile.registers_19[30] ),
    .A2(_09753_),
    .B1(_09791_),
    .C1(_09784_),
    .X(_02893_));
 sky130_fd_sc_hd__nand2_2 _26839_ (.A(_09443_),
    .B(_09751_),
    .Y(_09792_));
 sky130_fd_sc_hd__o211a_2 _26840_ (.A1(\decode.regfile.registers_19[31] ),
    .A2(_09753_),
    .B1(_09792_),
    .C1(_09784_),
    .X(_02894_));
 sky130_fd_sc_hd__and4_2 _26841_ (.A(_09929_),
    .B(_10149_),
    .C(_10196_),
    .D(_09935_),
    .X(_09793_));
 sky130_fd_sc_hd__buf_1 _26842_ (.A(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__buf_1 _26843_ (.A(_09794_),
    .X(_09795_));
 sky130_fd_sc_hd__buf_1 _26844_ (.A(_09794_),
    .X(_09796_));
 sky130_fd_sc_hd__nand2_2 _26845_ (.A(_10245_),
    .B(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__o211a_2 _26846_ (.A1(\decode.regfile.registers_20[0] ),
    .A2(_09795_),
    .B1(_09797_),
    .C1(_09784_),
    .X(_02895_));
 sky130_fd_sc_hd__nand2_2 _26847_ (.A(_09450_),
    .B(_09796_),
    .Y(_09798_));
 sky130_fd_sc_hd__buf_1 _26848_ (.A(_09701_),
    .X(_09799_));
 sky130_fd_sc_hd__o211a_2 _26849_ (.A1(\decode.regfile.registers_20[1] ),
    .A2(_09795_),
    .B1(_09798_),
    .C1(_09799_),
    .X(_02896_));
 sky130_fd_sc_hd__nand2_2 _26850_ (.A(_09377_),
    .B(_09796_),
    .Y(_09800_));
 sky130_fd_sc_hd__o211a_2 _26851_ (.A1(\decode.regfile.registers_20[2] ),
    .A2(_09795_),
    .B1(_09800_),
    .C1(_09799_),
    .X(_02897_));
 sky130_fd_sc_hd__nand2_2 _26852_ (.A(_09379_),
    .B(_09796_),
    .Y(_09801_));
 sky130_fd_sc_hd__o211a_2 _26853_ (.A1(\decode.regfile.registers_20[3] ),
    .A2(_09795_),
    .B1(_09801_),
    .C1(_09799_),
    .X(_02898_));
 sky130_fd_sc_hd__nand2_2 _26854_ (.A(_09381_),
    .B(_09796_),
    .Y(_09802_));
 sky130_fd_sc_hd__o211a_2 _26855_ (.A1(\decode.regfile.registers_20[4] ),
    .A2(_09795_),
    .B1(_09802_),
    .C1(_09799_),
    .X(_02899_));
 sky130_fd_sc_hd__nand2_2 _26856_ (.A(_09383_),
    .B(_09796_),
    .Y(_09803_));
 sky130_fd_sc_hd__o211a_2 _26857_ (.A1(\decode.regfile.registers_20[5] ),
    .A2(_09795_),
    .B1(_09803_),
    .C1(_09799_),
    .X(_02900_));
 sky130_fd_sc_hd__nand2_2 _26858_ (.A(_09385_),
    .B(_09796_),
    .Y(_09804_));
 sky130_fd_sc_hd__o211a_2 _26859_ (.A1(\decode.regfile.registers_20[6] ),
    .A2(_09795_),
    .B1(_09804_),
    .C1(_09799_),
    .X(_02901_));
 sky130_fd_sc_hd__nand2_2 _26860_ (.A(_09387_),
    .B(_09796_),
    .Y(_09805_));
 sky130_fd_sc_hd__o211a_2 _26861_ (.A1(\decode.regfile.registers_20[7] ),
    .A2(_09795_),
    .B1(_09805_),
    .C1(_09799_),
    .X(_02902_));
 sky130_fd_sc_hd__buf_1 _26862_ (.A(_09794_),
    .X(_09806_));
 sky130_fd_sc_hd__nand2_2 _26863_ (.A(_09389_),
    .B(_09806_),
    .Y(_09807_));
 sky130_fd_sc_hd__o211a_2 _26864_ (.A1(\decode.regfile.registers_20[8] ),
    .A2(_09795_),
    .B1(_09807_),
    .C1(_09799_),
    .X(_02903_));
 sky130_fd_sc_hd__nand2_2 _26865_ (.A(_09392_),
    .B(_09806_),
    .Y(_09808_));
 sky130_fd_sc_hd__o211a_2 _26866_ (.A1(\decode.regfile.registers_20[9] ),
    .A2(_09795_),
    .B1(_09808_),
    .C1(_09799_),
    .X(_02904_));
 sky130_fd_sc_hd__buf_1 _26867_ (.A(_09794_),
    .X(_09809_));
 sky130_fd_sc_hd__nand2_2 _26868_ (.A(_09396_),
    .B(_09806_),
    .Y(_09810_));
 sky130_fd_sc_hd__o211a_2 _26869_ (.A1(\decode.regfile.registers_20[10] ),
    .A2(_09809_),
    .B1(_09810_),
    .C1(_09799_),
    .X(_02905_));
 sky130_fd_sc_hd__nand2_2 _26870_ (.A(_09398_),
    .B(_09806_),
    .Y(_09811_));
 sky130_fd_sc_hd__buf_1 _26871_ (.A(_09701_),
    .X(_09812_));
 sky130_fd_sc_hd__o211a_2 _26872_ (.A1(\decode.regfile.registers_20[11] ),
    .A2(_09809_),
    .B1(_09811_),
    .C1(_09812_),
    .X(_02906_));
 sky130_fd_sc_hd__nand2_2 _26873_ (.A(_09400_),
    .B(_09806_),
    .Y(_09813_));
 sky130_fd_sc_hd__o211a_2 _26874_ (.A1(\decode.regfile.registers_20[12] ),
    .A2(_09809_),
    .B1(_09813_),
    .C1(_09812_),
    .X(_02907_));
 sky130_fd_sc_hd__nand2_2 _26875_ (.A(_09402_),
    .B(_09806_),
    .Y(_09814_));
 sky130_fd_sc_hd__o211a_2 _26876_ (.A1(\decode.regfile.registers_20[13] ),
    .A2(_09809_),
    .B1(_09814_),
    .C1(_09812_),
    .X(_02908_));
 sky130_fd_sc_hd__nand2_2 _26877_ (.A(_09404_),
    .B(_09806_),
    .Y(_09815_));
 sky130_fd_sc_hd__o211a_2 _26878_ (.A1(\decode.regfile.registers_20[14] ),
    .A2(_09809_),
    .B1(_09815_),
    .C1(_09812_),
    .X(_02909_));
 sky130_fd_sc_hd__nand2_2 _26879_ (.A(_09406_),
    .B(_09806_),
    .Y(_09816_));
 sky130_fd_sc_hd__o211a_2 _26880_ (.A1(\decode.regfile.registers_20[15] ),
    .A2(_09809_),
    .B1(_09816_),
    .C1(_09812_),
    .X(_02910_));
 sky130_fd_sc_hd__nand2_2 _26881_ (.A(_09408_),
    .B(_09806_),
    .Y(_09817_));
 sky130_fd_sc_hd__o211a_2 _26882_ (.A1(\decode.regfile.registers_20[16] ),
    .A2(_09809_),
    .B1(_09817_),
    .C1(_09812_),
    .X(_02911_));
 sky130_fd_sc_hd__nand2_2 _26883_ (.A(_09410_),
    .B(_09806_),
    .Y(_09818_));
 sky130_fd_sc_hd__o211a_2 _26884_ (.A1(\decode.regfile.registers_20[17] ),
    .A2(_09809_),
    .B1(_09818_),
    .C1(_09812_),
    .X(_02912_));
 sky130_fd_sc_hd__buf_1 _26885_ (.A(_09794_),
    .X(_09819_));
 sky130_fd_sc_hd__nand2_2 _26886_ (.A(_09412_),
    .B(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__o211a_2 _26887_ (.A1(\decode.regfile.registers_20[18] ),
    .A2(_09809_),
    .B1(_09820_),
    .C1(_09812_),
    .X(_02913_));
 sky130_fd_sc_hd__nand2_2 _26888_ (.A(_09415_),
    .B(_09819_),
    .Y(_09821_));
 sky130_fd_sc_hd__o211a_2 _26889_ (.A1(\decode.regfile.registers_20[19] ),
    .A2(_09809_),
    .B1(_09821_),
    .C1(_09812_),
    .X(_02914_));
 sky130_fd_sc_hd__buf_1 _26890_ (.A(_09794_),
    .X(_09822_));
 sky130_fd_sc_hd__nand2_2 _26891_ (.A(_09420_),
    .B(_09819_),
    .Y(_09823_));
 sky130_fd_sc_hd__o211a_2 _26892_ (.A1(\decode.regfile.registers_20[20] ),
    .A2(_09822_),
    .B1(_09823_),
    .C1(_09812_),
    .X(_02915_));
 sky130_fd_sc_hd__nand2_2 _26893_ (.A(_09422_),
    .B(_09819_),
    .Y(_09824_));
 sky130_fd_sc_hd__buf_1 _26894_ (.A(_09701_),
    .X(_09825_));
 sky130_fd_sc_hd__o211a_2 _26895_ (.A1(\decode.regfile.registers_20[21] ),
    .A2(_09822_),
    .B1(_09824_),
    .C1(_09825_),
    .X(_02916_));
 sky130_fd_sc_hd__nand2_2 _26896_ (.A(_09424_),
    .B(_09819_),
    .Y(_09826_));
 sky130_fd_sc_hd__o211a_2 _26897_ (.A1(\decode.regfile.registers_20[22] ),
    .A2(_09822_),
    .B1(_09826_),
    .C1(_09825_),
    .X(_02917_));
 sky130_fd_sc_hd__nand2_2 _26898_ (.A(_09426_),
    .B(_09819_),
    .Y(_09827_));
 sky130_fd_sc_hd__o211a_2 _26899_ (.A1(\decode.regfile.registers_20[23] ),
    .A2(_09822_),
    .B1(_09827_),
    .C1(_09825_),
    .X(_02918_));
 sky130_fd_sc_hd__nand2_2 _26900_ (.A(_09428_),
    .B(_09819_),
    .Y(_09828_));
 sky130_fd_sc_hd__o211a_2 _26901_ (.A1(\decode.regfile.registers_20[24] ),
    .A2(_09822_),
    .B1(_09828_),
    .C1(_09825_),
    .X(_02919_));
 sky130_fd_sc_hd__nand2_2 _26902_ (.A(_09430_),
    .B(_09819_),
    .Y(_09829_));
 sky130_fd_sc_hd__o211a_2 _26903_ (.A1(\decode.regfile.registers_20[25] ),
    .A2(_09822_),
    .B1(_09829_),
    .C1(_09825_),
    .X(_02920_));
 sky130_fd_sc_hd__nand2_2 _26904_ (.A(_09432_),
    .B(_09819_),
    .Y(_09830_));
 sky130_fd_sc_hd__o211a_2 _26905_ (.A1(\decode.regfile.registers_20[26] ),
    .A2(_09822_),
    .B1(_09830_),
    .C1(_09825_),
    .X(_02921_));
 sky130_fd_sc_hd__nand2_2 _26906_ (.A(_09434_),
    .B(_09819_),
    .Y(_09831_));
 sky130_fd_sc_hd__o211a_2 _26907_ (.A1(\decode.regfile.registers_20[27] ),
    .A2(_09822_),
    .B1(_09831_),
    .C1(_09825_),
    .X(_02922_));
 sky130_fd_sc_hd__nand2_2 _26908_ (.A(_09436_),
    .B(_09794_),
    .Y(_09832_));
 sky130_fd_sc_hd__o211a_2 _26909_ (.A1(\decode.regfile.registers_20[28] ),
    .A2(_09822_),
    .B1(_09832_),
    .C1(_09825_),
    .X(_02923_));
 sky130_fd_sc_hd__nand2_2 _26910_ (.A(_09438_),
    .B(_09794_),
    .Y(_09833_));
 sky130_fd_sc_hd__o211a_2 _26911_ (.A1(\decode.regfile.registers_20[29] ),
    .A2(_09822_),
    .B1(_09833_),
    .C1(_09825_),
    .X(_02924_));
 sky130_fd_sc_hd__nand2_2 _26912_ (.A(_09441_),
    .B(_09794_),
    .Y(_09834_));
 sky130_fd_sc_hd__o211a_2 _26913_ (.A1(\decode.regfile.registers_20[30] ),
    .A2(_09796_),
    .B1(_09834_),
    .C1(_09825_),
    .X(_02925_));
 sky130_fd_sc_hd__nand2_2 _26914_ (.A(_09443_),
    .B(_09794_),
    .Y(_09835_));
 sky130_fd_sc_hd__buf_1 _26915_ (.A(_09956_),
    .X(_09836_));
 sky130_fd_sc_hd__o211a_2 _26916_ (.A1(\decode.regfile.registers_20[31] ),
    .A2(_09796_),
    .B1(_09835_),
    .C1(_09836_),
    .X(_02926_));
 sky130_fd_sc_hd__and4_2 _26917_ (.A(_09929_),
    .B(_10240_),
    .C(_09935_),
    .D(_10149_),
    .X(_09837_));
 sky130_fd_sc_hd__buf_1 _26918_ (.A(_09837_),
    .X(_09838_));
 sky130_fd_sc_hd__buf_1 _26919_ (.A(_09838_),
    .X(_09839_));
 sky130_fd_sc_hd__buf_1 _26920_ (.A(_09838_),
    .X(_09840_));
 sky130_fd_sc_hd__nand2_2 _26921_ (.A(_10245_),
    .B(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__o211a_2 _26922_ (.A1(\decode.regfile.registers_21[0] ),
    .A2(_09839_),
    .B1(_09841_),
    .C1(_09836_),
    .X(_02927_));
 sky130_fd_sc_hd__nand2_2 _26923_ (.A(_09450_),
    .B(_09840_),
    .Y(_09842_));
 sky130_fd_sc_hd__o211a_2 _26924_ (.A1(\decode.regfile.registers_21[1] ),
    .A2(_09839_),
    .B1(_09842_),
    .C1(_09836_),
    .X(_02928_));
 sky130_fd_sc_hd__nand2_2 _26925_ (.A(_09969_),
    .B(_09840_),
    .Y(_09843_));
 sky130_fd_sc_hd__o211a_2 _26926_ (.A1(\decode.regfile.registers_21[2] ),
    .A2(_09839_),
    .B1(_09843_),
    .C1(_09836_),
    .X(_02929_));
 sky130_fd_sc_hd__nand2_2 _26927_ (.A(_09974_),
    .B(_09840_),
    .Y(_09844_));
 sky130_fd_sc_hd__o211a_2 _26928_ (.A1(\decode.regfile.registers_21[3] ),
    .A2(_09839_),
    .B1(_09844_),
    .C1(_09836_),
    .X(_02930_));
 sky130_fd_sc_hd__nand2_2 _26929_ (.A(_09983_),
    .B(_09840_),
    .Y(_09845_));
 sky130_fd_sc_hd__o211a_2 _26930_ (.A1(\decode.regfile.registers_21[4] ),
    .A2(_09839_),
    .B1(_09845_),
    .C1(_09836_),
    .X(_02931_));
 sky130_fd_sc_hd__nand2_2 _26931_ (.A(_09992_),
    .B(_09840_),
    .Y(_09846_));
 sky130_fd_sc_hd__o211a_2 _26932_ (.A1(\decode.regfile.registers_21[5] ),
    .A2(_09839_),
    .B1(_09846_),
    .C1(_09836_),
    .X(_02932_));
 sky130_fd_sc_hd__nand2_2 _26933_ (.A(_09998_),
    .B(_09840_),
    .Y(_09847_));
 sky130_fd_sc_hd__o211a_2 _26934_ (.A1(\decode.regfile.registers_21[6] ),
    .A2(_09839_),
    .B1(_09847_),
    .C1(_09836_),
    .X(_02933_));
 sky130_fd_sc_hd__nand2_2 _26935_ (.A(_10007_),
    .B(_09840_),
    .Y(_09848_));
 sky130_fd_sc_hd__o211a_2 _26936_ (.A1(\decode.regfile.registers_21[7] ),
    .A2(_09839_),
    .B1(_09848_),
    .C1(_09836_),
    .X(_02934_));
 sky130_fd_sc_hd__buf_1 _26937_ (.A(_09838_),
    .X(_09849_));
 sky130_fd_sc_hd__nand2_2 _26938_ (.A(_10014_),
    .B(_09849_),
    .Y(_09850_));
 sky130_fd_sc_hd__o211a_2 _26939_ (.A1(\decode.regfile.registers_21[8] ),
    .A2(_09839_),
    .B1(_09850_),
    .C1(_09836_),
    .X(_02935_));
 sky130_fd_sc_hd__nand2_2 _26940_ (.A(_10024_),
    .B(_09849_),
    .Y(_09851_));
 sky130_fd_sc_hd__buf_1 _26941_ (.A(_09956_),
    .X(_09852_));
 sky130_fd_sc_hd__o211a_2 _26942_ (.A1(\decode.regfile.registers_21[9] ),
    .A2(_09839_),
    .B1(_09851_),
    .C1(_09852_),
    .X(_02936_));
 sky130_fd_sc_hd__buf_1 _26943_ (.A(_09838_),
    .X(_09853_));
 sky130_fd_sc_hd__nand2_2 _26944_ (.A(_10030_),
    .B(_09849_),
    .Y(_09854_));
 sky130_fd_sc_hd__o211a_2 _26945_ (.A1(\decode.regfile.registers_21[10] ),
    .A2(_09853_),
    .B1(_09854_),
    .C1(_09852_),
    .X(_02937_));
 sky130_fd_sc_hd__nand2_2 _26946_ (.A(_10035_),
    .B(_09849_),
    .Y(_09855_));
 sky130_fd_sc_hd__o211a_2 _26947_ (.A1(\decode.regfile.registers_21[11] ),
    .A2(_09853_),
    .B1(_09855_),
    .C1(_09852_),
    .X(_02938_));
 sky130_fd_sc_hd__nand2_2 _26948_ (.A(_10041_),
    .B(_09849_),
    .Y(_09856_));
 sky130_fd_sc_hd__o211a_2 _26949_ (.A1(\decode.regfile.registers_21[12] ),
    .A2(_09853_),
    .B1(_09856_),
    .C1(_09852_),
    .X(_02939_));
 sky130_fd_sc_hd__nand2_2 _26950_ (.A(_10047_),
    .B(_09849_),
    .Y(_09857_));
 sky130_fd_sc_hd__o211a_2 _26951_ (.A1(\decode.regfile.registers_21[13] ),
    .A2(_09853_),
    .B1(_09857_),
    .C1(_09852_),
    .X(_02940_));
 sky130_fd_sc_hd__nand2_2 _26952_ (.A(_10052_),
    .B(_09849_),
    .Y(_09858_));
 sky130_fd_sc_hd__o211a_2 _26953_ (.A1(\decode.regfile.registers_21[14] ),
    .A2(_09853_),
    .B1(_09858_),
    .C1(_09852_),
    .X(_02941_));
 sky130_fd_sc_hd__nand2_2 _26954_ (.A(_10057_),
    .B(_09849_),
    .Y(_09859_));
 sky130_fd_sc_hd__o211a_2 _26955_ (.A1(\decode.regfile.registers_21[15] ),
    .A2(_09853_),
    .B1(_09859_),
    .C1(_09852_),
    .X(_02942_));
 sky130_fd_sc_hd__nand2_2 _26956_ (.A(_10063_),
    .B(_09849_),
    .Y(_09860_));
 sky130_fd_sc_hd__o211a_2 _26957_ (.A1(\decode.regfile.registers_21[16] ),
    .A2(_09853_),
    .B1(_09860_),
    .C1(_09852_),
    .X(_02943_));
 sky130_fd_sc_hd__nand2_2 _26958_ (.A(_10068_),
    .B(_09849_),
    .Y(_09861_));
 sky130_fd_sc_hd__o211a_2 _26959_ (.A1(\decode.regfile.registers_21[17] ),
    .A2(_09853_),
    .B1(_09861_),
    .C1(_09852_),
    .X(_02944_));
 sky130_fd_sc_hd__buf_1 _26960_ (.A(_09838_),
    .X(_09862_));
 sky130_fd_sc_hd__nand2_2 _26961_ (.A(_10073_),
    .B(_09862_),
    .Y(_09863_));
 sky130_fd_sc_hd__o211a_2 _26962_ (.A1(\decode.regfile.registers_21[18] ),
    .A2(_09853_),
    .B1(_09863_),
    .C1(_09852_),
    .X(_02945_));
 sky130_fd_sc_hd__nand2_2 _26963_ (.A(_10080_),
    .B(_09862_),
    .Y(_09864_));
 sky130_fd_sc_hd__buf_1 _26964_ (.A(_09956_),
    .X(_09865_));
 sky130_fd_sc_hd__o211a_2 _26965_ (.A1(\decode.regfile.registers_21[19] ),
    .A2(_09853_),
    .B1(_09864_),
    .C1(_09865_),
    .X(_02946_));
 sky130_fd_sc_hd__buf_1 _26966_ (.A(_09838_),
    .X(_09866_));
 sky130_fd_sc_hd__nand2_2 _26967_ (.A(_10086_),
    .B(_09862_),
    .Y(_09867_));
 sky130_fd_sc_hd__o211a_2 _26968_ (.A1(\decode.regfile.registers_21[20] ),
    .A2(_09866_),
    .B1(_09867_),
    .C1(_09865_),
    .X(_02947_));
 sky130_fd_sc_hd__nand2_2 _26969_ (.A(_10091_),
    .B(_09862_),
    .Y(_09868_));
 sky130_fd_sc_hd__o211a_2 _26970_ (.A1(\decode.regfile.registers_21[21] ),
    .A2(_09866_),
    .B1(_09868_),
    .C1(_09865_),
    .X(_02948_));
 sky130_fd_sc_hd__nand2_2 _26971_ (.A(_10096_),
    .B(_09862_),
    .Y(_09869_));
 sky130_fd_sc_hd__o211a_2 _26972_ (.A1(\decode.regfile.registers_21[22] ),
    .A2(_09866_),
    .B1(_09869_),
    .C1(_09865_),
    .X(_02949_));
 sky130_fd_sc_hd__nand2_2 _26973_ (.A(_10101_),
    .B(_09862_),
    .Y(_09870_));
 sky130_fd_sc_hd__o211a_2 _26974_ (.A1(\decode.regfile.registers_21[23] ),
    .A2(_09866_),
    .B1(_09870_),
    .C1(_09865_),
    .X(_02950_));
 sky130_fd_sc_hd__nand2_2 _26975_ (.A(_10106_),
    .B(_09862_),
    .Y(_09871_));
 sky130_fd_sc_hd__o211a_2 _26976_ (.A1(\decode.regfile.registers_21[24] ),
    .A2(_09866_),
    .B1(_09871_),
    .C1(_09865_),
    .X(_02951_));
 sky130_fd_sc_hd__nand2_2 _26977_ (.A(_10111_),
    .B(_09862_),
    .Y(_09872_));
 sky130_fd_sc_hd__o211a_2 _26978_ (.A1(\decode.regfile.registers_21[25] ),
    .A2(_09866_),
    .B1(_09872_),
    .C1(_09865_),
    .X(_02952_));
 sky130_fd_sc_hd__nand2_2 _26979_ (.A(_10116_),
    .B(_09862_),
    .Y(_09873_));
 sky130_fd_sc_hd__o211a_2 _26980_ (.A1(\decode.regfile.registers_21[26] ),
    .A2(_09866_),
    .B1(_09873_),
    .C1(_09865_),
    .X(_02953_));
 sky130_fd_sc_hd__nand2_2 _26981_ (.A(_10121_),
    .B(_09862_),
    .Y(_09874_));
 sky130_fd_sc_hd__o211a_2 _26982_ (.A1(\decode.regfile.registers_21[27] ),
    .A2(_09866_),
    .B1(_09874_),
    .C1(_09865_),
    .X(_02954_));
 sky130_fd_sc_hd__nand2_2 _26983_ (.A(_10127_),
    .B(_09838_),
    .Y(_09875_));
 sky130_fd_sc_hd__o211a_2 _26984_ (.A1(\decode.regfile.registers_21[28] ),
    .A2(_09866_),
    .B1(_09875_),
    .C1(_09865_),
    .X(_02955_));
 sky130_fd_sc_hd__nand2_2 _26985_ (.A(_10135_),
    .B(_09838_),
    .Y(_09876_));
 sky130_fd_sc_hd__o211a_2 _26986_ (.A1(\decode.regfile.registers_21[29] ),
    .A2(_09866_),
    .B1(_09876_),
    .C1(_06396_),
    .X(_02956_));
 sky130_fd_sc_hd__nand2_2 _26987_ (.A(_10141_),
    .B(_09838_),
    .Y(_09877_));
 sky130_fd_sc_hd__o211a_2 _26988_ (.A1(\decode.regfile.registers_21[30] ),
    .A2(_09840_),
    .B1(_09877_),
    .C1(_06396_),
    .X(_02957_));
 sky130_fd_sc_hd__nand2_2 _26989_ (.A(_10146_),
    .B(_09838_),
    .Y(_09878_));
 sky130_fd_sc_hd__o211a_2 _26990_ (.A1(\decode.regfile.registers_21[31] ),
    .A2(_09840_),
    .B1(_09878_),
    .C1(_06396_),
    .X(_02958_));
 sky130_fd_sc_hd__dfxtp_2 _26991_ (.CLK(clock),
    .D(_00020_),
    .Q(\decode.regfile.registers_22[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26992_ (.CLK(clock),
    .D(_00021_),
    .Q(\decode.regfile.registers_22[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26993_ (.CLK(clock),
    .D(_00022_),
    .Q(\decode.regfile.registers_22[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26994_ (.CLK(clock),
    .D(_00023_),
    .Q(\decode.regfile.registers_22[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26995_ (.CLK(clock),
    .D(_00024_),
    .Q(\decode.regfile.registers_22[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26996_ (.CLK(clock),
    .D(_00025_),
    .Q(\decode.regfile.registers_22[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26997_ (.CLK(clock),
    .D(_00026_),
    .Q(\decode.regfile.registers_22[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26998_ (.CLK(clock),
    .D(_00027_),
    .Q(\decode.regfile.registers_22[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26999_ (.CLK(clock),
    .D(_00028_),
    .Q(\decode.regfile.registers_22[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27000_ (.CLK(clock),
    .D(_00029_),
    .Q(\decode.regfile.registers_22[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27001_ (.CLK(clock),
    .D(_00030_),
    .Q(\decode.regfile.registers_22[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27002_ (.CLK(clock),
    .D(_00031_),
    .Q(\decode.regfile.registers_22[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27003_ (.CLK(clock),
    .D(_00032_),
    .Q(\decode.regfile.registers_22[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27004_ (.CLK(clock),
    .D(_00033_),
    .Q(\decode.regfile.registers_22[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27005_ (.CLK(clock),
    .D(_00034_),
    .Q(\decode.regfile.registers_22[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27006_ (.CLK(clock),
    .D(_00035_),
    .Q(\decode.regfile.registers_22[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27007_ (.CLK(clock),
    .D(_00036_),
    .Q(\decode.regfile.registers_22[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27008_ (.CLK(clock),
    .D(_00037_),
    .Q(\decode.regfile.registers_22[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27009_ (.CLK(clock),
    .D(_00038_),
    .Q(\decode.regfile.registers_22[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27010_ (.CLK(clock),
    .D(_00039_),
    .Q(\decode.regfile.registers_22[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27011_ (.CLK(clock),
    .D(_00040_),
    .Q(\decode.regfile.registers_22[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27012_ (.CLK(clock),
    .D(_00041_),
    .Q(\decode.regfile.registers_22[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27013_ (.CLK(clock),
    .D(_00042_),
    .Q(\decode.regfile.registers_22[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27014_ (.CLK(clock),
    .D(_00043_),
    .Q(\decode.regfile.registers_22[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27015_ (.CLK(clock),
    .D(_00044_),
    .Q(\decode.regfile.registers_22[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27016_ (.CLK(clock),
    .D(_00045_),
    .Q(\decode.regfile.registers_22[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27017_ (.CLK(clock),
    .D(_00046_),
    .Q(\decode.regfile.registers_22[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27018_ (.CLK(clock),
    .D(_00047_),
    .Q(\decode.regfile.registers_22[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27019_ (.CLK(clock),
    .D(_00048_),
    .Q(\decode.regfile.registers_22[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27020_ (.CLK(clock),
    .D(_00049_),
    .Q(\decode.regfile.registers_22[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27021_ (.CLK(clock),
    .D(_00050_),
    .Q(\decode.regfile.registers_22[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27022_ (.CLK(clock),
    .D(_00051_),
    .Q(\decode.regfile.registers_22[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27023_ (.CLK(clock),
    .D(_00052_),
    .Q(\decode.regfile.registers_23[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27024_ (.CLK(clock),
    .D(_00053_),
    .Q(\decode.regfile.registers_23[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27025_ (.CLK(clock),
    .D(_00054_),
    .Q(\decode.regfile.registers_23[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27026_ (.CLK(clock),
    .D(_00055_),
    .Q(\decode.regfile.registers_23[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27027_ (.CLK(clock),
    .D(_00056_),
    .Q(\decode.regfile.registers_23[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27028_ (.CLK(clock),
    .D(_00057_),
    .Q(\decode.regfile.registers_23[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27029_ (.CLK(clock),
    .D(_00058_),
    .Q(\decode.regfile.registers_23[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27030_ (.CLK(clock),
    .D(_00059_),
    .Q(\decode.regfile.registers_23[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27031_ (.CLK(clock),
    .D(_00060_),
    .Q(\decode.regfile.registers_23[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27032_ (.CLK(clock),
    .D(_00061_),
    .Q(\decode.regfile.registers_23[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27033_ (.CLK(clock),
    .D(_00062_),
    .Q(\decode.regfile.registers_23[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27034_ (.CLK(clock),
    .D(_00063_),
    .Q(\decode.regfile.registers_23[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27035_ (.CLK(clock),
    .D(_00064_),
    .Q(\decode.regfile.registers_23[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27036_ (.CLK(clock),
    .D(_00065_),
    .Q(\decode.regfile.registers_23[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27037_ (.CLK(clock),
    .D(_00066_),
    .Q(\decode.regfile.registers_23[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27038_ (.CLK(clock),
    .D(_00067_),
    .Q(\decode.regfile.registers_23[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27039_ (.CLK(clock),
    .D(_00068_),
    .Q(\decode.regfile.registers_23[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27040_ (.CLK(clock),
    .D(_00069_),
    .Q(\decode.regfile.registers_23[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27041_ (.CLK(clock),
    .D(_00070_),
    .Q(\decode.regfile.registers_23[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27042_ (.CLK(clock),
    .D(_00071_),
    .Q(\decode.regfile.registers_23[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27043_ (.CLK(clock),
    .D(_00072_),
    .Q(\decode.regfile.registers_23[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27044_ (.CLK(clock),
    .D(_00073_),
    .Q(\decode.regfile.registers_23[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27045_ (.CLK(clock),
    .D(_00074_),
    .Q(\decode.regfile.registers_23[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27046_ (.CLK(clock),
    .D(_00075_),
    .Q(\decode.regfile.registers_23[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27047_ (.CLK(clock),
    .D(_00076_),
    .Q(\decode.regfile.registers_23[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27048_ (.CLK(clock),
    .D(_00077_),
    .Q(\decode.regfile.registers_23[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27049_ (.CLK(clock),
    .D(_00078_),
    .Q(\decode.regfile.registers_23[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27050_ (.CLK(clock),
    .D(_00079_),
    .Q(\decode.regfile.registers_23[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27051_ (.CLK(clock),
    .D(_00080_),
    .Q(\decode.regfile.registers_23[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27052_ (.CLK(clock),
    .D(_00081_),
    .Q(\decode.regfile.registers_23[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27053_ (.CLK(clock),
    .D(_00082_),
    .Q(\decode.regfile.registers_23[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27054_ (.CLK(clock),
    .D(_00083_),
    .Q(\decode.regfile.registers_23[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27055_ (.CLK(clock),
    .D(_00084_),
    .Q(\decode.regfile.registers_24[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27056_ (.CLK(clock),
    .D(_00085_),
    .Q(\decode.regfile.registers_24[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27057_ (.CLK(clock),
    .D(_00086_),
    .Q(\decode.regfile.registers_24[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27058_ (.CLK(clock),
    .D(_00087_),
    .Q(\decode.regfile.registers_24[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27059_ (.CLK(clock),
    .D(_00088_),
    .Q(\decode.regfile.registers_24[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27060_ (.CLK(clock),
    .D(_00089_),
    .Q(\decode.regfile.registers_24[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27061_ (.CLK(clock),
    .D(_00090_),
    .Q(\decode.regfile.registers_24[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27062_ (.CLK(clock),
    .D(_00091_),
    .Q(\decode.regfile.registers_24[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27063_ (.CLK(clock),
    .D(_00092_),
    .Q(\decode.regfile.registers_24[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27064_ (.CLK(clock),
    .D(_00093_),
    .Q(\decode.regfile.registers_24[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27065_ (.CLK(clock),
    .D(_00094_),
    .Q(\decode.regfile.registers_24[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27066_ (.CLK(clock),
    .D(_00095_),
    .Q(\decode.regfile.registers_24[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27067_ (.CLK(clock),
    .D(_00096_),
    .Q(\decode.regfile.registers_24[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27068_ (.CLK(clock),
    .D(_00097_),
    .Q(\decode.regfile.registers_24[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27069_ (.CLK(clock),
    .D(_00098_),
    .Q(\decode.regfile.registers_24[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27070_ (.CLK(clock),
    .D(_00099_),
    .Q(\decode.regfile.registers_24[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27071_ (.CLK(clock),
    .D(_00100_),
    .Q(\decode.regfile.registers_24[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27072_ (.CLK(clock),
    .D(_00101_),
    .Q(\decode.regfile.registers_24[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27073_ (.CLK(clock),
    .D(_00102_),
    .Q(\decode.regfile.registers_24[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27074_ (.CLK(clock),
    .D(_00103_),
    .Q(\decode.regfile.registers_24[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27075_ (.CLK(clock),
    .D(_00104_),
    .Q(\decode.regfile.registers_24[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27076_ (.CLK(clock),
    .D(_00105_),
    .Q(\decode.regfile.registers_24[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27077_ (.CLK(clock),
    .D(_00106_),
    .Q(\decode.regfile.registers_24[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27078_ (.CLK(clock),
    .D(_00107_),
    .Q(\decode.regfile.registers_24[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27079_ (.CLK(clock),
    .D(_00108_),
    .Q(\decode.regfile.registers_24[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27080_ (.CLK(clock),
    .D(_00109_),
    .Q(\decode.regfile.registers_24[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27081_ (.CLK(clock),
    .D(_00110_),
    .Q(\decode.regfile.registers_24[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27082_ (.CLK(clock),
    .D(_00111_),
    .Q(\decode.regfile.registers_24[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27083_ (.CLK(clock),
    .D(_00112_),
    .Q(\decode.regfile.registers_24[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27084_ (.CLK(clock),
    .D(_00113_),
    .Q(\decode.regfile.registers_24[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27085_ (.CLK(clock),
    .D(_00114_),
    .Q(\decode.regfile.registers_24[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27086_ (.CLK(clock),
    .D(_00115_),
    .Q(\decode.regfile.registers_24[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27087_ (.CLK(clock),
    .D(_00116_),
    .Q(\decode.regfile.registers_25[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27088_ (.CLK(clock),
    .D(_00117_),
    .Q(\decode.regfile.registers_25[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27089_ (.CLK(clock),
    .D(_00118_),
    .Q(\decode.regfile.registers_25[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27090_ (.CLK(clock),
    .D(_00119_),
    .Q(\decode.regfile.registers_25[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27091_ (.CLK(clock),
    .D(_00120_),
    .Q(\decode.regfile.registers_25[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27092_ (.CLK(clock),
    .D(_00121_),
    .Q(\decode.regfile.registers_25[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27093_ (.CLK(clock),
    .D(_00122_),
    .Q(\decode.regfile.registers_25[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27094_ (.CLK(clock),
    .D(_00123_),
    .Q(\decode.regfile.registers_25[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27095_ (.CLK(clock),
    .D(_00124_),
    .Q(\decode.regfile.registers_25[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27096_ (.CLK(clock),
    .D(_00125_),
    .Q(\decode.regfile.registers_25[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27097_ (.CLK(clock),
    .D(_00126_),
    .Q(\decode.regfile.registers_25[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27098_ (.CLK(clock),
    .D(_00127_),
    .Q(\decode.regfile.registers_25[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27099_ (.CLK(clock),
    .D(_00128_),
    .Q(\decode.regfile.registers_25[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27100_ (.CLK(clock),
    .D(_00129_),
    .Q(\decode.regfile.registers_25[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27101_ (.CLK(clock),
    .D(_00130_),
    .Q(\decode.regfile.registers_25[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27102_ (.CLK(clock),
    .D(_00131_),
    .Q(\decode.regfile.registers_25[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27103_ (.CLK(clock),
    .D(_00132_),
    .Q(\decode.regfile.registers_25[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27104_ (.CLK(clock),
    .D(_00133_),
    .Q(\decode.regfile.registers_25[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27105_ (.CLK(clock),
    .D(_00134_),
    .Q(\decode.regfile.registers_25[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27106_ (.CLK(clock),
    .D(_00135_),
    .Q(\decode.regfile.registers_25[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27107_ (.CLK(clock),
    .D(_00136_),
    .Q(\decode.regfile.registers_25[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27108_ (.CLK(clock),
    .D(_00137_),
    .Q(\decode.regfile.registers_25[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27109_ (.CLK(clock),
    .D(_00138_),
    .Q(\decode.regfile.registers_25[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27110_ (.CLK(clock),
    .D(_00139_),
    .Q(\decode.regfile.registers_25[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27111_ (.CLK(clock),
    .D(_00140_),
    .Q(\decode.regfile.registers_25[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27112_ (.CLK(clock),
    .D(_00141_),
    .Q(\decode.regfile.registers_25[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27113_ (.CLK(clock),
    .D(_00142_),
    .Q(\decode.regfile.registers_25[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27114_ (.CLK(clock),
    .D(_00143_),
    .Q(\decode.regfile.registers_25[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27115_ (.CLK(clock),
    .D(_00144_),
    .Q(\decode.regfile.registers_25[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27116_ (.CLK(clock),
    .D(_00145_),
    .Q(\decode.regfile.registers_25[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27117_ (.CLK(clock),
    .D(_00146_),
    .Q(\decode.regfile.registers_25[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27118_ (.CLK(clock),
    .D(_00147_),
    .Q(\decode.regfile.registers_25[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27119_ (.CLK(clock),
    .D(_00148_),
    .Q(\decode.regfile.registers_26[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27120_ (.CLK(clock),
    .D(_00149_),
    .Q(\decode.regfile.registers_26[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27121_ (.CLK(clock),
    .D(_00150_),
    .Q(\decode.regfile.registers_26[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27122_ (.CLK(clock),
    .D(_00151_),
    .Q(\decode.regfile.registers_26[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27123_ (.CLK(clock),
    .D(_00152_),
    .Q(\decode.regfile.registers_26[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27124_ (.CLK(clock),
    .D(_00153_),
    .Q(\decode.regfile.registers_26[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27125_ (.CLK(clock),
    .D(_00154_),
    .Q(\decode.regfile.registers_26[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27126_ (.CLK(clock),
    .D(_00155_),
    .Q(\decode.regfile.registers_26[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27127_ (.CLK(clock),
    .D(_00156_),
    .Q(\decode.regfile.registers_26[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27128_ (.CLK(clock),
    .D(_00157_),
    .Q(\decode.regfile.registers_26[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27129_ (.CLK(clock),
    .D(_00158_),
    .Q(\decode.regfile.registers_26[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27130_ (.CLK(clock),
    .D(_00159_),
    .Q(\decode.regfile.registers_26[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27131_ (.CLK(clock),
    .D(_00160_),
    .Q(\decode.regfile.registers_26[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27132_ (.CLK(clock),
    .D(_00161_),
    .Q(\decode.regfile.registers_26[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27133_ (.CLK(clock),
    .D(_00162_),
    .Q(\decode.regfile.registers_26[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27134_ (.CLK(clock),
    .D(_00163_),
    .Q(\decode.regfile.registers_26[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27135_ (.CLK(clock),
    .D(_00164_),
    .Q(\decode.regfile.registers_26[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27136_ (.CLK(clock),
    .D(_00165_),
    .Q(\decode.regfile.registers_26[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27137_ (.CLK(clock),
    .D(_00166_),
    .Q(\decode.regfile.registers_26[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27138_ (.CLK(clock),
    .D(_00167_),
    .Q(\decode.regfile.registers_26[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27139_ (.CLK(clock),
    .D(_00168_),
    .Q(\decode.regfile.registers_26[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27140_ (.CLK(clock),
    .D(_00169_),
    .Q(\decode.regfile.registers_26[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27141_ (.CLK(clock),
    .D(_00170_),
    .Q(\decode.regfile.registers_26[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27142_ (.CLK(clock),
    .D(_00171_),
    .Q(\decode.regfile.registers_26[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27143_ (.CLK(clock),
    .D(_00172_),
    .Q(\decode.regfile.registers_26[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27144_ (.CLK(clock),
    .D(_00173_),
    .Q(\decode.regfile.registers_26[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27145_ (.CLK(clock),
    .D(_00174_),
    .Q(\decode.regfile.registers_26[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27146_ (.CLK(clock),
    .D(_00175_),
    .Q(\decode.regfile.registers_26[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27147_ (.CLK(clock),
    .D(_00176_),
    .Q(\decode.regfile.registers_26[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27148_ (.CLK(clock),
    .D(_00177_),
    .Q(\decode.regfile.registers_26[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27149_ (.CLK(clock),
    .D(_00178_),
    .Q(\decode.regfile.registers_26[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27150_ (.CLK(clock),
    .D(_00179_),
    .Q(\decode.regfile.registers_26[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27151_ (.CLK(clock),
    .D(_00180_),
    .Q(\decode.regfile.registers_27[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27152_ (.CLK(clock),
    .D(_00181_),
    .Q(\decode.regfile.registers_27[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27153_ (.CLK(clock),
    .D(_00182_),
    .Q(\decode.regfile.registers_27[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27154_ (.CLK(clock),
    .D(_00183_),
    .Q(\decode.regfile.registers_27[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27155_ (.CLK(clock),
    .D(_00184_),
    .Q(\decode.regfile.registers_27[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27156_ (.CLK(clock),
    .D(_00185_),
    .Q(\decode.regfile.registers_27[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27157_ (.CLK(clock),
    .D(_00186_),
    .Q(\decode.regfile.registers_27[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27158_ (.CLK(clock),
    .D(_00187_),
    .Q(\decode.regfile.registers_27[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27159_ (.CLK(clock),
    .D(_00188_),
    .Q(\decode.regfile.registers_27[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27160_ (.CLK(clock),
    .D(_00189_),
    .Q(\decode.regfile.registers_27[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27161_ (.CLK(clock),
    .D(_00190_),
    .Q(\decode.regfile.registers_27[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27162_ (.CLK(clock),
    .D(_00191_),
    .Q(\decode.regfile.registers_27[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27163_ (.CLK(clock),
    .D(_00192_),
    .Q(\decode.regfile.registers_27[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27164_ (.CLK(clock),
    .D(_00193_),
    .Q(\decode.regfile.registers_27[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27165_ (.CLK(clock),
    .D(_00194_),
    .Q(\decode.regfile.registers_27[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27166_ (.CLK(clock),
    .D(_00195_),
    .Q(\decode.regfile.registers_27[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27167_ (.CLK(clock),
    .D(_00196_),
    .Q(\decode.regfile.registers_27[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27168_ (.CLK(clock),
    .D(_00197_),
    .Q(\decode.regfile.registers_27[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27169_ (.CLK(clock),
    .D(_00198_),
    .Q(\decode.regfile.registers_27[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27170_ (.CLK(clock),
    .D(_00199_),
    .Q(\decode.regfile.registers_27[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27171_ (.CLK(clock),
    .D(_00200_),
    .Q(\decode.regfile.registers_27[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27172_ (.CLK(clock),
    .D(_00201_),
    .Q(\decode.regfile.registers_27[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27173_ (.CLK(clock),
    .D(_00202_),
    .Q(\decode.regfile.registers_27[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27174_ (.CLK(clock),
    .D(_00203_),
    .Q(\decode.regfile.registers_27[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27175_ (.CLK(clock),
    .D(_00204_),
    .Q(\decode.regfile.registers_27[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27176_ (.CLK(clock),
    .D(_00205_),
    .Q(\decode.regfile.registers_27[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27177_ (.CLK(clock),
    .D(_00206_),
    .Q(\decode.regfile.registers_27[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27178_ (.CLK(clock),
    .D(_00207_),
    .Q(\decode.regfile.registers_27[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27179_ (.CLK(clock),
    .D(_00208_),
    .Q(\decode.regfile.registers_27[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27180_ (.CLK(clock),
    .D(_00209_),
    .Q(\decode.regfile.registers_27[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27181_ (.CLK(clock),
    .D(_00210_),
    .Q(\decode.regfile.registers_27[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27182_ (.CLK(clock),
    .D(_00211_),
    .Q(\decode.regfile.registers_27[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27183_ (.CLK(clock),
    .D(_00212_),
    .Q(\decode.regfile.registers_28[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27184_ (.CLK(clock),
    .D(_00213_),
    .Q(\decode.regfile.registers_28[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27185_ (.CLK(clock),
    .D(_00214_),
    .Q(\decode.regfile.registers_28[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27186_ (.CLK(clock),
    .D(_00215_),
    .Q(\decode.regfile.registers_28[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27187_ (.CLK(clock),
    .D(_00216_),
    .Q(\decode.regfile.registers_28[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27188_ (.CLK(clock),
    .D(_00217_),
    .Q(\decode.regfile.registers_28[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27189_ (.CLK(clock),
    .D(_00218_),
    .Q(\decode.regfile.registers_28[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27190_ (.CLK(clock),
    .D(_00219_),
    .Q(\decode.regfile.registers_28[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27191_ (.CLK(clock),
    .D(_00220_),
    .Q(\decode.regfile.registers_28[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27192_ (.CLK(clock),
    .D(_00221_),
    .Q(\decode.regfile.registers_28[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27193_ (.CLK(clock),
    .D(_00222_),
    .Q(\decode.regfile.registers_28[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27194_ (.CLK(clock),
    .D(_00223_),
    .Q(\decode.regfile.registers_28[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27195_ (.CLK(clock),
    .D(_00224_),
    .Q(\decode.regfile.registers_28[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27196_ (.CLK(clock),
    .D(_00225_),
    .Q(\decode.regfile.registers_28[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27197_ (.CLK(clock),
    .D(_00226_),
    .Q(\decode.regfile.registers_28[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27198_ (.CLK(clock),
    .D(_00227_),
    .Q(\decode.regfile.registers_28[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27199_ (.CLK(clock),
    .D(_00228_),
    .Q(\decode.regfile.registers_28[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27200_ (.CLK(clock),
    .D(_00229_),
    .Q(\decode.regfile.registers_28[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27201_ (.CLK(clock),
    .D(_00230_),
    .Q(\decode.regfile.registers_28[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27202_ (.CLK(clock),
    .D(_00231_),
    .Q(\decode.regfile.registers_28[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27203_ (.CLK(clock),
    .D(_00232_),
    .Q(\decode.regfile.registers_28[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27204_ (.CLK(clock),
    .D(_00233_),
    .Q(\decode.regfile.registers_28[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27205_ (.CLK(clock),
    .D(_00234_),
    .Q(\decode.regfile.registers_28[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27206_ (.CLK(clock),
    .D(_00235_),
    .Q(\decode.regfile.registers_28[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27207_ (.CLK(clock),
    .D(_00236_),
    .Q(\decode.regfile.registers_28[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27208_ (.CLK(clock),
    .D(_00237_),
    .Q(\decode.regfile.registers_28[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27209_ (.CLK(clock),
    .D(_00238_),
    .Q(\decode.regfile.registers_28[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27210_ (.CLK(clock),
    .D(_00239_),
    .Q(\decode.regfile.registers_28[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27211_ (.CLK(clock),
    .D(_00240_),
    .Q(\decode.regfile.registers_28[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27212_ (.CLK(clock),
    .D(_00241_),
    .Q(\decode.regfile.registers_28[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27213_ (.CLK(clock),
    .D(_00242_),
    .Q(\decode.regfile.registers_28[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27214_ (.CLK(clock),
    .D(_00243_),
    .Q(\decode.regfile.registers_28[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27215_ (.CLK(clock),
    .D(_00244_),
    .Q(\decode.regfile.registers_29[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27216_ (.CLK(clock),
    .D(_00245_),
    .Q(\decode.regfile.registers_29[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27217_ (.CLK(clock),
    .D(_00246_),
    .Q(\decode.regfile.registers_29[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27218_ (.CLK(clock),
    .D(_00247_),
    .Q(\decode.regfile.registers_29[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27219_ (.CLK(clock),
    .D(_00248_),
    .Q(\decode.regfile.registers_29[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27220_ (.CLK(clock),
    .D(_00249_),
    .Q(\decode.regfile.registers_29[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27221_ (.CLK(clock),
    .D(_00250_),
    .Q(\decode.regfile.registers_29[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27222_ (.CLK(clock),
    .D(_00251_),
    .Q(\decode.regfile.registers_29[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27223_ (.CLK(clock),
    .D(_00252_),
    .Q(\decode.regfile.registers_29[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27224_ (.CLK(clock),
    .D(_00253_),
    .Q(\decode.regfile.registers_29[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27225_ (.CLK(clock),
    .D(_00254_),
    .Q(\decode.regfile.registers_29[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27226_ (.CLK(clock),
    .D(_00255_),
    .Q(\decode.regfile.registers_29[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27227_ (.CLK(clock),
    .D(_00256_),
    .Q(\decode.regfile.registers_29[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27228_ (.CLK(clock),
    .D(_00257_),
    .Q(\decode.regfile.registers_29[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27229_ (.CLK(clock),
    .D(_00258_),
    .Q(\decode.regfile.registers_29[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27230_ (.CLK(clock),
    .D(_00259_),
    .Q(\decode.regfile.registers_29[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27231_ (.CLK(clock),
    .D(_00260_),
    .Q(\decode.regfile.registers_29[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27232_ (.CLK(clock),
    .D(_00261_),
    .Q(\decode.regfile.registers_29[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27233_ (.CLK(clock),
    .D(_00262_),
    .Q(\decode.regfile.registers_29[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27234_ (.CLK(clock),
    .D(_00263_),
    .Q(\decode.regfile.registers_29[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27235_ (.CLK(clock),
    .D(_00264_),
    .Q(\decode.regfile.registers_29[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27236_ (.CLK(clock),
    .D(_00265_),
    .Q(\decode.regfile.registers_29[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27237_ (.CLK(clock),
    .D(_00266_),
    .Q(\decode.regfile.registers_29[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27238_ (.CLK(clock),
    .D(_00267_),
    .Q(\decode.regfile.registers_29[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27239_ (.CLK(clock),
    .D(_00268_),
    .Q(\decode.regfile.registers_29[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27240_ (.CLK(clock),
    .D(_00269_),
    .Q(\decode.regfile.registers_29[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27241_ (.CLK(clock),
    .D(_00270_),
    .Q(\decode.regfile.registers_29[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27242_ (.CLK(clock),
    .D(_00271_),
    .Q(\decode.regfile.registers_29[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27243_ (.CLK(clock),
    .D(_00272_),
    .Q(\decode.regfile.registers_29[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27244_ (.CLK(clock),
    .D(_00273_),
    .Q(\decode.regfile.registers_29[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27245_ (.CLK(clock),
    .D(_00274_),
    .Q(\decode.regfile.registers_29[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27246_ (.CLK(clock),
    .D(_00275_),
    .Q(\decode.regfile.registers_29[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27247_ (.CLK(clock),
    .D(_00276_),
    .Q(\decode.regfile.registers_30[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27248_ (.CLK(clock),
    .D(_00277_),
    .Q(\decode.regfile.registers_30[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27249_ (.CLK(clock),
    .D(_00278_),
    .Q(\decode.regfile.registers_30[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27250_ (.CLK(clock),
    .D(_00279_),
    .Q(\decode.regfile.registers_30[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27251_ (.CLK(clock),
    .D(_00280_),
    .Q(\decode.regfile.registers_30[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27252_ (.CLK(clock),
    .D(_00281_),
    .Q(\decode.regfile.registers_30[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27253_ (.CLK(clock),
    .D(_00282_),
    .Q(\decode.regfile.registers_30[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27254_ (.CLK(clock),
    .D(_00283_),
    .Q(\decode.regfile.registers_30[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27255_ (.CLK(clock),
    .D(_00284_),
    .Q(\decode.regfile.registers_30[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27256_ (.CLK(clock),
    .D(_00285_),
    .Q(\decode.regfile.registers_30[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27257_ (.CLK(clock),
    .D(_00286_),
    .Q(\decode.regfile.registers_30[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27258_ (.CLK(clock),
    .D(_00287_),
    .Q(\decode.regfile.registers_30[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27259_ (.CLK(clock),
    .D(_00288_),
    .Q(\decode.regfile.registers_30[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27260_ (.CLK(clock),
    .D(_00289_),
    .Q(\decode.regfile.registers_30[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27261_ (.CLK(clock),
    .D(_00290_),
    .Q(\decode.regfile.registers_30[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27262_ (.CLK(clock),
    .D(_00291_),
    .Q(\decode.regfile.registers_30[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27263_ (.CLK(clock),
    .D(_00292_),
    .Q(\decode.regfile.registers_30[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27264_ (.CLK(clock),
    .D(_00293_),
    .Q(\decode.regfile.registers_30[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27265_ (.CLK(clock),
    .D(_00294_),
    .Q(\decode.regfile.registers_30[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27266_ (.CLK(clock),
    .D(_00295_),
    .Q(\decode.regfile.registers_30[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27267_ (.CLK(clock),
    .D(_00296_),
    .Q(\decode.regfile.registers_30[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27268_ (.CLK(clock),
    .D(_00297_),
    .Q(\decode.regfile.registers_30[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27269_ (.CLK(clock),
    .D(_00298_),
    .Q(\decode.regfile.registers_30[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27270_ (.CLK(clock),
    .D(_00299_),
    .Q(\decode.regfile.registers_30[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27271_ (.CLK(clock),
    .D(_00300_),
    .Q(\decode.regfile.registers_30[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27272_ (.CLK(clock),
    .D(_00301_),
    .Q(\decode.regfile.registers_30[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27273_ (.CLK(clock),
    .D(_00302_),
    .Q(\decode.regfile.registers_30[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27274_ (.CLK(clock),
    .D(_00303_),
    .Q(\decode.regfile.registers_30[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27275_ (.CLK(clock),
    .D(_00304_),
    .Q(\decode.regfile.registers_30[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27276_ (.CLK(clock),
    .D(_00305_),
    .Q(\decode.regfile.registers_30[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27277_ (.CLK(clock),
    .D(_00306_),
    .Q(\decode.regfile.registers_30[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27278_ (.CLK(clock),
    .D(_00307_),
    .Q(\decode.regfile.registers_30[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27279_ (.CLK(clock),
    .D(_00308_),
    .Q(\decode.regfile.registers_31[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27280_ (.CLK(clock),
    .D(_00309_),
    .Q(\decode.regfile.registers_31[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27281_ (.CLK(clock),
    .D(_00310_),
    .Q(\decode.regfile.registers_31[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27282_ (.CLK(clock),
    .D(_00311_),
    .Q(\decode.regfile.registers_31[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27283_ (.CLK(clock),
    .D(_00312_),
    .Q(\decode.regfile.registers_31[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27284_ (.CLK(clock),
    .D(_00313_),
    .Q(\decode.regfile.registers_31[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27285_ (.CLK(clock),
    .D(_00314_),
    .Q(\decode.regfile.registers_31[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27286_ (.CLK(clock),
    .D(_00315_),
    .Q(\decode.regfile.registers_31[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27287_ (.CLK(clock),
    .D(_00316_),
    .Q(\decode.regfile.registers_31[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27288_ (.CLK(clock),
    .D(_00317_),
    .Q(\decode.regfile.registers_31[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27289_ (.CLK(clock),
    .D(_00318_),
    .Q(\decode.regfile.registers_31[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27290_ (.CLK(clock),
    .D(_00319_),
    .Q(\decode.regfile.registers_31[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27291_ (.CLK(clock),
    .D(_00320_),
    .Q(\decode.regfile.registers_31[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27292_ (.CLK(clock),
    .D(_00321_),
    .Q(\decode.regfile.registers_31[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27293_ (.CLK(clock),
    .D(_00322_),
    .Q(\decode.regfile.registers_31[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27294_ (.CLK(clock),
    .D(_00323_),
    .Q(\decode.regfile.registers_31[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27295_ (.CLK(clock),
    .D(_00324_),
    .Q(\decode.regfile.registers_31[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27296_ (.CLK(clock),
    .D(_00325_),
    .Q(\decode.regfile.registers_31[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27297_ (.CLK(clock),
    .D(_00326_),
    .Q(\decode.regfile.registers_31[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27298_ (.CLK(clock),
    .D(_00327_),
    .Q(\decode.regfile.registers_31[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27299_ (.CLK(clock),
    .D(_00328_),
    .Q(\decode.regfile.registers_31[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27300_ (.CLK(clock),
    .D(_00329_),
    .Q(\decode.regfile.registers_31[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27301_ (.CLK(clock),
    .D(_00330_),
    .Q(\decode.regfile.registers_31[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27302_ (.CLK(clock),
    .D(_00331_),
    .Q(\decode.regfile.registers_31[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27303_ (.CLK(clock),
    .D(_00332_),
    .Q(\decode.regfile.registers_31[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27304_ (.CLK(clock),
    .D(_00333_),
    .Q(\decode.regfile.registers_31[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27305_ (.CLK(clock),
    .D(_00334_),
    .Q(\decode.regfile.registers_31[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27306_ (.CLK(clock),
    .D(_00335_),
    .Q(\decode.regfile.registers_31[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27307_ (.CLK(clock),
    .D(_00336_),
    .Q(\decode.regfile.registers_31[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27308_ (.CLK(clock),
    .D(_00337_),
    .Q(\decode.regfile.registers_31[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27309_ (.CLK(clock),
    .D(_00338_),
    .Q(\decode.regfile.registers_31[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27310_ (.CLK(clock),
    .D(_00339_),
    .Q(\decode.regfile.registers_31[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27311_ (.CLK(clock),
    .D(_00340_),
    .Q(\fetch.btb.btbTable[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27312_ (.CLK(clock),
    .D(_00341_),
    .Q(\fetch.btb.btbTable[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27313_ (.CLK(clock),
    .D(_00342_),
    .Q(\decode.id_ex_ex_use_rs1_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27314_ (.CLK(clock),
    .D(_00343_),
    .Q(\decode.id_ex_ex_rd_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27315_ (.CLK(clock),
    .D(_00344_),
    .Q(\decode.id_ex_ex_rd_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27316_ (.CLK(clock),
    .D(_00345_),
    .Q(\decode.id_ex_ex_rd_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27317_ (.CLK(clock),
    .D(_00346_),
    .Q(\decode.id_ex_ex_rd_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27318_ (.CLK(clock),
    .D(_00347_),
    .Q(\decode.id_ex_ex_rd_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27319_ (.CLK(clock),
    .D(_00348_),
    .Q(\decode.id_ex_ex_rs1_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27320_ (.CLK(clock),
    .D(_00349_),
    .Q(\decode.id_ex_ex_rs1_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27321_ (.CLK(clock),
    .D(_00350_),
    .Q(\decode.id_ex_ex_rs1_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27322_ (.CLK(clock),
    .D(_00351_),
    .Q(\decode.id_ex_ex_rs1_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27323_ (.CLK(clock),
    .D(_00352_),
    .Q(\decode.id_ex_ex_rs1_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27324_ (.CLK(clock),
    .D(_00353_),
    .Q(\decode.id_ex_funct3_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27325_ (.CLK(clock),
    .D(_00354_),
    .Q(\decode.id_ex_funct3_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27326_ (.CLK(clock),
    .D(_00355_),
    .Q(\decode.id_ex_funct3_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27327_ (.CLK(clock),
    .D(_00356_),
    .Q(\decode.id_ex_imm_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27328_ (.CLK(clock),
    .D(_00357_),
    .Q(\decode.id_ex_imm_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27329_ (.CLK(clock),
    .D(_00358_),
    .Q(\decode.id_ex_imm_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27330_ (.CLK(clock),
    .D(_00359_),
    .Q(\decode.id_ex_imm_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27331_ (.CLK(clock),
    .D(_00360_),
    .Q(\decode.id_ex_imm_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27332_ (.CLK(clock),
    .D(_00361_),
    .Q(\decode.id_ex_imm_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27333_ (.CLK(clock),
    .D(_00362_),
    .Q(\decode.id_ex_imm_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27334_ (.CLK(clock),
    .D(_00363_),
    .Q(\decode.id_ex_imm_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27335_ (.CLK(clock),
    .D(_00364_),
    .Q(\decode.id_ex_imm_reg[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27336_ (.CLK(clock),
    .D(_00365_),
    .Q(\decode.id_ex_imm_reg[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27337_ (.CLK(clock),
    .D(_00366_),
    .Q(\decode.id_ex_imm_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27338_ (.CLK(clock),
    .D(_00367_),
    .Q(\decode.id_ex_imm_reg[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27339_ (.CLK(clock),
    .D(_00368_),
    .Q(\decode.id_ex_imm_reg[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27340_ (.CLK(clock),
    .D(_00369_),
    .Q(\decode.id_ex_imm_reg[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27341_ (.CLK(clock),
    .D(_00370_),
    .Q(\decode.id_ex_imm_reg[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27342_ (.CLK(clock),
    .D(_00371_),
    .Q(\decode.id_ex_imm_reg[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27343_ (.CLK(clock),
    .D(_00372_),
    .Q(\decode.id_ex_imm_reg[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27344_ (.CLK(clock),
    .D(_00373_),
    .Q(\decode.id_ex_imm_reg[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27345_ (.CLK(clock),
    .D(_00374_),
    .Q(\decode.id_ex_imm_reg[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27346_ (.CLK(clock),
    .D(_00375_),
    .Q(\decode.id_ex_imm_reg[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27347_ (.CLK(clock),
    .D(_00376_),
    .Q(\decode.id_ex_imm_reg[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27348_ (.CLK(clock),
    .D(_00377_),
    .Q(\decode.id_ex_imm_reg[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27349_ (.CLK(clock),
    .D(_00378_),
    .Q(\decode.id_ex_imm_reg[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27350_ (.CLK(clock),
    .D(_00379_),
    .Q(\decode.id_ex_imm_reg[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27351_ (.CLK(clock),
    .D(_00380_),
    .Q(\decode.id_ex_imm_reg[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27352_ (.CLK(clock),
    .D(_00381_),
    .Q(\decode.id_ex_imm_reg[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27353_ (.CLK(clock),
    .D(_00382_),
    .Q(\decode.id_ex_imm_reg[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27354_ (.CLK(clock),
    .D(_00383_),
    .Q(\decode.id_ex_imm_reg[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27355_ (.CLK(clock),
    .D(_00384_),
    .Q(\decode.id_ex_imm_reg[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27356_ (.CLK(clock),
    .D(_00385_),
    .Q(\decode.id_ex_imm_reg[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27357_ (.CLK(clock),
    .D(_00386_),
    .Q(\decode.id_ex_imm_reg[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27358_ (.CLK(clock),
    .D(_00387_),
    .Q(\decode.id_ex_imm_reg[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27359_ (.CLK(clock),
    .D(_00388_),
    .Q(\decode.id_ex_rs2_data_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27360_ (.CLK(clock),
    .D(_00389_),
    .Q(\decode.id_ex_rs2_data_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27361_ (.CLK(clock),
    .D(_00390_),
    .Q(\decode.id_ex_rs2_data_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27362_ (.CLK(clock),
    .D(_00391_),
    .Q(\decode.id_ex_rs2_data_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27363_ (.CLK(clock),
    .D(_00392_),
    .Q(\decode.id_ex_rs2_data_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27364_ (.CLK(clock),
    .D(_00393_),
    .Q(\decode.id_ex_rs2_data_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27365_ (.CLK(clock),
    .D(_00394_),
    .Q(\decode.id_ex_rs2_data_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27366_ (.CLK(clock),
    .D(_00395_),
    .Q(\decode.id_ex_rs2_data_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27367_ (.CLK(clock),
    .D(_00396_),
    .Q(\decode.id_ex_rs2_data_reg[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27368_ (.CLK(clock),
    .D(_00397_),
    .Q(\decode.id_ex_rs2_data_reg[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27369_ (.CLK(clock),
    .D(_00398_),
    .Q(\decode.id_ex_rs2_data_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27370_ (.CLK(clock),
    .D(_00399_),
    .Q(\decode.id_ex_rs2_data_reg[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27371_ (.CLK(clock),
    .D(_00400_),
    .Q(\decode.id_ex_rs2_data_reg[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27372_ (.CLK(clock),
    .D(_00401_),
    .Q(\decode.id_ex_rs2_data_reg[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27373_ (.CLK(clock),
    .D(_00402_),
    .Q(\decode.id_ex_rs2_data_reg[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27374_ (.CLK(clock),
    .D(_00403_),
    .Q(\decode.id_ex_rs2_data_reg[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27375_ (.CLK(clock),
    .D(_00404_),
    .Q(\decode.id_ex_rs2_data_reg[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27376_ (.CLK(clock),
    .D(_00405_),
    .Q(\decode.id_ex_rs2_data_reg[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27377_ (.CLK(clock),
    .D(_00406_),
    .Q(\decode.id_ex_rs2_data_reg[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27378_ (.CLK(clock),
    .D(_00407_),
    .Q(\decode.id_ex_rs2_data_reg[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27379_ (.CLK(clock),
    .D(_00408_),
    .Q(\decode.id_ex_rs2_data_reg[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27380_ (.CLK(clock),
    .D(_00409_),
    .Q(\decode.id_ex_rs2_data_reg[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27381_ (.CLK(clock),
    .D(_00410_),
    .Q(\decode.id_ex_rs2_data_reg[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27382_ (.CLK(clock),
    .D(_00411_),
    .Q(\decode.id_ex_rs2_data_reg[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27383_ (.CLK(clock),
    .D(_00412_),
    .Q(\decode.id_ex_rs2_data_reg[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27384_ (.CLK(clock),
    .D(_00413_),
    .Q(\decode.id_ex_rs2_data_reg[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27385_ (.CLK(clock),
    .D(_00414_),
    .Q(\decode.id_ex_rs2_data_reg[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27386_ (.CLK(clock),
    .D(_00415_),
    .Q(\decode.id_ex_rs2_data_reg[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27387_ (.CLK(clock),
    .D(_00416_),
    .Q(\decode.id_ex_rs2_data_reg[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27388_ (.CLK(clock),
    .D(_00417_),
    .Q(\decode.id_ex_rs2_data_reg[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27389_ (.CLK(clock),
    .D(_00418_),
    .Q(\decode.id_ex_rs2_data_reg[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27390_ (.CLK(clock),
    .D(_00419_),
    .Q(\decode.id_ex_rs2_data_reg[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27391_ (.CLK(clock),
    .D(_00420_),
    .Q(\decode.id_ex_rs1_data_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27392_ (.CLK(clock),
    .D(_00421_),
    .Q(\decode.id_ex_rs1_data_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27393_ (.CLK(clock),
    .D(_00422_),
    .Q(\decode.id_ex_rs1_data_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27394_ (.CLK(clock),
    .D(_00423_),
    .Q(\decode.id_ex_rs1_data_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27395_ (.CLK(clock),
    .D(_00424_),
    .Q(\decode.id_ex_rs1_data_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27396_ (.CLK(clock),
    .D(_00425_),
    .Q(\decode.id_ex_rs1_data_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27397_ (.CLK(clock),
    .D(_00426_),
    .Q(\decode.id_ex_rs1_data_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27398_ (.CLK(clock),
    .D(_00427_),
    .Q(\decode.id_ex_rs1_data_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27399_ (.CLK(clock),
    .D(_00428_),
    .Q(\decode.id_ex_rs1_data_reg[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27400_ (.CLK(clock),
    .D(_00429_),
    .Q(\decode.id_ex_rs1_data_reg[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27401_ (.CLK(clock),
    .D(_00430_),
    .Q(\decode.id_ex_rs1_data_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27402_ (.CLK(clock),
    .D(_00431_),
    .Q(\decode.id_ex_rs1_data_reg[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27403_ (.CLK(clock),
    .D(_00432_),
    .Q(\decode.id_ex_rs1_data_reg[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27404_ (.CLK(clock),
    .D(_00433_),
    .Q(\decode.id_ex_rs1_data_reg[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27405_ (.CLK(clock),
    .D(_00434_),
    .Q(\decode.id_ex_rs1_data_reg[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27406_ (.CLK(clock),
    .D(_00435_),
    .Q(\decode.id_ex_rs1_data_reg[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27407_ (.CLK(clock),
    .D(_00436_),
    .Q(\decode.id_ex_rs1_data_reg[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27408_ (.CLK(clock),
    .D(_00437_),
    .Q(\decode.id_ex_rs1_data_reg[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27409_ (.CLK(clock),
    .D(_00438_),
    .Q(\decode.id_ex_rs1_data_reg[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27410_ (.CLK(clock),
    .D(_00439_),
    .Q(\decode.id_ex_rs1_data_reg[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27411_ (.CLK(clock),
    .D(_00440_),
    .Q(\decode.id_ex_rs1_data_reg[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27412_ (.CLK(clock),
    .D(_00441_),
    .Q(\decode.id_ex_rs1_data_reg[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27413_ (.CLK(clock),
    .D(_00442_),
    .Q(\decode.id_ex_rs1_data_reg[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27414_ (.CLK(clock),
    .D(_00443_),
    .Q(\decode.id_ex_rs1_data_reg[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27415_ (.CLK(clock),
    .D(_00444_),
    .Q(\decode.id_ex_rs1_data_reg[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27416_ (.CLK(clock),
    .D(_00445_),
    .Q(\decode.id_ex_rs1_data_reg[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27417_ (.CLK(clock),
    .D(_00446_),
    .Q(\decode.id_ex_rs1_data_reg[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27418_ (.CLK(clock),
    .D(_00447_),
    .Q(\decode.id_ex_rs1_data_reg[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27419_ (.CLK(clock),
    .D(_00448_),
    .Q(\decode.id_ex_rs1_data_reg[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27420_ (.CLK(clock),
    .D(_00449_),
    .Q(\decode.id_ex_rs1_data_reg[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27421_ (.CLK(clock),
    .D(_00450_),
    .Q(\decode.id_ex_rs1_data_reg[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27422_ (.CLK(clock),
    .D(_00451_),
    .Q(\decode.id_ex_rs1_data_reg[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27423_ (.CLK(clock),
    .D(_00452_),
    .Q(\decode.id_ex_islui_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27424_ (.CLK(clock),
    .D(_00453_),
    .Q(\decode.id_ex_isjump_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27425_ (.CLK(clock),
    .D(_00454_),
    .Q(\decode.id_ex_rdsel_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27426_ (.CLK(clock),
    .D(_00455_),
    .Q(\decode.id_ex_pcsel_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27427_ (.CLK(clock),
    .D(_00456_),
    .Q(\decode.id_ex_memtoreg_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27428_ (.CLK(clock),
    .D(_00457_),
    .Q(\decode.id_ex_memtoreg_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27429_ (.CLK(clock),
    .D(_00458_),
    .Q(\decode.id_ex_regwrite_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27430_ (.CLK(clock),
    .D(_00459_),
    .Q(\decode.id_ex_memwrite_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27431_ (.CLK(clock),
    .D(_00460_),
    .Q(\decode.id_ex_memread_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27432_ (.CLK(clock),
    .D(_00461_),
    .Q(\decode.id_ex_isbranch_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27433_ (.CLK(clock),
    .D(_00462_),
    .Q(\decode.id_ex_immsrc_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27434_ (.CLK(clock),
    .D(_00463_),
    .Q(\decode.id_ex_pc_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27435_ (.CLK(clock),
    .D(_00464_),
    .Q(\decode.id_ex_pc_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27436_ (.CLK(clock),
    .D(_00465_),
    .Q(\decode.id_ex_pc_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27437_ (.CLK(clock),
    .D(_00466_),
    .Q(\decode.id_ex_pc_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27438_ (.CLK(clock),
    .D(_00467_),
    .Q(\decode.id_ex_pc_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27439_ (.CLK(clock),
    .D(_00468_),
    .Q(\decode.id_ex_pc_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27440_ (.CLK(clock),
    .D(_00469_),
    .Q(\decode.id_ex_pc_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27441_ (.CLK(clock),
    .D(_00470_),
    .Q(\decode.id_ex_pc_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27442_ (.CLK(clock),
    .D(_00471_),
    .Q(\decode.id_ex_pc_reg[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27443_ (.CLK(clock),
    .D(_00472_),
    .Q(\decode.id_ex_pc_reg[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27444_ (.CLK(clock),
    .D(_00473_),
    .Q(\decode.id_ex_pc_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27445_ (.CLK(clock),
    .D(_00474_),
    .Q(\decode.id_ex_pc_reg[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27446_ (.CLK(clock),
    .D(_00475_),
    .Q(\decode.id_ex_pc_reg[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27447_ (.CLK(clock),
    .D(_00476_),
    .Q(\decode.id_ex_pc_reg[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27448_ (.CLK(clock),
    .D(_00477_),
    .Q(\decode.id_ex_pc_reg[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27449_ (.CLK(clock),
    .D(_00478_),
    .Q(\decode.id_ex_pc_reg[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27450_ (.CLK(clock),
    .D(_00479_),
    .Q(\decode.id_ex_pc_reg[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27451_ (.CLK(clock),
    .D(_00480_),
    .Q(\decode.id_ex_pc_reg[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27452_ (.CLK(clock),
    .D(_00481_),
    .Q(\decode.id_ex_pc_reg[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27453_ (.CLK(clock),
    .D(_00482_),
    .Q(\decode.id_ex_pc_reg[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27454_ (.CLK(clock),
    .D(_00483_),
    .Q(\decode.id_ex_pc_reg[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27455_ (.CLK(clock),
    .D(_00484_),
    .Q(\decode.id_ex_pc_reg[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27456_ (.CLK(clock),
    .D(_00485_),
    .Q(\decode.id_ex_pc_reg[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27457_ (.CLK(clock),
    .D(_00486_),
    .Q(\decode.id_ex_pc_reg[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27458_ (.CLK(clock),
    .D(_00487_),
    .Q(\decode.id_ex_pc_reg[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27459_ (.CLK(clock),
    .D(_00488_),
    .Q(\decode.id_ex_pc_reg[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27460_ (.CLK(clock),
    .D(_00489_),
    .Q(\decode.id_ex_pc_reg[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27461_ (.CLK(clock),
    .D(_00490_),
    .Q(\decode.id_ex_pc_reg[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27462_ (.CLK(clock),
    .D(_00491_),
    .Q(\decode.id_ex_pc_reg[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27463_ (.CLK(clock),
    .D(_00492_),
    .Q(\decode.id_ex_pc_reg[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27464_ (.CLK(clock),
    .D(_00493_),
    .Q(\decode.id_ex_pc_reg[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27465_ (.CLK(clock),
    .D(_00494_),
    .Q(\decode.id_ex_pc_reg[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27466_ (.CLK(clock),
    .D(_00495_),
    .Q(\csr.io_csr_address[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27467_ (.CLK(clock),
    .D(_00496_),
    .Q(\csr.io_csr_address[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27468_ (.CLK(clock),
    .D(_00497_),
    .Q(\csr.io_csr_address[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27469_ (.CLK(clock),
    .D(_00498_),
    .Q(\csr.io_csr_address[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27470_ (.CLK(clock),
    .D(_00499_),
    .Q(\csr.io_csr_address[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27471_ (.CLK(clock),
    .D(_00500_),
    .Q(\csr.io_csr_address[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27472_ (.CLK(clock),
    .D(_00501_),
    .Q(\csr.io_csr_address[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27473_ (.CLK(clock),
    .D(_00502_),
    .Q(\csr.io_csr_address[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27474_ (.CLK(clock),
    .D(_00503_),
    .Q(\csr.io_csr_address[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27475_ (.CLK(clock),
    .D(_00504_),
    .Q(\csr.io_csr_address[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27476_ (.CLK(clock),
    .D(_00505_),
    .Q(\csr.io_csr_address[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27477_ (.CLK(clock),
    .D(_00506_),
    .Q(\csr.io_csr_address[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27478_ (.CLK(clock),
    .D(_00507_),
    .Q(\decode.csr_write_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27479_ (.CLK(clock),
    .D(_00508_),
    .Q(\decode.csr_read_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27480_ (.CLK(clock),
    .D(_00509_),
    .Q(\decode.exception_out_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27481_ (.CLK(clock),
    .D(_00510_),
    .Q(\decode.io_wfi_out ));
 sky130_fd_sc_hd__dfxtp_2 _27482_ (.CLK(clock),
    .D(_00511_),
    .Q(\decode.io_mret_out ));
 sky130_fd_sc_hd__dfxtp_2 _27483_ (.CLK(clock),
    .D(_00512_),
    .Q(\csr.mtip ));
 sky130_fd_sc_hd__dfxtp_2 _27484_ (.CLK(clock),
    .D(_00513_),
    .Q(io_memory_size[0]));
 sky130_fd_sc_hd__dfxtp_2 _27485_ (.CLK(clock),
    .D(_00514_),
    .Q(io_memory_size[1]));
 sky130_fd_sc_hd__dfxtp_2 _27486_ (.CLK(clock),
    .D(_00515_),
    .Q(io_load_store_unsigned));
 sky130_fd_sc_hd__dfxtp_2 _27487_ (.CLK(clock),
    .D(_00516_),
    .Q(io_memory_write_data[0]));
 sky130_fd_sc_hd__dfxtp_2 _27488_ (.CLK(clock),
    .D(_00517_),
    .Q(io_memory_write_data[1]));
 sky130_fd_sc_hd__dfxtp_2 _27489_ (.CLK(clock),
    .D(_00518_),
    .Q(io_memory_write_data[2]));
 sky130_fd_sc_hd__dfxtp_2 _27490_ (.CLK(clock),
    .D(_00519_),
    .Q(io_memory_write_data[3]));
 sky130_fd_sc_hd__dfxtp_2 _27491_ (.CLK(clock),
    .D(_00520_),
    .Q(io_memory_write_data[4]));
 sky130_fd_sc_hd__dfxtp_2 _27492_ (.CLK(clock),
    .D(_00521_),
    .Q(io_memory_write_data[5]));
 sky130_fd_sc_hd__dfxtp_2 _27493_ (.CLK(clock),
    .D(_00522_),
    .Q(io_memory_write_data[6]));
 sky130_fd_sc_hd__dfxtp_2 _27494_ (.CLK(clock),
    .D(_00523_),
    .Q(io_memory_write_data[7]));
 sky130_fd_sc_hd__dfxtp_2 _27495_ (.CLK(clock),
    .D(_00524_),
    .Q(io_memory_write_data[8]));
 sky130_fd_sc_hd__dfxtp_2 _27496_ (.CLK(clock),
    .D(_00525_),
    .Q(io_memory_write_data[9]));
 sky130_fd_sc_hd__dfxtp_2 _27497_ (.CLK(clock),
    .D(_00526_),
    .Q(io_memory_write_data[10]));
 sky130_fd_sc_hd__dfxtp_2 _27498_ (.CLK(clock),
    .D(_00527_),
    .Q(io_memory_write_data[11]));
 sky130_fd_sc_hd__dfxtp_2 _27499_ (.CLK(clock),
    .D(_00528_),
    .Q(io_memory_write_data[12]));
 sky130_fd_sc_hd__dfxtp_2 _27500_ (.CLK(clock),
    .D(_00529_),
    .Q(io_memory_write_data[13]));
 sky130_fd_sc_hd__dfxtp_2 _27501_ (.CLK(clock),
    .D(_00530_),
    .Q(io_memory_write_data[14]));
 sky130_fd_sc_hd__dfxtp_2 _27502_ (.CLK(clock),
    .D(_00531_),
    .Q(io_memory_write_data[15]));
 sky130_fd_sc_hd__dfxtp_2 _27503_ (.CLK(clock),
    .D(_00532_),
    .Q(io_memory_write_data[16]));
 sky130_fd_sc_hd__dfxtp_2 _27504_ (.CLK(clock),
    .D(_00533_),
    .Q(io_memory_write_data[17]));
 sky130_fd_sc_hd__dfxtp_2 _27505_ (.CLK(clock),
    .D(_00534_),
    .Q(io_memory_write_data[18]));
 sky130_fd_sc_hd__dfxtp_2 _27506_ (.CLK(clock),
    .D(_00535_),
    .Q(io_memory_write_data[19]));
 sky130_fd_sc_hd__dfxtp_2 _27507_ (.CLK(clock),
    .D(_00536_),
    .Q(io_memory_write_data[20]));
 sky130_fd_sc_hd__dfxtp_2 _27508_ (.CLK(clock),
    .D(_00537_),
    .Q(io_memory_write_data[21]));
 sky130_fd_sc_hd__dfxtp_2 _27509_ (.CLK(clock),
    .D(_00538_),
    .Q(io_memory_write_data[22]));
 sky130_fd_sc_hd__dfxtp_2 _27510_ (.CLK(clock),
    .D(_00539_),
    .Q(io_memory_write_data[23]));
 sky130_fd_sc_hd__dfxtp_2 _27511_ (.CLK(clock),
    .D(_00540_),
    .Q(io_memory_write_data[24]));
 sky130_fd_sc_hd__dfxtp_2 _27512_ (.CLK(clock),
    .D(_00541_),
    .Q(io_memory_write_data[25]));
 sky130_fd_sc_hd__dfxtp_2 _27513_ (.CLK(clock),
    .D(_00542_),
    .Q(io_memory_write_data[26]));
 sky130_fd_sc_hd__dfxtp_2 _27514_ (.CLK(clock),
    .D(_00543_),
    .Q(io_memory_write_data[27]));
 sky130_fd_sc_hd__dfxtp_2 _27515_ (.CLK(clock),
    .D(_00544_),
    .Q(io_memory_write_data[28]));
 sky130_fd_sc_hd__dfxtp_2 _27516_ (.CLK(clock),
    .D(_00545_),
    .Q(io_memory_write_data[29]));
 sky130_fd_sc_hd__dfxtp_2 _27517_ (.CLK(clock),
    .D(_00546_),
    .Q(io_memory_write_data[30]));
 sky130_fd_sc_hd__dfxtp_2 _27518_ (.CLK(clock),
    .D(_00547_),
    .Q(io_memory_write_data[31]));
 sky130_fd_sc_hd__dfxtp_2 _27519_ (.CLK(clock),
    .D(_00548_),
    .Q(io_memory_address[0]));
 sky130_fd_sc_hd__dfxtp_2 _27520_ (.CLK(clock),
    .D(_00549_),
    .Q(io_memory_address[1]));
 sky130_fd_sc_hd__dfxtp_2 _27521_ (.CLK(clock),
    .D(_00550_),
    .Q(io_memory_address[2]));
 sky130_fd_sc_hd__dfxtp_2 _27522_ (.CLK(clock),
    .D(_00551_),
    .Q(io_memory_address[3]));
 sky130_fd_sc_hd__dfxtp_2 _27523_ (.CLK(clock),
    .D(_00552_),
    .Q(io_memory_address[4]));
 sky130_fd_sc_hd__dfxtp_2 _27524_ (.CLK(clock),
    .D(_00553_),
    .Q(io_memory_address[5]));
 sky130_fd_sc_hd__dfxtp_2 _27525_ (.CLK(clock),
    .D(_00554_),
    .Q(io_memory_address[6]));
 sky130_fd_sc_hd__dfxtp_2 _27526_ (.CLK(clock),
    .D(_00555_),
    .Q(io_memory_address[7]));
 sky130_fd_sc_hd__dfxtp_2 _27527_ (.CLK(clock),
    .D(_00556_),
    .Q(io_memory_address[8]));
 sky130_fd_sc_hd__dfxtp_2 _27528_ (.CLK(clock),
    .D(_00557_),
    .Q(io_memory_address[9]));
 sky130_fd_sc_hd__dfxtp_2 _27529_ (.CLK(clock),
    .D(_00558_),
    .Q(io_memory_address[10]));
 sky130_fd_sc_hd__dfxtp_2 _27530_ (.CLK(clock),
    .D(_00559_),
    .Q(io_memory_address[11]));
 sky130_fd_sc_hd__dfxtp_2 _27531_ (.CLK(clock),
    .D(_00560_),
    .Q(io_memory_address[12]));
 sky130_fd_sc_hd__dfxtp_2 _27532_ (.CLK(clock),
    .D(_00561_),
    .Q(io_memory_address[13]));
 sky130_fd_sc_hd__dfxtp_2 _27533_ (.CLK(clock),
    .D(_00562_),
    .Q(io_memory_address[14]));
 sky130_fd_sc_hd__dfxtp_2 _27534_ (.CLK(clock),
    .D(_00563_),
    .Q(io_memory_address[15]));
 sky130_fd_sc_hd__dfxtp_2 _27535_ (.CLK(clock),
    .D(_00564_),
    .Q(io_memory_address[16]));
 sky130_fd_sc_hd__dfxtp_2 _27536_ (.CLK(clock),
    .D(_00565_),
    .Q(io_memory_address[17]));
 sky130_fd_sc_hd__dfxtp_2 _27537_ (.CLK(clock),
    .D(_00566_),
    .Q(io_memory_address[18]));
 sky130_fd_sc_hd__dfxtp_2 _27538_ (.CLK(clock),
    .D(_00567_),
    .Q(io_memory_address[19]));
 sky130_fd_sc_hd__dfxtp_2 _27539_ (.CLK(clock),
    .D(_00568_),
    .Q(io_memory_address[20]));
 sky130_fd_sc_hd__dfxtp_2 _27540_ (.CLK(clock),
    .D(_00569_),
    .Q(io_memory_address[21]));
 sky130_fd_sc_hd__dfxtp_2 _27541_ (.CLK(clock),
    .D(_00570_),
    .Q(io_memory_address[22]));
 sky130_fd_sc_hd__dfxtp_2 _27542_ (.CLK(clock),
    .D(_00571_),
    .Q(io_memory_address[23]));
 sky130_fd_sc_hd__dfxtp_2 _27543_ (.CLK(clock),
    .D(_00572_),
    .Q(io_memory_address[24]));
 sky130_fd_sc_hd__dfxtp_2 _27544_ (.CLK(clock),
    .D(_00573_),
    .Q(io_memory_address[25]));
 sky130_fd_sc_hd__dfxtp_2 _27545_ (.CLK(clock),
    .D(_00574_),
    .Q(io_memory_address[26]));
 sky130_fd_sc_hd__dfxtp_2 _27546_ (.CLK(clock),
    .D(_00575_),
    .Q(io_memory_address[27]));
 sky130_fd_sc_hd__dfxtp_2 _27547_ (.CLK(clock),
    .D(_00576_),
    .Q(io_memory_address[28]));
 sky130_fd_sc_hd__dfxtp_2 _27548_ (.CLK(clock),
    .D(_00577_),
    .Q(io_memory_address[29]));
 sky130_fd_sc_hd__dfxtp_2 _27549_ (.CLK(clock),
    .D(_00578_),
    .Q(io_memory_address[30]));
 sky130_fd_sc_hd__dfxtp_2 _27550_ (.CLK(clock),
    .D(_00579_),
    .Q(io_memory_address[31]));
 sky130_fd_sc_hd__dfxtp_2 _27551_ (.CLK(clock),
    .D(_00580_),
    .Q(\execute.io_mem_zero ));
 sky130_fd_sc_hd__dfxtp_2 _27552_ (.CLK(clock),
    .D(_00581_),
    .Q(\execute.io_mem_memtoreg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27553_ (.CLK(clock),
    .D(_00582_),
    .Q(\execute.io_mem_memtoreg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27554_ (.CLK(clock),
    .D(_00583_),
    .Q(\execute.io_mem_regwrite ));
 sky130_fd_sc_hd__dfxtp_2 _27555_ (.CLK(clock),
    .D(_00584_),
    .Q(\execute.io_mem_memwrite ));
 sky130_fd_sc_hd__dfxtp_2 _27556_ (.CLK(clock),
    .D(_00585_),
    .Q(io_memory_read));
 sky130_fd_sc_hd__dfxtp_2 _27557_ (.CLK(clock),
    .D(_00586_),
    .Q(\execute.io_mem_isjump ));
 sky130_fd_sc_hd__dfxtp_2 _27558_ (.CLK(clock),
    .D(_00587_),
    .Q(\execute.io_mem_isbranch ));
 sky130_fd_sc_hd__dfxtp_2 _27559_ (.CLK(clock),
    .D(_00588_),
    .Q(\csr.io_mem_pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27560_ (.CLK(clock),
    .D(_00589_),
    .Q(\csr.io_mem_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27561_ (.CLK(clock),
    .D(_00590_),
    .Q(\csr.io_mem_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27562_ (.CLK(clock),
    .D(_00591_),
    .Q(\csr.io_mem_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27563_ (.CLK(clock),
    .D(_00592_),
    .Q(\csr.io_mem_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27564_ (.CLK(clock),
    .D(_00593_),
    .Q(\csr.io_mem_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27565_ (.CLK(clock),
    .D(_00594_),
    .Q(\csr.io_mem_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27566_ (.CLK(clock),
    .D(_00595_),
    .Q(\csr.io_mem_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27567_ (.CLK(clock),
    .D(_00596_),
    .Q(\csr.io_mem_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27568_ (.CLK(clock),
    .D(_00597_),
    .Q(\csr.io_mem_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27569_ (.CLK(clock),
    .D(_00598_),
    .Q(\csr.io_mem_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27570_ (.CLK(clock),
    .D(_00599_),
    .Q(\csr.io_mem_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27571_ (.CLK(clock),
    .D(_00600_),
    .Q(\csr.io_mem_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27572_ (.CLK(clock),
    .D(_00601_),
    .Q(\csr.io_mem_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27573_ (.CLK(clock),
    .D(_00602_),
    .Q(\csr.io_mem_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27574_ (.CLK(clock),
    .D(_00603_),
    .Q(\csr.io_mem_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27575_ (.CLK(clock),
    .D(_00604_),
    .Q(\csr.io_mem_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27576_ (.CLK(clock),
    .D(_00605_),
    .Q(\csr.io_mem_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27577_ (.CLK(clock),
    .D(_00606_),
    .Q(\csr.io_mem_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27578_ (.CLK(clock),
    .D(_00607_),
    .Q(\csr.io_mem_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27579_ (.CLK(clock),
    .D(_00608_),
    .Q(\csr.io_mem_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27580_ (.CLK(clock),
    .D(_00609_),
    .Q(\csr.io_mem_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27581_ (.CLK(clock),
    .D(_00610_),
    .Q(\csr.io_mem_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27582_ (.CLK(clock),
    .D(_00611_),
    .Q(\csr.io_mem_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27583_ (.CLK(clock),
    .D(_00612_),
    .Q(\csr.io_mem_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27584_ (.CLK(clock),
    .D(_00613_),
    .Q(\csr.io_mem_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27585_ (.CLK(clock),
    .D(_00614_),
    .Q(\csr.io_mem_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27586_ (.CLK(clock),
    .D(_00615_),
    .Q(\csr.io_mem_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27587_ (.CLK(clock),
    .D(_00616_),
    .Q(\csr.io_mem_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27588_ (.CLK(clock),
    .D(_00617_),
    .Q(\csr.io_mem_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27589_ (.CLK(clock),
    .D(_00618_),
    .Q(\csr.io_mem_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27590_ (.CLK(clock),
    .D(_00619_),
    .Q(\csr.io_mem_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27591_ (.CLK(clock),
    .D(_00620_),
    .Q(\execute.io_target_pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27592_ (.CLK(clock),
    .D(_00621_),
    .Q(\execute.io_target_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27593_ (.CLK(clock),
    .D(_00622_),
    .Q(\execute.io_target_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27594_ (.CLK(clock),
    .D(_00623_),
    .Q(\execute.io_target_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27595_ (.CLK(clock),
    .D(_00624_),
    .Q(\execute.io_target_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27596_ (.CLK(clock),
    .D(_00625_),
    .Q(\execute.io_target_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27597_ (.CLK(clock),
    .D(_00626_),
    .Q(\execute.io_target_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27598_ (.CLK(clock),
    .D(_00627_),
    .Q(\execute.io_target_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27599_ (.CLK(clock),
    .D(_00628_),
    .Q(\execute.io_target_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27600_ (.CLK(clock),
    .D(_00629_),
    .Q(\execute.io_target_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27601_ (.CLK(clock),
    .D(_00630_),
    .Q(\execute.io_target_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27602_ (.CLK(clock),
    .D(_00631_),
    .Q(\execute.io_target_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27603_ (.CLK(clock),
    .D(_00632_),
    .Q(\execute.io_target_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27604_ (.CLK(clock),
    .D(_00633_),
    .Q(\execute.io_target_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27605_ (.CLK(clock),
    .D(_00634_),
    .Q(\execute.io_target_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27606_ (.CLK(clock),
    .D(_00635_),
    .Q(\execute.io_target_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27607_ (.CLK(clock),
    .D(_00636_),
    .Q(\execute.io_target_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27608_ (.CLK(clock),
    .D(_00637_),
    .Q(\execute.io_target_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27609_ (.CLK(clock),
    .D(_00638_),
    .Q(\execute.io_target_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27610_ (.CLK(clock),
    .D(_00639_),
    .Q(\execute.io_target_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27611_ (.CLK(clock),
    .D(_00640_),
    .Q(\execute.io_target_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27612_ (.CLK(clock),
    .D(_00641_),
    .Q(\execute.io_target_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27613_ (.CLK(clock),
    .D(_00642_),
    .Q(\execute.io_target_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27614_ (.CLK(clock),
    .D(_00643_),
    .Q(\execute.io_target_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27615_ (.CLK(clock),
    .D(_00644_),
    .Q(\execute.io_target_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27616_ (.CLK(clock),
    .D(_00645_),
    .Q(\execute.io_target_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27617_ (.CLK(clock),
    .D(_00646_),
    .Q(\execute.io_target_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27618_ (.CLK(clock),
    .D(_00647_),
    .Q(\execute.io_target_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27619_ (.CLK(clock),
    .D(_00648_),
    .Q(\execute.io_target_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27620_ (.CLK(clock),
    .D(_00649_),
    .Q(\execute.io_target_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27621_ (.CLK(clock),
    .D(_00650_),
    .Q(\execute.io_target_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27622_ (.CLK(clock),
    .D(_00651_),
    .Q(\execute.io_target_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27623_ (.CLK(clock),
    .D(_00652_),
    .Q(\execute.io_reg_pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27624_ (.CLK(clock),
    .D(_00653_),
    .Q(\execute.io_reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27625_ (.CLK(clock),
    .D(_00654_),
    .Q(\execute.io_reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27626_ (.CLK(clock),
    .D(_00655_),
    .Q(\execute.io_reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27627_ (.CLK(clock),
    .D(_00656_),
    .Q(\execute.io_reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27628_ (.CLK(clock),
    .D(_00657_),
    .Q(\execute.io_reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27629_ (.CLK(clock),
    .D(_00658_),
    .Q(\execute.io_reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27630_ (.CLK(clock),
    .D(_00659_),
    .Q(\execute.io_reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27631_ (.CLK(clock),
    .D(_00660_),
    .Q(\execute.io_reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27632_ (.CLK(clock),
    .D(_00661_),
    .Q(\execute.io_reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27633_ (.CLK(clock),
    .D(_00662_),
    .Q(\execute.io_reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27634_ (.CLK(clock),
    .D(_00663_),
    .Q(\execute.io_reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27635_ (.CLK(clock),
    .D(_00664_),
    .Q(\execute.io_reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27636_ (.CLK(clock),
    .D(_00665_),
    .Q(\execute.io_reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27637_ (.CLK(clock),
    .D(_00666_),
    .Q(\execute.io_reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27638_ (.CLK(clock),
    .D(_00667_),
    .Q(\execute.io_reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27639_ (.CLK(clock),
    .D(_00668_),
    .Q(\execute.io_reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27640_ (.CLK(clock),
    .D(_00669_),
    .Q(\execute.io_reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27641_ (.CLK(clock),
    .D(_00670_),
    .Q(\execute.io_reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27642_ (.CLK(clock),
    .D(_00671_),
    .Q(\execute.io_reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27643_ (.CLK(clock),
    .D(_00672_),
    .Q(\execute.io_reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27644_ (.CLK(clock),
    .D(_00673_),
    .Q(\execute.io_reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27645_ (.CLK(clock),
    .D(_00674_),
    .Q(\execute.io_reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27646_ (.CLK(clock),
    .D(_00675_),
    .Q(\execute.io_reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27647_ (.CLK(clock),
    .D(_00676_),
    .Q(\execute.io_reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27648_ (.CLK(clock),
    .D(_00677_),
    .Q(\execute.io_reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27649_ (.CLK(clock),
    .D(_00678_),
    .Q(\execute.io_reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27650_ (.CLK(clock),
    .D(_00679_),
    .Q(\execute.io_reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27651_ (.CLK(clock),
    .D(_00680_),
    .Q(\execute.io_reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27652_ (.CLK(clock),
    .D(_00681_),
    .Q(\execute.io_reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27653_ (.CLK(clock),
    .D(_00682_),
    .Q(\execute.io_reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27654_ (.CLK(clock),
    .D(_00683_),
    .Q(\execute.io_reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27655_ (.CLK(clock),
    .D(_00684_),
    .Q(\execute.exception_out_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27656_ (.CLK(clock),
    .D(_00685_),
    .Q(\execute.io_wfi_out ));
 sky130_fd_sc_hd__dfxtp_2 _27657_ (.CLK(clock),
    .D(_00686_),
    .Q(\execute.io_mret_out ));
 sky130_fd_sc_hd__dfxtp_2 _27658_ (.CLK(clock),
    .D(_00687_),
    .Q(\execute.csr_read_data_out_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27659_ (.CLK(clock),
    .D(_00688_),
    .Q(\execute.csr_read_data_out_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27660_ (.CLK(clock),
    .D(_00689_),
    .Q(\execute.csr_read_data_out_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27661_ (.CLK(clock),
    .D(_00690_),
    .Q(\execute.csr_read_data_out_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27662_ (.CLK(clock),
    .D(_00691_),
    .Q(\execute.csr_read_data_out_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27663_ (.CLK(clock),
    .D(_00692_),
    .Q(\execute.csr_read_data_out_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27664_ (.CLK(clock),
    .D(_00693_),
    .Q(\execute.csr_read_data_out_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27665_ (.CLK(clock),
    .D(_00694_),
    .Q(\execute.csr_read_data_out_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27666_ (.CLK(clock),
    .D(_00695_),
    .Q(\execute.csr_read_data_out_reg[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27667_ (.CLK(clock),
    .D(_00696_),
    .Q(\execute.csr_read_data_out_reg[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27668_ (.CLK(clock),
    .D(_00697_),
    .Q(\execute.csr_read_data_out_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27669_ (.CLK(clock),
    .D(_00698_),
    .Q(\execute.csr_read_data_out_reg[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27670_ (.CLK(clock),
    .D(_00699_),
    .Q(\execute.csr_read_data_out_reg[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27671_ (.CLK(clock),
    .D(_00700_),
    .Q(\execute.csr_read_data_out_reg[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27672_ (.CLK(clock),
    .D(_00701_),
    .Q(\execute.csr_read_data_out_reg[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27673_ (.CLK(clock),
    .D(_00702_),
    .Q(\execute.csr_read_data_out_reg[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27674_ (.CLK(clock),
    .D(_00703_),
    .Q(\execute.csr_read_data_out_reg[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27675_ (.CLK(clock),
    .D(_00704_),
    .Q(\execute.csr_read_data_out_reg[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27676_ (.CLK(clock),
    .D(_00705_),
    .Q(\execute.csr_read_data_out_reg[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27677_ (.CLK(clock),
    .D(_00706_),
    .Q(\execute.csr_read_data_out_reg[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27678_ (.CLK(clock),
    .D(_00707_),
    .Q(\execute.csr_read_data_out_reg[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27679_ (.CLK(clock),
    .D(_00708_),
    .Q(\execute.csr_read_data_out_reg[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27680_ (.CLK(clock),
    .D(_00709_),
    .Q(\execute.csr_read_data_out_reg[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27681_ (.CLK(clock),
    .D(_00710_),
    .Q(\execute.csr_read_data_out_reg[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27682_ (.CLK(clock),
    .D(_00711_),
    .Q(\execute.csr_read_data_out_reg[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27683_ (.CLK(clock),
    .D(_00712_),
    .Q(\execute.csr_read_data_out_reg[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27684_ (.CLK(clock),
    .D(_00713_),
    .Q(\execute.csr_read_data_out_reg[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27685_ (.CLK(clock),
    .D(_00714_),
    .Q(\execute.csr_read_data_out_reg[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27686_ (.CLK(clock),
    .D(_00715_),
    .Q(\execute.csr_read_data_out_reg[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27687_ (.CLK(clock),
    .D(_00716_),
    .Q(\execute.csr_read_data_out_reg[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27688_ (.CLK(clock),
    .D(_00717_),
    .Q(\execute.csr_read_data_out_reg[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27689_ (.CLK(clock),
    .D(_00718_),
    .Q(\execute.csr_read_data_out_reg[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27690_ (.CLK(clock),
    .D(_00719_),
    .Q(\execute.csr_write_data_out_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27691_ (.CLK(clock),
    .D(_00720_),
    .Q(\execute.csr_write_data_out_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27692_ (.CLK(clock),
    .D(_00721_),
    .Q(\execute.csr_write_data_out_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27693_ (.CLK(clock),
    .D(_00722_),
    .Q(\execute.csr_write_data_out_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27694_ (.CLK(clock),
    .D(_00723_),
    .Q(\execute.csr_write_data_out_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27695_ (.CLK(clock),
    .D(_00724_),
    .Q(\execute.csr_write_data_out_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27696_ (.CLK(clock),
    .D(_00725_),
    .Q(\execute.csr_write_data_out_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27697_ (.CLK(clock),
    .D(_00726_),
    .Q(\execute.csr_write_data_out_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27698_ (.CLK(clock),
    .D(_00727_),
    .Q(\execute.csr_write_data_out_reg[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27699_ (.CLK(clock),
    .D(_00728_),
    .Q(\execute.csr_write_data_out_reg[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27700_ (.CLK(clock),
    .D(_00729_),
    .Q(\execute.csr_write_data_out_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27701_ (.CLK(clock),
    .D(_00730_),
    .Q(\execute.csr_write_data_out_reg[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27702_ (.CLK(clock),
    .D(_00731_),
    .Q(\execute.csr_write_data_out_reg[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27703_ (.CLK(clock),
    .D(_00732_),
    .Q(\execute.csr_write_data_out_reg[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27704_ (.CLK(clock),
    .D(_00733_),
    .Q(\execute.csr_write_data_out_reg[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27705_ (.CLK(clock),
    .D(_00734_),
    .Q(\execute.csr_write_data_out_reg[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27706_ (.CLK(clock),
    .D(_00735_),
    .Q(\execute.csr_write_data_out_reg[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27707_ (.CLK(clock),
    .D(_00736_),
    .Q(\execute.csr_write_data_out_reg[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27708_ (.CLK(clock),
    .D(_00737_),
    .Q(\execute.csr_write_data_out_reg[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27709_ (.CLK(clock),
    .D(_00738_),
    .Q(\execute.csr_write_data_out_reg[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27710_ (.CLK(clock),
    .D(_00739_),
    .Q(\execute.csr_write_data_out_reg[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27711_ (.CLK(clock),
    .D(_00740_),
    .Q(\execute.csr_write_data_out_reg[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27712_ (.CLK(clock),
    .D(_00741_),
    .Q(\execute.csr_write_data_out_reg[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27713_ (.CLK(clock),
    .D(_00742_),
    .Q(\execute.csr_write_data_out_reg[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27714_ (.CLK(clock),
    .D(_00743_),
    .Q(\execute.csr_write_data_out_reg[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27715_ (.CLK(clock),
    .D(_00744_),
    .Q(\execute.csr_write_data_out_reg[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27716_ (.CLK(clock),
    .D(_00745_),
    .Q(\execute.csr_write_data_out_reg[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27717_ (.CLK(clock),
    .D(_00746_),
    .Q(\execute.csr_write_data_out_reg[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27718_ (.CLK(clock),
    .D(_00747_),
    .Q(\execute.csr_write_data_out_reg[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27719_ (.CLK(clock),
    .D(_00748_),
    .Q(\execute.csr_write_data_out_reg[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27720_ (.CLK(clock),
    .D(_00749_),
    .Q(\execute.csr_write_data_out_reg[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27721_ (.CLK(clock),
    .D(_00750_),
    .Q(\execute.csr_write_data_out_reg[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27722_ (.CLK(clock),
    .D(_00751_),
    .Q(\execute.csr_write_address_out_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27723_ (.CLK(clock),
    .D(_00752_),
    .Q(\execute.csr_write_address_out_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27724_ (.CLK(clock),
    .D(_00753_),
    .Q(\execute.csr_write_address_out_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27725_ (.CLK(clock),
    .D(_00754_),
    .Q(\execute.csr_write_address_out_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27726_ (.CLK(clock),
    .D(_00755_),
    .Q(\execute.csr_write_address_out_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27727_ (.CLK(clock),
    .D(_00756_),
    .Q(\execute.csr_write_address_out_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27728_ (.CLK(clock),
    .D(_00757_),
    .Q(\execute.csr_write_address_out_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27729_ (.CLK(clock),
    .D(_00758_),
    .Q(\execute.csr_write_address_out_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27730_ (.CLK(clock),
    .D(_00759_),
    .Q(\execute.csr_write_address_out_reg[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27731_ (.CLK(clock),
    .D(_00760_),
    .Q(\execute.csr_write_address_out_reg[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27732_ (.CLK(clock),
    .D(_00761_),
    .Q(\execute.csr_write_address_out_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27733_ (.CLK(clock),
    .D(_00762_),
    .Q(\execute.csr_write_address_out_reg[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27734_ (.CLK(clock),
    .D(_00763_),
    .Q(\execute.csr_write_enable_out_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27735_ (.CLK(clock),
    .D(_00764_),
    .Q(\decode.id_ex_ex_use_rs2_reg ));
 sky130_fd_sc_hd__dfxtp_2 _27736_ (.CLK(clock),
    .D(_00765_),
    .Q(\fetch.bht.bhtTable_tag_MPORT_en ));
 sky130_fd_sc_hd__dfxtp_2 _27737_ (.CLK(clock),
    .D(_00766_),
    .Q(\decode.io_wb_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27738_ (.CLK(clock),
    .D(_00767_),
    .Q(\decode.io_wb_rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27739_ (.CLK(clock),
    .D(_00768_),
    .Q(\decode.io_wb_rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27740_ (.CLK(clock),
    .D(_00769_),
    .Q(\decode.io_wb_rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27741_ (.CLK(clock),
    .D(_00770_),
    .Q(\decode.io_wb_rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27742_ (.CLK(clock),
    .D(_00771_),
    .Q(\decode.io_wb_regwrite ));
 sky130_fd_sc_hd__dfxtp_2 _27743_ (.CLK(clock),
    .D(_00772_),
    .Q(\memory.io_wb_memtoreg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27744_ (.CLK(clock),
    .D(_00773_),
    .Q(\memory.io_wb_memtoreg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27745_ (.CLK(clock),
    .D(_00774_),
    .Q(\memory.io_wb_aluresult[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27746_ (.CLK(clock),
    .D(_00775_),
    .Q(\memory.io_wb_aluresult[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27747_ (.CLK(clock),
    .D(_00776_),
    .Q(\memory.io_wb_aluresult[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27748_ (.CLK(clock),
    .D(_00777_),
    .Q(\memory.io_wb_aluresult[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27749_ (.CLK(clock),
    .D(_00778_),
    .Q(\memory.io_wb_aluresult[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27750_ (.CLK(clock),
    .D(_00779_),
    .Q(\memory.io_wb_aluresult[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27751_ (.CLK(clock),
    .D(_00780_),
    .Q(\memory.io_wb_aluresult[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27752_ (.CLK(clock),
    .D(_00781_),
    .Q(\memory.io_wb_aluresult[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27753_ (.CLK(clock),
    .D(_00782_),
    .Q(\memory.io_wb_aluresult[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27754_ (.CLK(clock),
    .D(_00783_),
    .Q(\memory.io_wb_aluresult[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27755_ (.CLK(clock),
    .D(_00784_),
    .Q(\memory.io_wb_aluresult[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27756_ (.CLK(clock),
    .D(_00785_),
    .Q(\memory.io_wb_aluresult[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27757_ (.CLK(clock),
    .D(_00786_),
    .Q(\memory.io_wb_aluresult[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27758_ (.CLK(clock),
    .D(_00787_),
    .Q(\memory.io_wb_aluresult[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27759_ (.CLK(clock),
    .D(_00788_),
    .Q(\memory.io_wb_aluresult[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27760_ (.CLK(clock),
    .D(_00789_),
    .Q(\memory.io_wb_aluresult[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27761_ (.CLK(clock),
    .D(_00790_),
    .Q(\memory.io_wb_aluresult[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27762_ (.CLK(clock),
    .D(_00791_),
    .Q(\memory.io_wb_aluresult[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27763_ (.CLK(clock),
    .D(_00792_),
    .Q(\memory.io_wb_aluresult[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27764_ (.CLK(clock),
    .D(_00793_),
    .Q(\memory.io_wb_aluresult[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27765_ (.CLK(clock),
    .D(_00794_),
    .Q(\memory.io_wb_aluresult[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27766_ (.CLK(clock),
    .D(_00795_),
    .Q(\memory.io_wb_aluresult[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27767_ (.CLK(clock),
    .D(_00796_),
    .Q(\memory.io_wb_aluresult[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27768_ (.CLK(clock),
    .D(_00797_),
    .Q(\memory.io_wb_aluresult[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27769_ (.CLK(clock),
    .D(_00798_),
    .Q(\memory.io_wb_aluresult[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27770_ (.CLK(clock),
    .D(_00799_),
    .Q(\memory.io_wb_aluresult[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27771_ (.CLK(clock),
    .D(_00800_),
    .Q(\memory.io_wb_aluresult[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27772_ (.CLK(clock),
    .D(_00801_),
    .Q(\memory.io_wb_aluresult[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27773_ (.CLK(clock),
    .D(_00802_),
    .Q(\memory.io_wb_aluresult[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27774_ (.CLK(clock),
    .D(_00803_),
    .Q(\memory.io_wb_aluresult[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27775_ (.CLK(clock),
    .D(_00804_),
    .Q(\memory.io_wb_aluresult[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27776_ (.CLK(clock),
    .D(_00805_),
    .Q(\memory.io_wb_aluresult[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27777_ (.CLK(clock),
    .D(_00806_),
    .Q(\memory.io_wb_readdata[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27778_ (.CLK(clock),
    .D(_00807_),
    .Q(\memory.io_wb_readdata[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27779_ (.CLK(clock),
    .D(_00808_),
    .Q(\memory.io_wb_readdata[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27780_ (.CLK(clock),
    .D(_00809_),
    .Q(\memory.io_wb_readdata[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27781_ (.CLK(clock),
    .D(_00810_),
    .Q(\memory.io_wb_readdata[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27782_ (.CLK(clock),
    .D(_00811_),
    .Q(\memory.io_wb_readdata[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27783_ (.CLK(clock),
    .D(_00812_),
    .Q(\memory.io_wb_readdata[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27784_ (.CLK(clock),
    .D(_00813_),
    .Q(\memory.io_wb_readdata[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27785_ (.CLK(clock),
    .D(_00814_),
    .Q(\memory.io_wb_readdata[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27786_ (.CLK(clock),
    .D(_00815_),
    .Q(\memory.io_wb_readdata[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27787_ (.CLK(clock),
    .D(_00816_),
    .Q(\memory.io_wb_readdata[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27788_ (.CLK(clock),
    .D(_00817_),
    .Q(\memory.io_wb_readdata[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27789_ (.CLK(clock),
    .D(_00818_),
    .Q(\memory.io_wb_readdata[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27790_ (.CLK(clock),
    .D(_00819_),
    .Q(\memory.io_wb_readdata[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27791_ (.CLK(clock),
    .D(_00820_),
    .Q(\memory.io_wb_readdata[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27792_ (.CLK(clock),
    .D(_00821_),
    .Q(\memory.io_wb_readdata[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27793_ (.CLK(clock),
    .D(_00822_),
    .Q(\memory.io_wb_readdata[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27794_ (.CLK(clock),
    .D(_00823_),
    .Q(\memory.io_wb_readdata[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27795_ (.CLK(clock),
    .D(_00824_),
    .Q(\memory.io_wb_readdata[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27796_ (.CLK(clock),
    .D(_00825_),
    .Q(\memory.io_wb_readdata[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27797_ (.CLK(clock),
    .D(_00826_),
    .Q(\memory.io_wb_readdata[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27798_ (.CLK(clock),
    .D(_00827_),
    .Q(\memory.io_wb_readdata[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27799_ (.CLK(clock),
    .D(_00828_),
    .Q(\memory.io_wb_readdata[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27800_ (.CLK(clock),
    .D(_00829_),
    .Q(\memory.io_wb_readdata[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27801_ (.CLK(clock),
    .D(_00830_),
    .Q(\memory.io_wb_readdata[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27802_ (.CLK(clock),
    .D(_00831_),
    .Q(\memory.io_wb_readdata[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27803_ (.CLK(clock),
    .D(_00832_),
    .Q(\memory.io_wb_readdata[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27804_ (.CLK(clock),
    .D(_00833_),
    .Q(\memory.io_wb_readdata[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27805_ (.CLK(clock),
    .D(_00834_),
    .Q(\memory.io_wb_readdata[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27806_ (.CLK(clock),
    .D(_00835_),
    .Q(\memory.io_wb_readdata[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27807_ (.CLK(clock),
    .D(_00836_),
    .Q(\memory.io_wb_readdata[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27808_ (.CLK(clock),
    .D(_00837_),
    .Q(\memory.io_wb_readdata[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27809_ (.CLK(clock),
    .D(_00838_),
    .Q(\memory.io_wb_reg_pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27810_ (.CLK(clock),
    .D(_00839_),
    .Q(\memory.io_wb_reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27811_ (.CLK(clock),
    .D(_00840_),
    .Q(\memory.io_wb_reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27812_ (.CLK(clock),
    .D(_00841_),
    .Q(\memory.io_wb_reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27813_ (.CLK(clock),
    .D(_00842_),
    .Q(\memory.io_wb_reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27814_ (.CLK(clock),
    .D(_00843_),
    .Q(\memory.io_wb_reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27815_ (.CLK(clock),
    .D(_00844_),
    .Q(\memory.io_wb_reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27816_ (.CLK(clock),
    .D(_00845_),
    .Q(\memory.io_wb_reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27817_ (.CLK(clock),
    .D(_00846_),
    .Q(\memory.io_wb_reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27818_ (.CLK(clock),
    .D(_00847_),
    .Q(\memory.io_wb_reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27819_ (.CLK(clock),
    .D(_00848_),
    .Q(\memory.io_wb_reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27820_ (.CLK(clock),
    .D(_00849_),
    .Q(\memory.io_wb_reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27821_ (.CLK(clock),
    .D(_00850_),
    .Q(\memory.io_wb_reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27822_ (.CLK(clock),
    .D(_00851_),
    .Q(\memory.io_wb_reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27823_ (.CLK(clock),
    .D(_00852_),
    .Q(\memory.io_wb_reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27824_ (.CLK(clock),
    .D(_00853_),
    .Q(\memory.io_wb_reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27825_ (.CLK(clock),
    .D(_00854_),
    .Q(\memory.io_wb_reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27826_ (.CLK(clock),
    .D(_00855_),
    .Q(\memory.io_wb_reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27827_ (.CLK(clock),
    .D(_00856_),
    .Q(\memory.io_wb_reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27828_ (.CLK(clock),
    .D(_00857_),
    .Q(\memory.io_wb_reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27829_ (.CLK(clock),
    .D(_00858_),
    .Q(\memory.io_wb_reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27830_ (.CLK(clock),
    .D(_00859_),
    .Q(\memory.io_wb_reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27831_ (.CLK(clock),
    .D(_00860_),
    .Q(\memory.io_wb_reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27832_ (.CLK(clock),
    .D(_00861_),
    .Q(\memory.io_wb_reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27833_ (.CLK(clock),
    .D(_00862_),
    .Q(\memory.io_wb_reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27834_ (.CLK(clock),
    .D(_00863_),
    .Q(\memory.io_wb_reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27835_ (.CLK(clock),
    .D(_00864_),
    .Q(\memory.io_wb_reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27836_ (.CLK(clock),
    .D(_00865_),
    .Q(\memory.io_wb_reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27837_ (.CLK(clock),
    .D(_00866_),
    .Q(\memory.io_wb_reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27838_ (.CLK(clock),
    .D(_00867_),
    .Q(\memory.io_wb_reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27839_ (.CLK(clock),
    .D(_00868_),
    .Q(\memory.io_wb_reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27840_ (.CLK(clock),
    .D(_00869_),
    .Q(\memory.io_wb_reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27841_ (.CLK(clock),
    .D(_00870_),
    .Q(\csr.io_mret ));
 sky130_fd_sc_hd__dfxtp_2 _27842_ (.CLK(clock),
    .D(_00871_),
    .Q(\memory.csr_read_data_out_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27843_ (.CLK(clock),
    .D(_00872_),
    .Q(\memory.csr_read_data_out_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27844_ (.CLK(clock),
    .D(_00873_),
    .Q(\memory.csr_read_data_out_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27845_ (.CLK(clock),
    .D(_00874_),
    .Q(\memory.csr_read_data_out_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27846_ (.CLK(clock),
    .D(_00875_),
    .Q(\memory.csr_read_data_out_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27847_ (.CLK(clock),
    .D(_00876_),
    .Q(\memory.csr_read_data_out_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27848_ (.CLK(clock),
    .D(_00877_),
    .Q(\memory.csr_read_data_out_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27849_ (.CLK(clock),
    .D(_00878_),
    .Q(\memory.csr_read_data_out_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27850_ (.CLK(clock),
    .D(_00879_),
    .Q(\memory.csr_read_data_out_reg[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27851_ (.CLK(clock),
    .D(_00880_),
    .Q(\memory.csr_read_data_out_reg[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27852_ (.CLK(clock),
    .D(_00881_),
    .Q(\memory.csr_read_data_out_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27853_ (.CLK(clock),
    .D(_00882_),
    .Q(\memory.csr_read_data_out_reg[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27854_ (.CLK(clock),
    .D(_00883_),
    .Q(\memory.csr_read_data_out_reg[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27855_ (.CLK(clock),
    .D(_00884_),
    .Q(\memory.csr_read_data_out_reg[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27856_ (.CLK(clock),
    .D(_00885_),
    .Q(\memory.csr_read_data_out_reg[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27857_ (.CLK(clock),
    .D(_00886_),
    .Q(\memory.csr_read_data_out_reg[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27858_ (.CLK(clock),
    .D(_00887_),
    .Q(\memory.csr_read_data_out_reg[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27859_ (.CLK(clock),
    .D(_00888_),
    .Q(\memory.csr_read_data_out_reg[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27860_ (.CLK(clock),
    .D(_00889_),
    .Q(\memory.csr_read_data_out_reg[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27861_ (.CLK(clock),
    .D(_00890_),
    .Q(\memory.csr_read_data_out_reg[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27862_ (.CLK(clock),
    .D(_00891_),
    .Q(\memory.csr_read_data_out_reg[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27863_ (.CLK(clock),
    .D(_00892_),
    .Q(\memory.csr_read_data_out_reg[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27864_ (.CLK(clock),
    .D(_00893_),
    .Q(\memory.csr_read_data_out_reg[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27865_ (.CLK(clock),
    .D(_00894_),
    .Q(\memory.csr_read_data_out_reg[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27866_ (.CLK(clock),
    .D(_00895_),
    .Q(\memory.csr_read_data_out_reg[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27867_ (.CLK(clock),
    .D(_00896_),
    .Q(\memory.csr_read_data_out_reg[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27868_ (.CLK(clock),
    .D(_00897_),
    .Q(\memory.csr_read_data_out_reg[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27869_ (.CLK(clock),
    .D(_00898_),
    .Q(\memory.csr_read_data_out_reg[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27870_ (.CLK(clock),
    .D(_00899_),
    .Q(\memory.csr_read_data_out_reg[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27871_ (.CLK(clock),
    .D(_00900_),
    .Q(\memory.csr_read_data_out_reg[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27872_ (.CLK(clock),
    .D(_00901_),
    .Q(\memory.csr_read_data_out_reg[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27873_ (.CLK(clock),
    .D(_00902_),
    .Q(\memory.csr_read_data_out_reg[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27874_ (.CLK(clock),
    .D(_00903_),
    .Q(\csr.io_inst_retired ));
 sky130_fd_sc_hd__dfxtp_2 _27875_ (.CLK(clock),
    .D(_00904_),
    .Q(\csr.io_interrupt ));
 sky130_fd_sc_hd__dfxtp_2 _27876_ (.CLK(clock),
    .D(_00905_),
    .Q(\csr.io_trapped ));
 sky130_fd_sc_hd__dfxtp_2 _27877_ (.CLK(clock),
    .D(_00906_),
    .Q(\csr.io_ecause[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27878_ (.CLK(clock),
    .D(_00907_),
    .Q(\csr.io_ecause[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27879_ (.CLK(clock),
    .D(_00908_),
    .Q(\csr._mcycle_T_2[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27880_ (.CLK(clock),
    .D(_00909_),
    .Q(\csr._mcycle_T_2[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27881_ (.CLK(clock),
    .D(_00910_),
    .Q(\csr._mcycle_T_2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27882_ (.CLK(clock),
    .D(_00911_),
    .Q(\csr._mcycle_T_2[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27883_ (.CLK(clock),
    .D(_00912_),
    .Q(\csr._mcycle_T_2[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27884_ (.CLK(clock),
    .D(_00913_),
    .Q(\csr._mcycle_T_2[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27885_ (.CLK(clock),
    .D(_00914_),
    .Q(\csr._mcycle_T_2[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27886_ (.CLK(clock),
    .D(_00915_),
    .Q(\csr._mcycle_T_2[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27887_ (.CLK(clock),
    .D(_00916_),
    .Q(\csr._mcycle_T_2[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27888_ (.CLK(clock),
    .D(_00917_),
    .Q(\csr._mcycle_T_2[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27889_ (.CLK(clock),
    .D(_00918_),
    .Q(\csr._mcycle_T_2[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27890_ (.CLK(clock),
    .D(_00919_),
    .Q(\csr._mcycle_T_2[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27891_ (.CLK(clock),
    .D(_00920_),
    .Q(\csr._mcycle_T_2[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27892_ (.CLK(clock),
    .D(_00921_),
    .Q(\csr._mcycle_T_2[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27893_ (.CLK(clock),
    .D(_00922_),
    .Q(\csr._mcycle_T_2[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27894_ (.CLK(clock),
    .D(_00923_),
    .Q(\csr._mcycle_T_2[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27895_ (.CLK(clock),
    .D(_00924_),
    .Q(\csr._mcycle_T_2[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27896_ (.CLK(clock),
    .D(_00925_),
    .Q(\csr._mcycle_T_2[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27897_ (.CLK(clock),
    .D(_00926_),
    .Q(\csr._mcycle_T_2[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27898_ (.CLK(clock),
    .D(_00927_),
    .Q(\csr._mcycle_T_2[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27899_ (.CLK(clock),
    .D(_00928_),
    .Q(\csr._mcycle_T_2[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27900_ (.CLK(clock),
    .D(_00929_),
    .Q(\csr._mcycle_T_2[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27901_ (.CLK(clock),
    .D(_00930_),
    .Q(\csr._mcycle_T_2[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27902_ (.CLK(clock),
    .D(_00931_),
    .Q(\csr._mcycle_T_2[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27903_ (.CLK(clock),
    .D(_00932_),
    .Q(\csr._mcycle_T_2[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27904_ (.CLK(clock),
    .D(_00933_),
    .Q(\csr._mcycle_T_2[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27905_ (.CLK(clock),
    .D(_00934_),
    .Q(\csr._mcycle_T_2[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27906_ (.CLK(clock),
    .D(_00935_),
    .Q(\csr._mcycle_T_2[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27907_ (.CLK(clock),
    .D(_00936_),
    .Q(\csr._mcycle_T_2[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27908_ (.CLK(clock),
    .D(_00937_),
    .Q(\csr._mcycle_T_2[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27909_ (.CLK(clock),
    .D(_00938_),
    .Q(\csr._mcycle_T_2[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27910_ (.CLK(clock),
    .D(_00939_),
    .Q(\csr._mcycle_T_2[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27911_ (.CLK(clock),
    .D(_00940_),
    .Q(\csr.io_csr_write_address[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27912_ (.CLK(clock),
    .D(_00941_),
    .Q(\csr.io_csr_write_address[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27913_ (.CLK(clock),
    .D(_00942_),
    .Q(\csr.io_csr_write_address[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27914_ (.CLK(clock),
    .D(_00943_),
    .Q(\csr.io_csr_write_address[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27915_ (.CLK(clock),
    .D(_00944_),
    .Q(\csr.io_csr_write_address[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27916_ (.CLK(clock),
    .D(_00945_),
    .Q(\csr.io_csr_write_address[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27917_ (.CLK(clock),
    .D(_00946_),
    .Q(\csr.io_csr_write_address[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27918_ (.CLK(clock),
    .D(_00947_),
    .Q(\csr.io_csr_write_address[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27919_ (.CLK(clock),
    .D(_00948_),
    .Q(\csr.io_csr_write_address[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27920_ (.CLK(clock),
    .D(_00949_),
    .Q(\csr.io_csr_write_address[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27921_ (.CLK(clock),
    .D(_00950_),
    .Q(\csr.io_csr_write_address[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27922_ (.CLK(clock),
    .D(_00951_),
    .Q(\csr.io_csr_write_address[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27923_ (.CLK(clock),
    .D(_00952_),
    .Q(\csr.io_csr_write_enable ));
 sky130_fd_sc_hd__dfxtp_2 _27924_ (.CLK(clock),
    .D(_00953_),
    .Q(\execute.io_mem_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27925_ (.CLK(clock),
    .D(_00954_),
    .Q(\execute.io_mem_rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27926_ (.CLK(clock),
    .D(_00955_),
    .Q(\execute.io_mem_rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27927_ (.CLK(clock),
    .D(_00956_),
    .Q(\execute.io_mem_rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27928_ (.CLK(clock),
    .D(_00957_),
    .Q(\execute.io_mem_rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27929_ (.CLK(clock),
    .D(_00010_),
    .Q(\fetch.bht.bhtTable_valid[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27930_ (.CLK(clock),
    .D(_00009_),
    .Q(\fetch.bht.bhtTable_valid[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27931_ (.CLK(clock),
    .D(_00008_),
    .Q(\fetch.bht.bhtTable_valid[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27932_ (.CLK(clock),
    .D(_00007_),
    .Q(\fetch.bht.bhtTable_valid[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27933_ (.CLK(clock),
    .D(_00006_),
    .Q(\fetch.bht.bhtTable_valid[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27934_ (.CLK(clock),
    .D(_00005_),
    .Q(\fetch.bht.bhtTable_valid[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27935_ (.CLK(clock),
    .D(_00019_),
    .Q(\fetch.bht.bhtTable_valid[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27936_ (.CLK(clock),
    .D(_00958_),
    .Q(\fetch.bht.bhtTable_tag[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27937_ (.CLK(clock),
    .D(_00959_),
    .Q(\fetch.bht.bhtTable_tag[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27938_ (.CLK(clock),
    .D(_00960_),
    .Q(\fetch.bht.bhtTable_tag[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27939_ (.CLK(clock),
    .D(_00961_),
    .Q(\fetch.bht.bhtTable_tag[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27940_ (.CLK(clock),
    .D(_00962_),
    .Q(\fetch.bht.bhtTable_tag[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27941_ (.CLK(clock),
    .D(_00963_),
    .Q(\fetch.bht.bhtTable_tag[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27942_ (.CLK(clock),
    .D(_00964_),
    .Q(\fetch.bht.bhtTable_tag[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27943_ (.CLK(clock),
    .D(_00965_),
    .Q(\fetch.bht.bhtTable_tag[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27944_ (.CLK(clock),
    .D(_00966_),
    .Q(\fetch.bht.bhtTable_tag[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27945_ (.CLK(clock),
    .D(_00967_),
    .Q(\fetch.bht.bhtTable_tag[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27946_ (.CLK(clock),
    .D(_00968_),
    .Q(\fetch.bht.bhtTable_tag[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27947_ (.CLK(clock),
    .D(_00969_),
    .Q(\fetch.bht.bhtTable_tag[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27948_ (.CLK(clock),
    .D(_00970_),
    .Q(\fetch.bht.bhtTable_tag[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27949_ (.CLK(clock),
    .D(_00971_),
    .Q(\fetch.bht.bhtTable_tag[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27950_ (.CLK(clock),
    .D(_00972_),
    .Q(\fetch.bht.bhtTable_tag[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27951_ (.CLK(clock),
    .D(_00973_),
    .Q(\fetch.bht.bhtTable_tag[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27952_ (.CLK(clock),
    .D(_00974_),
    .Q(\fetch.bht.bhtTable_tag[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27953_ (.CLK(clock),
    .D(_00975_),
    .Q(\fetch.bht.bhtTable_tag[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27954_ (.CLK(clock),
    .D(_00976_),
    .Q(\fetch.bht.bhtTable_tag[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27955_ (.CLK(clock),
    .D(_00977_),
    .Q(\fetch.bht.bhtTable_tag[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27956_ (.CLK(clock),
    .D(_00978_),
    .Q(\fetch.bht.bhtTable_tag[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27957_ (.CLK(clock),
    .D(_00979_),
    .Q(\fetch.bht.bhtTable_tag[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27958_ (.CLK(clock),
    .D(_00980_),
    .Q(\fetch.bht.bhtTable_tag[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27959_ (.CLK(clock),
    .D(_00981_),
    .Q(\fetch.bht.bhtTable_tag[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27960_ (.CLK(clock),
    .D(_00982_),
    .Q(\fetch.bht.bhtTable_tag[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27961_ (.CLK(clock),
    .D(_00983_),
    .Q(\fetch.bht.bhtTable_tag[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27962_ (.CLK(clock),
    .D(_00984_),
    .Q(\fetch.bht.bhtTable_tag[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27963_ (.CLK(clock),
    .D(_00985_),
    .Q(\fetch.bht.bhtTable_tag[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27964_ (.CLK(clock),
    .D(_00986_),
    .Q(\fetch.bht.bhtTable_tag[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27965_ (.CLK(clock),
    .D(_00987_),
    .Q(\fetch.bht.bhtTable_tag[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27966_ (.CLK(clock),
    .D(_00988_),
    .Q(\fetch.bht.bhtTable_tag[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27967_ (.CLK(clock),
    .D(_00989_),
    .Q(\fetch.bht.bhtTable_tag[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27968_ (.CLK(clock),
    .D(_00990_),
    .Q(\fetch.bht.bhtTable_tag[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27969_ (.CLK(clock),
    .D(_00991_),
    .Q(\fetch.bht.bhtTable_tag[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27970_ (.CLK(clock),
    .D(_00992_),
    .Q(\fetch.bht.bhtTable_tag[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27971_ (.CLK(clock),
    .D(_00993_),
    .Q(\fetch.bht.bhtTable_tag[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27972_ (.CLK(clock),
    .D(_00994_),
    .Q(\fetch.bht.bhtTable_tag[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27973_ (.CLK(clock),
    .D(_00995_),
    .Q(\fetch.bht.bhtTable_tag[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27974_ (.CLK(clock),
    .D(_00996_),
    .Q(\fetch.bht.bhtTable_tag[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27975_ (.CLK(clock),
    .D(_00997_),
    .Q(\fetch.bht.bhtTable_tag[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27976_ (.CLK(clock),
    .D(_00998_),
    .Q(\fetch.bht.bhtTable_tag[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27977_ (.CLK(clock),
    .D(_00999_),
    .Q(\fetch.bht.bhtTable_tag[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27978_ (.CLK(clock),
    .D(_01000_),
    .Q(\fetch.bht.bhtTable_tag[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27979_ (.CLK(clock),
    .D(_01001_),
    .Q(\fetch.bht.bhtTable_tag[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27980_ (.CLK(clock),
    .D(_01002_),
    .Q(\fetch.bht.bhtTable_tag[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27981_ (.CLK(clock),
    .D(_01003_),
    .Q(\fetch.bht.bhtTable_tag[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27982_ (.CLK(clock),
    .D(_01004_),
    .Q(\fetch.bht.bhtTable_tag[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27983_ (.CLK(clock),
    .D(_01005_),
    .Q(\fetch.bht.bhtTable_tag[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27984_ (.CLK(clock),
    .D(_01006_),
    .Q(\fetch.bht.bhtTable_tag[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27985_ (.CLK(clock),
    .D(_01007_),
    .Q(\fetch.bht.bhtTable_tag[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27986_ (.CLK(clock),
    .D(_01008_),
    .Q(\fetch.bht.bhtTable_tag[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27987_ (.CLK(clock),
    .D(_01009_),
    .Q(\fetch.bht.bhtTable_tag[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27988_ (.CLK(clock),
    .D(_01010_),
    .Q(\fetch.bht.bhtTable_tag[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27989_ (.CLK(clock),
    .D(_01011_),
    .Q(\fetch.bht.bhtTable_tag[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27990_ (.CLK(clock),
    .D(_01012_),
    .Q(\fetch.bht.bhtTable_tag[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27991_ (.CLK(clock),
    .D(_01013_),
    .Q(\fetch.bht.bhtTable_tag[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27992_ (.CLK(clock),
    .D(_01014_),
    .Q(\fetch.bht.bhtTable_tag[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27993_ (.CLK(clock),
    .D(_01015_),
    .Q(\fetch.bht.bhtTable_tag[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27994_ (.CLK(clock),
    .D(_01016_),
    .Q(\fetch.bht.bhtTable_tag[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27995_ (.CLK(clock),
    .D(_01017_),
    .Q(\fetch.bht.bhtTable_tag[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27996_ (.CLK(clock),
    .D(_01018_),
    .Q(\fetch.bht.bhtTable_tag[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27997_ (.CLK(clock),
    .D(_01019_),
    .Q(\fetch.bht.bhtTable_tag[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27998_ (.CLK(clock),
    .D(_01020_),
    .Q(\fetch.bht.bhtTable_tag[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27999_ (.CLK(clock),
    .D(_01021_),
    .Q(\fetch.bht.bhtTable_tag[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28000_ (.CLK(clock),
    .D(_01022_),
    .Q(\fetch.bht.bhtTable_tag[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28001_ (.CLK(clock),
    .D(_01023_),
    .Q(\fetch.bht.bhtTable_tag[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28002_ (.CLK(clock),
    .D(_01024_),
    .Q(\fetch.bht.bhtTable_tag[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28003_ (.CLK(clock),
    .D(_01025_),
    .Q(\fetch.bht.bhtTable_tag[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28004_ (.CLK(clock),
    .D(_01026_),
    .Q(\fetch.bht.bhtTable_tag[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28005_ (.CLK(clock),
    .D(_01027_),
    .Q(\fetch.bht.bhtTable_tag[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28006_ (.CLK(clock),
    .D(_01028_),
    .Q(\fetch.bht.bhtTable_tag[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28007_ (.CLK(clock),
    .D(_01029_),
    .Q(\fetch.bht.bhtTable_tag[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28008_ (.CLK(clock),
    .D(_01030_),
    .Q(\fetch.bht.bhtTable_tag[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28009_ (.CLK(clock),
    .D(_01031_),
    .Q(\fetch.bht.bhtTable_tag[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28010_ (.CLK(clock),
    .D(_01032_),
    .Q(\fetch.bht.bhtTable_tag[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28011_ (.CLK(clock),
    .D(_01033_),
    .Q(\fetch.bht.bhtTable_tag[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28012_ (.CLK(clock),
    .D(_01034_),
    .Q(\fetch.bht.bhtTable_tag[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28013_ (.CLK(clock),
    .D(_01035_),
    .Q(\fetch.bht.bhtTable_tag[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28014_ (.CLK(clock),
    .D(_01036_),
    .Q(\fetch.bht.bhtTable_tag[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28015_ (.CLK(clock),
    .D(_01037_),
    .Q(\fetch.bht.bhtTable_tag[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28016_ (.CLK(clock),
    .D(_01038_),
    .Q(\fetch.bht.bhtTable_tag[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28017_ (.CLK(clock),
    .D(_01039_),
    .Q(\fetch.bht.bhtTable_tag[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28018_ (.CLK(clock),
    .D(_01040_),
    .Q(\fetch.bht.bhtTable_tag[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28019_ (.CLK(clock),
    .D(_01041_),
    .Q(\fetch.bht.bhtTable_tag[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28020_ (.CLK(clock),
    .D(_01042_),
    .Q(\fetch.bht.bhtTable_tag[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28021_ (.CLK(clock),
    .D(_01043_),
    .Q(\fetch.bht.bhtTable_tag[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28022_ (.CLK(clock),
    .D(_01044_),
    .Q(\fetch.bht.bhtTable_tag[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28023_ (.CLK(clock),
    .D(_01045_),
    .Q(\fetch.bht.bhtTable_tag[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28024_ (.CLK(clock),
    .D(_01046_),
    .Q(\fetch.bht.bhtTable_tag[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28025_ (.CLK(clock),
    .D(_01047_),
    .Q(\fetch.bht.bhtTable_tag[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28026_ (.CLK(clock),
    .D(_01048_),
    .Q(\fetch.bht.bhtTable_tag[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28027_ (.CLK(clock),
    .D(_01049_),
    .Q(\fetch.bht.bhtTable_tag[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28028_ (.CLK(clock),
    .D(_01050_),
    .Q(\fetch.bht.bhtTable_tag[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28029_ (.CLK(clock),
    .D(_01051_),
    .Q(\fetch.bht.bhtTable_tag[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28030_ (.CLK(clock),
    .D(_01052_),
    .Q(\fetch.bht.bhtTable_tag[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28031_ (.CLK(clock),
    .D(_01053_),
    .Q(\fetch.bht.bhtTable_tag[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28032_ (.CLK(clock),
    .D(_01054_),
    .Q(\fetch.bht.bhtTable_tag[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28033_ (.CLK(clock),
    .D(_01055_),
    .Q(\fetch.bht.bhtTable_tag[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28034_ (.CLK(clock),
    .D(_01056_),
    .Q(\fetch.bht.bhtTable_tag[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28035_ (.CLK(clock),
    .D(_01057_),
    .Q(\fetch.bht.bhtTable_tag[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28036_ (.CLK(clock),
    .D(_01058_),
    .Q(\fetch.bht.bhtTable_tag[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28037_ (.CLK(clock),
    .D(_01059_),
    .Q(\fetch.bht.bhtTable_tag[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28038_ (.CLK(clock),
    .D(_01060_),
    .Q(\fetch.bht.bhtTable_tag[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28039_ (.CLK(clock),
    .D(_01061_),
    .Q(\fetch.bht.bhtTable_tag[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28040_ (.CLK(clock),
    .D(_01062_),
    .Q(\decode.control.io_opcode[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28041_ (.CLK(clock),
    .D(_01063_),
    .Q(\decode.control.io_opcode[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28042_ (.CLK(clock),
    .D(_01064_),
    .Q(\decode.control.io_opcode[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28043_ (.CLK(clock),
    .D(_01065_),
    .Q(\fetch.bht.bhtTable_tag[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28044_ (.CLK(clock),
    .D(_01066_),
    .Q(\fetch.bht.bhtTable_tag[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28045_ (.CLK(clock),
    .D(_01067_),
    .Q(\fetch.bht.bhtTable_tag[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28046_ (.CLK(clock),
    .D(_01068_),
    .Q(\fetch.bht.bhtTable_tag[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28047_ (.CLK(clock),
    .D(_01069_),
    .Q(\fetch.bht.bhtTable_tag[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28048_ (.CLK(clock),
    .D(_01070_),
    .Q(\fetch.bht.bhtTable_tag[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28049_ (.CLK(clock),
    .D(_01071_),
    .Q(\fetch.bht.bhtTable_tag[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28050_ (.CLK(clock),
    .D(_01072_),
    .Q(\fetch.bht.bhtTable_tag[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28051_ (.CLK(clock),
    .D(_01073_),
    .Q(\fetch.bht.bhtTable_tag[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28052_ (.CLK(clock),
    .D(_01074_),
    .Q(\fetch.bht.bhtTable_tag[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28053_ (.CLK(clock),
    .D(_01075_),
    .Q(\fetch.bht.bhtTable_tag[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28054_ (.CLK(clock),
    .D(_01076_),
    .Q(\fetch.bht.bhtTable_tag[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28055_ (.CLK(clock),
    .D(_01077_),
    .Q(\fetch.bht.bhtTable_tag[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28056_ (.CLK(clock),
    .D(_01078_),
    .Q(\fetch.bht.bhtTable_tag[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28057_ (.CLK(clock),
    .D(_01079_),
    .Q(\fetch.bht.bhtTable_tag[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28058_ (.CLK(clock),
    .D(_01080_),
    .Q(\fetch.bht.bhtTable_tag[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28059_ (.CLK(clock),
    .D(_01081_),
    .Q(\fetch.bht.bhtTable_tag[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28060_ (.CLK(clock),
    .D(_01082_),
    .Q(\fetch.bht.bhtTable_tag[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28061_ (.CLK(clock),
    .D(_01083_),
    .Q(\fetch.bht.bhtTable_tag[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28062_ (.CLK(clock),
    .D(_01084_),
    .Q(\fetch.bht.bhtTable_tag[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28063_ (.CLK(clock),
    .D(_01085_),
    .Q(\fetch.bht.bhtTable_tag[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28064_ (.CLK(clock),
    .D(_01086_),
    .Q(\fetch.bht.bhtTable_tag[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28065_ (.CLK(clock),
    .D(_01087_),
    .Q(\fetch.bht.bhtTable_tag[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28066_ (.CLK(clock),
    .D(_01088_),
    .Q(\fetch.bht.bhtTable_tag[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28067_ (.CLK(clock),
    .D(_01089_),
    .Q(\fetch.bht.bhtTable_tag[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28068_ (.CLK(clock),
    .D(_01090_),
    .Q(\fetch.bht.bhtTable_tag[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28069_ (.CLK(clock),
    .D(_01091_),
    .Q(\fetch.bht.bhtTable_tag[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28070_ (.CLK(clock),
    .D(_01092_),
    .Q(\fetch.bht.bhtTable_tag[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28071_ (.CLK(clock),
    .D(_01093_),
    .Q(\fetch.bht.bhtTable_tag[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28072_ (.CLK(clock),
    .D(_01094_),
    .Q(\fetch.bht.bhtTable_tag[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28073_ (.CLK(clock),
    .D(_01095_),
    .Q(\fetch.bht.bhtTable_tag[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28074_ (.CLK(clock),
    .D(_01096_),
    .Q(\fetch.bht.bhtTable_tag[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28075_ (.CLK(clock),
    .D(_01097_),
    .Q(\fetch.bht.bhtTable_tag[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28076_ (.CLK(clock),
    .D(_01098_),
    .Q(\fetch.bht.bhtTable_tag[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28077_ (.CLK(clock),
    .D(_01099_),
    .Q(\fetch.bht.bhtTable_tag[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28078_ (.CLK(clock),
    .D(_01100_),
    .Q(\fetch.bht.bhtTable_tag[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28079_ (.CLK(clock),
    .D(_01101_),
    .Q(\fetch.bht.bhtTable_tag[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28080_ (.CLK(clock),
    .D(_01102_),
    .Q(\fetch.bht.bhtTable_tag[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28081_ (.CLK(clock),
    .D(_01103_),
    .Q(\fetch.bht.bhtTable_tag[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28082_ (.CLK(clock),
    .D(_01104_),
    .Q(\fetch.bht.bhtTable_tag[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28083_ (.CLK(clock),
    .D(_01105_),
    .Q(\fetch.bht.bhtTable_tag[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28084_ (.CLK(clock),
    .D(_01106_),
    .Q(\fetch.bht.bhtTable_tag[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28085_ (.CLK(clock),
    .D(_01107_),
    .Q(\fetch.bht.bhtTable_tag[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28086_ (.CLK(clock),
    .D(_01108_),
    .Q(\fetch.bht.bhtTable_tag[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28087_ (.CLK(clock),
    .D(_01109_),
    .Q(\fetch.bht.bhtTable_tag[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28088_ (.CLK(clock),
    .D(_01110_),
    .Q(\fetch.bht.bhtTable_tag[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28089_ (.CLK(clock),
    .D(_01111_),
    .Q(\fetch.bht.bhtTable_tag[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28090_ (.CLK(clock),
    .D(_01112_),
    .Q(\fetch.bht.bhtTable_tag[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28091_ (.CLK(clock),
    .D(_01113_),
    .Q(\fetch.bht.bhtTable_tag[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28092_ (.CLK(clock),
    .D(_01114_),
    .Q(\fetch.bht.bhtTable_tag[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28093_ (.CLK(clock),
    .D(_01115_),
    .Q(\fetch.bht.bhtTable_tag[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28094_ (.CLK(clock),
    .D(_01116_),
    .Q(\fetch.bht.bhtTable_tag[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28095_ (.CLK(clock),
    .D(_01117_),
    .Q(\csr.minstret[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28096_ (.CLK(clock),
    .D(_01118_),
    .Q(\csr.minstret[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28097_ (.CLK(clock),
    .D(_01119_),
    .Q(\csr.minstret[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28098_ (.CLK(clock),
    .D(_01120_),
    .Q(\csr.minstret[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28099_ (.CLK(clock),
    .D(_01121_),
    .Q(\csr.minstret[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28100_ (.CLK(clock),
    .D(_01122_),
    .Q(\csr.minstret[5] ));
 sky130_fd_sc_hd__dfxtp_2 _28101_ (.CLK(clock),
    .D(_01123_),
    .Q(\csr.minstret[6] ));
 sky130_fd_sc_hd__dfxtp_2 _28102_ (.CLK(clock),
    .D(_01124_),
    .Q(\csr.minstret[7] ));
 sky130_fd_sc_hd__dfxtp_2 _28103_ (.CLK(clock),
    .D(_01125_),
    .Q(\csr.minstret[8] ));
 sky130_fd_sc_hd__dfxtp_2 _28104_ (.CLK(clock),
    .D(_01126_),
    .Q(\csr.minstret[9] ));
 sky130_fd_sc_hd__dfxtp_2 _28105_ (.CLK(clock),
    .D(_01127_),
    .Q(\csr.minstret[10] ));
 sky130_fd_sc_hd__dfxtp_2 _28106_ (.CLK(clock),
    .D(_01128_),
    .Q(\csr.minstret[11] ));
 sky130_fd_sc_hd__dfxtp_2 _28107_ (.CLK(clock),
    .D(_01129_),
    .Q(\csr.minstret[12] ));
 sky130_fd_sc_hd__dfxtp_2 _28108_ (.CLK(clock),
    .D(_01130_),
    .Q(\csr.minstret[13] ));
 sky130_fd_sc_hd__dfxtp_2 _28109_ (.CLK(clock),
    .D(_01131_),
    .Q(\csr.minstret[14] ));
 sky130_fd_sc_hd__dfxtp_2 _28110_ (.CLK(clock),
    .D(_01132_),
    .Q(\csr.minstret[15] ));
 sky130_fd_sc_hd__dfxtp_2 _28111_ (.CLK(clock),
    .D(_01133_),
    .Q(\csr.minstret[16] ));
 sky130_fd_sc_hd__dfxtp_2 _28112_ (.CLK(clock),
    .D(_01134_),
    .Q(\csr.minstret[17] ));
 sky130_fd_sc_hd__dfxtp_2 _28113_ (.CLK(clock),
    .D(_01135_),
    .Q(\csr.minstret[18] ));
 sky130_fd_sc_hd__dfxtp_2 _28114_ (.CLK(clock),
    .D(_01136_),
    .Q(\csr.minstret[19] ));
 sky130_fd_sc_hd__dfxtp_2 _28115_ (.CLK(clock),
    .D(_01137_),
    .Q(\csr.minstret[20] ));
 sky130_fd_sc_hd__dfxtp_2 _28116_ (.CLK(clock),
    .D(_01138_),
    .Q(\csr.minstret[21] ));
 sky130_fd_sc_hd__dfxtp_2 _28117_ (.CLK(clock),
    .D(_01139_),
    .Q(\csr.minstret[22] ));
 sky130_fd_sc_hd__dfxtp_2 _28118_ (.CLK(clock),
    .D(_01140_),
    .Q(\csr.minstret[23] ));
 sky130_fd_sc_hd__dfxtp_2 _28119_ (.CLK(clock),
    .D(_01141_),
    .Q(\csr.minstret[24] ));
 sky130_fd_sc_hd__dfxtp_2 _28120_ (.CLK(clock),
    .D(_01142_),
    .Q(\csr.minstret[25] ));
 sky130_fd_sc_hd__dfxtp_2 _28121_ (.CLK(clock),
    .D(_01143_),
    .Q(\csr.minstret[26] ));
 sky130_fd_sc_hd__dfxtp_2 _28122_ (.CLK(clock),
    .D(_01144_),
    .Q(\csr.minstret[27] ));
 sky130_fd_sc_hd__dfxtp_2 _28123_ (.CLK(clock),
    .D(_01145_),
    .Q(\csr.minstret[28] ));
 sky130_fd_sc_hd__dfxtp_2 _28124_ (.CLK(clock),
    .D(_01146_),
    .Q(\csr.minstret[29] ));
 sky130_fd_sc_hd__dfxtp_2 _28125_ (.CLK(clock),
    .D(_01147_),
    .Q(\csr.minstret[30] ));
 sky130_fd_sc_hd__dfxtp_2 _28126_ (.CLK(clock),
    .D(_01148_),
    .Q(\csr.minstret[31] ));
 sky130_fd_sc_hd__dfxtp_2 _28127_ (.CLK(clock),
    .D(_01149_),
    .Q(\csr.io_ecause[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28128_ (.CLK(clock),
    .D(_01150_),
    .Q(\fetch.bht.bhtTable_tag[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28129_ (.CLK(clock),
    .D(_01151_),
    .Q(\fetch.bht.bhtTable_tag[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28130_ (.CLK(clock),
    .D(_01152_),
    .Q(\fetch.bht.bhtTable_tag[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28131_ (.CLK(clock),
    .D(_01153_),
    .Q(\fetch.bht.bhtTable_tag[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28132_ (.CLK(clock),
    .D(_01154_),
    .Q(\fetch.bht.bhtTable_tag[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28133_ (.CLK(clock),
    .D(_01155_),
    .Q(\fetch.bht.bhtTable_tag[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28134_ (.CLK(clock),
    .D(_01156_),
    .Q(\fetch.bht.bhtTable_tag[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28135_ (.CLK(clock),
    .D(_01157_),
    .Q(\fetch.bht.bhtTable_tag[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28136_ (.CLK(clock),
    .D(_01158_),
    .Q(\fetch.bht.bhtTable_tag[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28137_ (.CLK(clock),
    .D(_01159_),
    .Q(\fetch.bht.bhtTable_tag[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28138_ (.CLK(clock),
    .D(_01160_),
    .Q(\fetch.bht.bhtTable_tag[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28139_ (.CLK(clock),
    .D(_01161_),
    .Q(\fetch.bht.bhtTable_tag[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28140_ (.CLK(clock),
    .D(_01162_),
    .Q(\fetch.bht.bhtTable_tag[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28141_ (.CLK(clock),
    .D(_01163_),
    .Q(\fetch.bht.bhtTable_tag[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28142_ (.CLK(clock),
    .D(_01164_),
    .Q(\fetch.bht.bhtTable_tag[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28143_ (.CLK(clock),
    .D(_01165_),
    .Q(\fetch.bht.bhtTable_tag[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28144_ (.CLK(clock),
    .D(_01166_),
    .Q(\fetch.bht.bhtTable_tag[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28145_ (.CLK(clock),
    .D(_01167_),
    .Q(\fetch.bht.bhtTable_tag[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28146_ (.CLK(clock),
    .D(_01168_),
    .Q(\fetch.bht.bhtTable_tag[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28147_ (.CLK(clock),
    .D(_01169_),
    .Q(\fetch.bht.bhtTable_tag[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28148_ (.CLK(clock),
    .D(_01170_),
    .Q(\fetch.bht.bhtTable_tag[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28149_ (.CLK(clock),
    .D(_01171_),
    .Q(\fetch.bht.bhtTable_tag[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28150_ (.CLK(clock),
    .D(_01172_),
    .Q(\fetch.bht.bhtTable_tag[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28151_ (.CLK(clock),
    .D(_01173_),
    .Q(\fetch.bht.bhtTable_tag[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28152_ (.CLK(clock),
    .D(_01174_),
    .Q(\fetch.bht.bhtTable_tag[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28153_ (.CLK(clock),
    .D(_01175_),
    .Q(\fetch.bht.bhtTable_tag[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28154_ (.CLK(clock),
    .D(_01176_),
    .Q(\fetch.btb.io_branch ));
 sky130_fd_sc_hd__dfxtp_2 _28155_ (.CLK(clock),
    .D(_01177_),
    .Q(\csr.ie ));
 sky130_fd_sc_hd__dfxtp_2 _28156_ (.CLK(clock),
    .D(_01178_),
    .Q(\csr.mtie ));
 sky130_fd_sc_hd__dfxtp_2 _28157_ (.CLK(clock),
    .D(_01179_),
    .Q(\csr.msip ));
 sky130_fd_sc_hd__dfxtp_2 _28158_ (.CLK(clock),
    .D(_01180_),
    .Q(\csr.msie ));
 sky130_fd_sc_hd__dfxtp_2 _28159_ (.CLK(clock),
    .D(_01181_),
    .Q(\csr.meie ));
 sky130_fd_sc_hd__dfxtp_2 _28160_ (.CLK(clock),
    .D(_01182_),
    .Q(\csr.pie ));
 sky130_fd_sc_hd__dfxtp_2 _28161_ (.CLK(clock),
    .D(_01183_),
    .Q(\csr._csr_read_data_T_9[31] ));
 sky130_fd_sc_hd__dfxtp_2 _28162_ (.CLK(clock),
    .D(_01184_),
    .Q(\csr._csr_read_data_T_9[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28163_ (.CLK(clock),
    .D(_01185_),
    .Q(\csr._csr_read_data_T_9[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28164_ (.CLK(clock),
    .D(_01186_),
    .Q(\csr._csr_read_data_T_9[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28165_ (.CLK(clock),
    .D(_01187_),
    .Q(\csr._csr_read_data_T_9[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28166_ (.CLK(clock),
    .D(_01188_),
    .Q(\csr.io_mret_vector[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28167_ (.CLK(clock),
    .D(_01189_),
    .Q(\csr.io_mret_vector[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28168_ (.CLK(clock),
    .D(_01190_),
    .Q(\csr.io_mret_vector[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28169_ (.CLK(clock),
    .D(_01191_),
    .Q(\csr.io_mret_vector[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28170_ (.CLK(clock),
    .D(_01192_),
    .Q(\csr.io_mret_vector[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28171_ (.CLK(clock),
    .D(_01193_),
    .Q(\csr.io_mret_vector[5] ));
 sky130_fd_sc_hd__dfxtp_2 _28172_ (.CLK(clock),
    .D(_01194_),
    .Q(\csr.io_mret_vector[6] ));
 sky130_fd_sc_hd__dfxtp_2 _28173_ (.CLK(clock),
    .D(_01195_),
    .Q(\csr.io_mret_vector[7] ));
 sky130_fd_sc_hd__dfxtp_2 _28174_ (.CLK(clock),
    .D(_01196_),
    .Q(\csr.io_mret_vector[8] ));
 sky130_fd_sc_hd__dfxtp_2 _28175_ (.CLK(clock),
    .D(_01197_),
    .Q(\csr.io_mret_vector[9] ));
 sky130_fd_sc_hd__dfxtp_2 _28176_ (.CLK(clock),
    .D(_01198_),
    .Q(\csr.io_mret_vector[10] ));
 sky130_fd_sc_hd__dfxtp_2 _28177_ (.CLK(clock),
    .D(_01199_),
    .Q(\csr.io_mret_vector[11] ));
 sky130_fd_sc_hd__dfxtp_2 _28178_ (.CLK(clock),
    .D(_01200_),
    .Q(\csr.io_mret_vector[12] ));
 sky130_fd_sc_hd__dfxtp_2 _28179_ (.CLK(clock),
    .D(_01201_),
    .Q(\csr.io_mret_vector[13] ));
 sky130_fd_sc_hd__dfxtp_2 _28180_ (.CLK(clock),
    .D(_01202_),
    .Q(\csr.io_mret_vector[14] ));
 sky130_fd_sc_hd__dfxtp_2 _28181_ (.CLK(clock),
    .D(_01203_),
    .Q(\csr.io_mret_vector[15] ));
 sky130_fd_sc_hd__dfxtp_2 _28182_ (.CLK(clock),
    .D(_01204_),
    .Q(\csr.io_mret_vector[16] ));
 sky130_fd_sc_hd__dfxtp_2 _28183_ (.CLK(clock),
    .D(_01205_),
    .Q(\csr.io_mret_vector[17] ));
 sky130_fd_sc_hd__dfxtp_2 _28184_ (.CLK(clock),
    .D(_01206_),
    .Q(\csr.io_mret_vector[18] ));
 sky130_fd_sc_hd__dfxtp_2 _28185_ (.CLK(clock),
    .D(_01207_),
    .Q(\csr.io_mret_vector[19] ));
 sky130_fd_sc_hd__dfxtp_2 _28186_ (.CLK(clock),
    .D(_01208_),
    .Q(\csr.io_mret_vector[20] ));
 sky130_fd_sc_hd__dfxtp_2 _28187_ (.CLK(clock),
    .D(_01209_),
    .Q(\csr.io_mret_vector[21] ));
 sky130_fd_sc_hd__dfxtp_2 _28188_ (.CLK(clock),
    .D(_01210_),
    .Q(\csr.io_mret_vector[22] ));
 sky130_fd_sc_hd__dfxtp_2 _28189_ (.CLK(clock),
    .D(_01211_),
    .Q(\csr.io_mret_vector[23] ));
 sky130_fd_sc_hd__dfxtp_2 _28190_ (.CLK(clock),
    .D(_01212_),
    .Q(\csr.io_mret_vector[24] ));
 sky130_fd_sc_hd__dfxtp_2 _28191_ (.CLK(clock),
    .D(_01213_),
    .Q(\csr.io_mret_vector[25] ));
 sky130_fd_sc_hd__dfxtp_2 _28192_ (.CLK(clock),
    .D(_01214_),
    .Q(\csr.io_mret_vector[26] ));
 sky130_fd_sc_hd__dfxtp_2 _28193_ (.CLK(clock),
    .D(_01215_),
    .Q(\csr.io_mret_vector[27] ));
 sky130_fd_sc_hd__dfxtp_2 _28194_ (.CLK(clock),
    .D(_01216_),
    .Q(\csr.io_mret_vector[28] ));
 sky130_fd_sc_hd__dfxtp_2 _28195_ (.CLK(clock),
    .D(_01217_),
    .Q(\csr.io_mret_vector[29] ));
 sky130_fd_sc_hd__dfxtp_2 _28196_ (.CLK(clock),
    .D(_01218_),
    .Q(\csr.io_mret_vector[30] ));
 sky130_fd_sc_hd__dfxtp_2 _28197_ (.CLK(clock),
    .D(_01219_),
    .Q(\csr.io_mret_vector[31] ));
 sky130_fd_sc_hd__dfxtp_2 _28198_ (.CLK(clock),
    .D(_01220_),
    .Q(\csr.mscratch[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28199_ (.CLK(clock),
    .D(_01221_),
    .Q(\csr.mscratch[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28200_ (.CLK(clock),
    .D(_01222_),
    .Q(\csr.mscratch[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28201_ (.CLK(clock),
    .D(_01223_),
    .Q(\csr.mscratch[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28202_ (.CLK(clock),
    .D(_01224_),
    .Q(\csr.mscratch[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28203_ (.CLK(clock),
    .D(_01225_),
    .Q(\csr.mscratch[5] ));
 sky130_fd_sc_hd__dfxtp_2 _28204_ (.CLK(clock),
    .D(_01226_),
    .Q(\csr.mscratch[6] ));
 sky130_fd_sc_hd__dfxtp_2 _28205_ (.CLK(clock),
    .D(_01227_),
    .Q(\csr.mscratch[7] ));
 sky130_fd_sc_hd__dfxtp_2 _28206_ (.CLK(clock),
    .D(_01228_),
    .Q(\csr.mscratch[8] ));
 sky130_fd_sc_hd__dfxtp_2 _28207_ (.CLK(clock),
    .D(_01229_),
    .Q(\csr.mscratch[9] ));
 sky130_fd_sc_hd__dfxtp_2 _28208_ (.CLK(clock),
    .D(_01230_),
    .Q(\csr.mscratch[10] ));
 sky130_fd_sc_hd__dfxtp_2 _28209_ (.CLK(clock),
    .D(_01231_),
    .Q(\csr.mscratch[11] ));
 sky130_fd_sc_hd__dfxtp_2 _28210_ (.CLK(clock),
    .D(_01232_),
    .Q(\csr.mscratch[12] ));
 sky130_fd_sc_hd__dfxtp_2 _28211_ (.CLK(clock),
    .D(_01233_),
    .Q(\csr.mscratch[13] ));
 sky130_fd_sc_hd__dfxtp_2 _28212_ (.CLK(clock),
    .D(_01234_),
    .Q(\csr.mscratch[14] ));
 sky130_fd_sc_hd__dfxtp_2 _28213_ (.CLK(clock),
    .D(_01235_),
    .Q(\csr.mscratch[15] ));
 sky130_fd_sc_hd__dfxtp_2 _28214_ (.CLK(clock),
    .D(_01236_),
    .Q(\csr.mscratch[16] ));
 sky130_fd_sc_hd__dfxtp_2 _28215_ (.CLK(clock),
    .D(_01237_),
    .Q(\csr.mscratch[17] ));
 sky130_fd_sc_hd__dfxtp_2 _28216_ (.CLK(clock),
    .D(_01238_),
    .Q(\csr.mscratch[18] ));
 sky130_fd_sc_hd__dfxtp_2 _28217_ (.CLK(clock),
    .D(_01239_),
    .Q(\csr.mscratch[19] ));
 sky130_fd_sc_hd__dfxtp_2 _28218_ (.CLK(clock),
    .D(_01240_),
    .Q(\csr.mscratch[20] ));
 sky130_fd_sc_hd__dfxtp_2 _28219_ (.CLK(clock),
    .D(_01241_),
    .Q(\csr.mscratch[21] ));
 sky130_fd_sc_hd__dfxtp_2 _28220_ (.CLK(clock),
    .D(_01242_),
    .Q(\csr.mscratch[22] ));
 sky130_fd_sc_hd__dfxtp_2 _28221_ (.CLK(clock),
    .D(_01243_),
    .Q(\csr.mscratch[23] ));
 sky130_fd_sc_hd__dfxtp_2 _28222_ (.CLK(clock),
    .D(_01244_),
    .Q(\csr.mscratch[24] ));
 sky130_fd_sc_hd__dfxtp_2 _28223_ (.CLK(clock),
    .D(_01245_),
    .Q(\csr.mscratch[25] ));
 sky130_fd_sc_hd__dfxtp_2 _28224_ (.CLK(clock),
    .D(_01246_),
    .Q(\csr.mscratch[26] ));
 sky130_fd_sc_hd__dfxtp_2 _28225_ (.CLK(clock),
    .D(_01247_),
    .Q(\csr.mscratch[27] ));
 sky130_fd_sc_hd__dfxtp_2 _28226_ (.CLK(clock),
    .D(_01248_),
    .Q(\csr.mscratch[28] ));
 sky130_fd_sc_hd__dfxtp_2 _28227_ (.CLK(clock),
    .D(_01249_),
    .Q(\csr.mscratch[29] ));
 sky130_fd_sc_hd__dfxtp_2 _28228_ (.CLK(clock),
    .D(_01250_),
    .Q(\csr.mscratch[30] ));
 sky130_fd_sc_hd__dfxtp_2 _28229_ (.CLK(clock),
    .D(_01251_),
    .Q(\csr.mscratch[31] ));
 sky130_fd_sc_hd__dfxtp_2 _28230_ (.CLK(clock),
    .D(_01252_),
    .Q(io_fetch_address[0]));
 sky130_fd_sc_hd__dfxtp_2 _28231_ (.CLK(clock),
    .D(_01253_),
    .Q(io_fetch_address[1]));
 sky130_fd_sc_hd__dfxtp_2 _28232_ (.CLK(clock),
    .D(_01254_),
    .Q(\csr._minstret_T_3[32] ));
 sky130_fd_sc_hd__dfxtp_2 _28233_ (.CLK(clock),
    .D(_01255_),
    .Q(\csr._minstret_T_3[33] ));
 sky130_fd_sc_hd__dfxtp_2 _28234_ (.CLK(clock),
    .D(_01256_),
    .Q(\csr._minstret_T_3[34] ));
 sky130_fd_sc_hd__dfxtp_2 _28235_ (.CLK(clock),
    .D(_01257_),
    .Q(\csr._minstret_T_3[35] ));
 sky130_fd_sc_hd__dfxtp_2 _28236_ (.CLK(clock),
    .D(_01258_),
    .Q(\csr._minstret_T_3[36] ));
 sky130_fd_sc_hd__dfxtp_2 _28237_ (.CLK(clock),
    .D(_01259_),
    .Q(\csr._minstret_T_3[37] ));
 sky130_fd_sc_hd__dfxtp_2 _28238_ (.CLK(clock),
    .D(_01260_),
    .Q(\csr._minstret_T_3[38] ));
 sky130_fd_sc_hd__dfxtp_2 _28239_ (.CLK(clock),
    .D(_01261_),
    .Q(\csr._minstret_T_3[39] ));
 sky130_fd_sc_hd__dfxtp_2 _28240_ (.CLK(clock),
    .D(_01262_),
    .Q(\csr._minstret_T_3[40] ));
 sky130_fd_sc_hd__dfxtp_2 _28241_ (.CLK(clock),
    .D(_01263_),
    .Q(\csr._minstret_T_3[41] ));
 sky130_fd_sc_hd__dfxtp_2 _28242_ (.CLK(clock),
    .D(_01264_),
    .Q(\csr._minstret_T_3[42] ));
 sky130_fd_sc_hd__dfxtp_2 _28243_ (.CLK(clock),
    .D(_01265_),
    .Q(\csr._minstret_T_3[43] ));
 sky130_fd_sc_hd__dfxtp_2 _28244_ (.CLK(clock),
    .D(_01266_),
    .Q(\csr._minstret_T_3[44] ));
 sky130_fd_sc_hd__dfxtp_2 _28245_ (.CLK(clock),
    .D(_01267_),
    .Q(\csr._minstret_T_3[45] ));
 sky130_fd_sc_hd__dfxtp_2 _28246_ (.CLK(clock),
    .D(_01268_),
    .Q(\csr._minstret_T_3[46] ));
 sky130_fd_sc_hd__dfxtp_2 _28247_ (.CLK(clock),
    .D(_01269_),
    .Q(\csr._minstret_T_3[47] ));
 sky130_fd_sc_hd__dfxtp_2 _28248_ (.CLK(clock),
    .D(_01270_),
    .Q(\csr._minstret_T_3[48] ));
 sky130_fd_sc_hd__dfxtp_2 _28249_ (.CLK(clock),
    .D(_01271_),
    .Q(\csr._minstret_T_3[49] ));
 sky130_fd_sc_hd__dfxtp_2 _28250_ (.CLK(clock),
    .D(_01272_),
    .Q(\csr._minstret_T_3[50] ));
 sky130_fd_sc_hd__dfxtp_2 _28251_ (.CLK(clock),
    .D(_01273_),
    .Q(\csr._minstret_T_3[51] ));
 sky130_fd_sc_hd__dfxtp_2 _28252_ (.CLK(clock),
    .D(_01274_),
    .Q(\csr._minstret_T_3[52] ));
 sky130_fd_sc_hd__dfxtp_2 _28253_ (.CLK(clock),
    .D(_01275_),
    .Q(\csr._minstret_T_3[53] ));
 sky130_fd_sc_hd__dfxtp_2 _28254_ (.CLK(clock),
    .D(_01276_),
    .Q(\csr._minstret_T_3[54] ));
 sky130_fd_sc_hd__dfxtp_2 _28255_ (.CLK(clock),
    .D(_01277_),
    .Q(\csr._minstret_T_3[55] ));
 sky130_fd_sc_hd__dfxtp_2 _28256_ (.CLK(clock),
    .D(_01278_),
    .Q(\csr._minstret_T_3[56] ));
 sky130_fd_sc_hd__dfxtp_2 _28257_ (.CLK(clock),
    .D(_01279_),
    .Q(\csr._minstret_T_3[57] ));
 sky130_fd_sc_hd__dfxtp_2 _28258_ (.CLK(clock),
    .D(_01280_),
    .Q(\csr._minstret_T_3[58] ));
 sky130_fd_sc_hd__dfxtp_2 _28259_ (.CLK(clock),
    .D(_01281_),
    .Q(\csr._minstret_T_3[59] ));
 sky130_fd_sc_hd__dfxtp_2 _28260_ (.CLK(clock),
    .D(_01282_),
    .Q(\csr._minstret_T_3[60] ));
 sky130_fd_sc_hd__dfxtp_2 _28261_ (.CLK(clock),
    .D(_01283_),
    .Q(\csr._minstret_T_3[61] ));
 sky130_fd_sc_hd__dfxtp_2 _28262_ (.CLK(clock),
    .D(_01284_),
    .Q(\csr._minstret_T_3[62] ));
 sky130_fd_sc_hd__dfxtp_2 _28263_ (.CLK(clock),
    .D(_01285_),
    .Q(\csr._minstret_T_3[63] ));
 sky130_fd_sc_hd__dfxtp_2 _28264_ (.CLK(clock),
    .D(_01286_),
    .Q(\csr._csr_read_data_T_8[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28265_ (.CLK(clock),
    .D(_01287_),
    .Q(\csr._csr_read_data_T_8[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28266_ (.CLK(clock),
    .D(_01288_),
    .Q(\csr._csr_read_data_T_8[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28267_ (.CLK(clock),
    .D(_01289_),
    .Q(\csr._csr_read_data_T_8[5] ));
 sky130_fd_sc_hd__dfxtp_2 _28268_ (.CLK(clock),
    .D(_01290_),
    .Q(\csr._csr_read_data_T_8[6] ));
 sky130_fd_sc_hd__dfxtp_2 _28269_ (.CLK(clock),
    .D(_01291_),
    .Q(\csr._csr_read_data_T_8[7] ));
 sky130_fd_sc_hd__dfxtp_2 _28270_ (.CLK(clock),
    .D(_01292_),
    .Q(\csr._csr_read_data_T_8[8] ));
 sky130_fd_sc_hd__dfxtp_2 _28271_ (.CLK(clock),
    .D(_01293_),
    .Q(\csr._csr_read_data_T_8[9] ));
 sky130_fd_sc_hd__dfxtp_2 _28272_ (.CLK(clock),
    .D(_01294_),
    .Q(\csr._csr_read_data_T_8[10] ));
 sky130_fd_sc_hd__dfxtp_2 _28273_ (.CLK(clock),
    .D(_01295_),
    .Q(\csr._csr_read_data_T_8[11] ));
 sky130_fd_sc_hd__dfxtp_2 _28274_ (.CLK(clock),
    .D(_01296_),
    .Q(\csr._csr_read_data_T_8[12] ));
 sky130_fd_sc_hd__dfxtp_2 _28275_ (.CLK(clock),
    .D(_01297_),
    .Q(\csr._csr_read_data_T_8[13] ));
 sky130_fd_sc_hd__dfxtp_2 _28276_ (.CLK(clock),
    .D(_01298_),
    .Q(\csr._csr_read_data_T_8[14] ));
 sky130_fd_sc_hd__dfxtp_2 _28277_ (.CLK(clock),
    .D(_01299_),
    .Q(\csr._csr_read_data_T_8[15] ));
 sky130_fd_sc_hd__dfxtp_2 _28278_ (.CLK(clock),
    .D(_01300_),
    .Q(\csr._csr_read_data_T_8[16] ));
 sky130_fd_sc_hd__dfxtp_2 _28279_ (.CLK(clock),
    .D(_01301_),
    .Q(\csr._csr_read_data_T_8[17] ));
 sky130_fd_sc_hd__dfxtp_2 _28280_ (.CLK(clock),
    .D(_01302_),
    .Q(\csr._csr_read_data_T_8[18] ));
 sky130_fd_sc_hd__dfxtp_2 _28281_ (.CLK(clock),
    .D(_01303_),
    .Q(\csr._csr_read_data_T_8[19] ));
 sky130_fd_sc_hd__dfxtp_2 _28282_ (.CLK(clock),
    .D(_01304_),
    .Q(\csr._csr_read_data_T_8[20] ));
 sky130_fd_sc_hd__dfxtp_2 _28283_ (.CLK(clock),
    .D(_01305_),
    .Q(\csr._csr_read_data_T_8[21] ));
 sky130_fd_sc_hd__dfxtp_2 _28284_ (.CLK(clock),
    .D(_01306_),
    .Q(\csr._csr_read_data_T_8[22] ));
 sky130_fd_sc_hd__dfxtp_2 _28285_ (.CLK(clock),
    .D(_01307_),
    .Q(\csr._csr_read_data_T_8[23] ));
 sky130_fd_sc_hd__dfxtp_2 _28286_ (.CLK(clock),
    .D(_01308_),
    .Q(\csr._csr_read_data_T_8[24] ));
 sky130_fd_sc_hd__dfxtp_2 _28287_ (.CLK(clock),
    .D(_01309_),
    .Q(\csr._csr_read_data_T_8[25] ));
 sky130_fd_sc_hd__dfxtp_2 _28288_ (.CLK(clock),
    .D(_01310_),
    .Q(\csr._csr_read_data_T_8[26] ));
 sky130_fd_sc_hd__dfxtp_2 _28289_ (.CLK(clock),
    .D(_01311_),
    .Q(\csr._csr_read_data_T_8[27] ));
 sky130_fd_sc_hd__dfxtp_2 _28290_ (.CLK(clock),
    .D(_01312_),
    .Q(\csr._csr_read_data_T_8[28] ));
 sky130_fd_sc_hd__dfxtp_2 _28291_ (.CLK(clock),
    .D(_01313_),
    .Q(\csr._csr_read_data_T_8[29] ));
 sky130_fd_sc_hd__dfxtp_2 _28292_ (.CLK(clock),
    .D(_01314_),
    .Q(\csr._csr_read_data_T_8[30] ));
 sky130_fd_sc_hd__dfxtp_2 _28293_ (.CLK(clock),
    .D(_01315_),
    .Q(\csr._csr_read_data_T_8[31] ));
 sky130_fd_sc_hd__dfxtp_2 _28294_ (.CLK(clock),
    .D(_00018_),
    .Q(\fetch.bht.bhtTable_valid[8] ));
 sky130_fd_sc_hd__dfxtp_2 _28295_ (.CLK(clock),
    .D(_00017_),
    .Q(\fetch.bht.bhtTable_valid[7] ));
 sky130_fd_sc_hd__dfxtp_2 _28296_ (.CLK(clock),
    .D(_00016_),
    .Q(\fetch.bht.bhtTable_valid[6] ));
 sky130_fd_sc_hd__dfxtp_2 _28297_ (.CLK(clock),
    .D(_00015_),
    .Q(\fetch.bht.bhtTable_valid[5] ));
 sky130_fd_sc_hd__dfxtp_2 _28298_ (.CLK(clock),
    .D(_00014_),
    .Q(\fetch.bht.bhtTable_valid[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28299_ (.CLK(clock),
    .D(_00013_),
    .Q(\fetch.bht.bhtTable_valid[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28300_ (.CLK(clock),
    .D(_00012_),
    .Q(\fetch.bht.bhtTable_valid[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28301_ (.CLK(clock),
    .D(_00011_),
    .Q(\fetch.bht.bhtTable_valid[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28302_ (.CLK(clock),
    .D(_00004_),
    .Q(\fetch.bht.bhtTable_valid[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28303_ (.CLK(clock),
    .D(_01316_),
    .Q(\decode.id_ex_aluop_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28304_ (.CLK(clock),
    .D(_01317_),
    .Q(\decode.id_ex_aluop_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28305_ (.CLK(clock),
    .D(_01318_),
    .Q(\fetch.bht.bhtTable_tag[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28306_ (.CLK(clock),
    .D(_01319_),
    .Q(\fetch.bht.bhtTable_tag[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28307_ (.CLK(clock),
    .D(_01320_),
    .Q(\fetch.bht.bhtTable_tag[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28308_ (.CLK(clock),
    .D(_01321_),
    .Q(\fetch.bht.bhtTable_tag[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28309_ (.CLK(clock),
    .D(_01322_),
    .Q(\fetch.bht.bhtTable_tag[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28310_ (.CLK(clock),
    .D(_01323_),
    .Q(\fetch.bht.bhtTable_tag[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28311_ (.CLK(clock),
    .D(_01324_),
    .Q(\fetch.bht.bhtTable_tag[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28312_ (.CLK(clock),
    .D(_01325_),
    .Q(\fetch.bht.bhtTable_tag[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28313_ (.CLK(clock),
    .D(_01326_),
    .Q(\fetch.bht.bhtTable_tag[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28314_ (.CLK(clock),
    .D(_01327_),
    .Q(\fetch.bht.bhtTable_tag[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28315_ (.CLK(clock),
    .D(_01328_),
    .Q(\fetch.bht.bhtTable_tag[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28316_ (.CLK(clock),
    .D(_01329_),
    .Q(\fetch.bht.bhtTable_tag[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28317_ (.CLK(clock),
    .D(_01330_),
    .Q(\fetch.bht.bhtTable_tag[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28318_ (.CLK(clock),
    .D(_01331_),
    .Q(\fetch.bht.bhtTable_tag[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28319_ (.CLK(clock),
    .D(_01332_),
    .Q(\fetch.bht.bhtTable_tag[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28320_ (.CLK(clock),
    .D(_01333_),
    .Q(\fetch.bht.bhtTable_tag[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28321_ (.CLK(clock),
    .D(_01334_),
    .Q(\fetch.bht.bhtTable_tag[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28322_ (.CLK(clock),
    .D(_01335_),
    .Q(\fetch.bht.bhtTable_tag[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28323_ (.CLK(clock),
    .D(_01336_),
    .Q(\fetch.bht.bhtTable_tag[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28324_ (.CLK(clock),
    .D(_01337_),
    .Q(\fetch.bht.bhtTable_tag[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28325_ (.CLK(clock),
    .D(_01338_),
    .Q(\fetch.bht.bhtTable_tag[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28326_ (.CLK(clock),
    .D(_01339_),
    .Q(\fetch.bht.bhtTable_tag[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28327_ (.CLK(clock),
    .D(_01340_),
    .Q(\fetch.bht.bhtTable_tag[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28328_ (.CLK(clock),
    .D(_01341_),
    .Q(\fetch.bht.bhtTable_tag[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28329_ (.CLK(clock),
    .D(_01342_),
    .Q(\fetch.bht.bhtTable_tag[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28330_ (.CLK(clock),
    .D(_01343_),
    .Q(\fetch.bht.bhtTable_tag[10][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28331_ (.CLK(clock),
    .D(_01344_),
    .Q(\fetch.bht.bhtTable_tag[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28332_ (.CLK(clock),
    .D(_01345_),
    .Q(\fetch.bht.bhtTable_tag[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28333_ (.CLK(clock),
    .D(_01346_),
    .Q(\fetch.bht.bhtTable_tag[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28334_ (.CLK(clock),
    .D(_01347_),
    .Q(\fetch.bht.bhtTable_tag[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28335_ (.CLK(clock),
    .D(_01348_),
    .Q(\fetch.bht.bhtTable_tag[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28336_ (.CLK(clock),
    .D(_01349_),
    .Q(\fetch.bht.bhtTable_tag[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28337_ (.CLK(clock),
    .D(_01350_),
    .Q(\fetch.bht.bhtTable_tag[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28338_ (.CLK(clock),
    .D(_01351_),
    .Q(\fetch.bht.bhtTable_tag[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28339_ (.CLK(clock),
    .D(_01352_),
    .Q(\fetch.bht.bhtTable_tag[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28340_ (.CLK(clock),
    .D(_01353_),
    .Q(\fetch.bht.bhtTable_tag[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28341_ (.CLK(clock),
    .D(_01354_),
    .Q(\fetch.bht.bhtTable_tag[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28342_ (.CLK(clock),
    .D(_01355_),
    .Q(\fetch.bht.bhtTable_tag[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28343_ (.CLK(clock),
    .D(_01356_),
    .Q(\fetch.bht.bhtTable_tag[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28344_ (.CLK(clock),
    .D(_01357_),
    .Q(\fetch.bht.bhtTable_tag[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28345_ (.CLK(clock),
    .D(_01358_),
    .Q(\fetch.bht.bhtTable_tag[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28346_ (.CLK(clock),
    .D(_01359_),
    .Q(\fetch.bht.bhtTable_tag[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28347_ (.CLK(clock),
    .D(_01360_),
    .Q(\fetch.bht.bhtTable_tag[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28348_ (.CLK(clock),
    .D(_01361_),
    .Q(\fetch.bht.bhtTable_tag[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28349_ (.CLK(clock),
    .D(_01362_),
    .Q(\fetch.bht.bhtTable_tag[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28350_ (.CLK(clock),
    .D(_01363_),
    .Q(\fetch.bht.bhtTable_tag[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28351_ (.CLK(clock),
    .D(_01364_),
    .Q(\fetch.bht.bhtTable_tag[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28352_ (.CLK(clock),
    .D(_01365_),
    .Q(\fetch.bht.bhtTable_tag[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28353_ (.CLK(clock),
    .D(_01366_),
    .Q(\fetch.bht.bhtTable_tag[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28354_ (.CLK(clock),
    .D(_01367_),
    .Q(\fetch.bht.bhtTable_tag[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28355_ (.CLK(clock),
    .D(_01368_),
    .Q(\fetch.bht.bhtTable_tag[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28356_ (.CLK(clock),
    .D(_01369_),
    .Q(\fetch.bht.bhtTable_tag[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28357_ (.CLK(clock),
    .D(_01370_),
    .Q(\fetch.bht.bhtTable_tag[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28358_ (.CLK(clock),
    .D(_01371_),
    .Q(\fetch.bht.bhtTable_tag[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28359_ (.CLK(clock),
    .D(_01372_),
    .Q(\fetch.bht.bhtTable_tag[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28360_ (.CLK(clock),
    .D(_01373_),
    .Q(\fetch.bht.bhtTable_tag[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28361_ (.CLK(clock),
    .D(_01374_),
    .Q(\fetch.bht.bhtTable_tag[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28362_ (.CLK(clock),
    .D(_01375_),
    .Q(\fetch.bht.bhtTable_tag[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28363_ (.CLK(clock),
    .D(_01376_),
    .Q(\fetch.bht.bhtTable_tag[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28364_ (.CLK(clock),
    .D(_01377_),
    .Q(\fetch.bht.bhtTable_tag[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28365_ (.CLK(clock),
    .D(_01378_),
    .Q(\fetch.bht.bhtTable_tag[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28366_ (.CLK(clock),
    .D(_01379_),
    .Q(\fetch.bht.bhtTable_tag[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28367_ (.CLK(clock),
    .D(_01380_),
    .Q(\fetch.bht.bhtTable_tag[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28368_ (.CLK(clock),
    .D(_01381_),
    .Q(\fetch.bht.bhtTable_tag[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28369_ (.CLK(clock),
    .D(_01382_),
    .Q(\fetch.bht.bhtTable_tag[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28370_ (.CLK(clock),
    .D(_01383_),
    .Q(\fetch.bht.bhtTable_tag[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28371_ (.CLK(clock),
    .D(_01384_),
    .Q(\fetch.bht.bhtTable_tag[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28372_ (.CLK(clock),
    .D(_01385_),
    .Q(\fetch.bht.bhtTable_tag[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28373_ (.CLK(clock),
    .D(_01386_),
    .Q(\fetch.bht.bhtTable_tag[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28374_ (.CLK(clock),
    .D(_01387_),
    .Q(\fetch.bht.bhtTable_tag[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28375_ (.CLK(clock),
    .D(_01388_),
    .Q(\fetch.bht.bhtTable_tag[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28376_ (.CLK(clock),
    .D(_01389_),
    .Q(\fetch.bht.bhtTable_tag[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28377_ (.CLK(clock),
    .D(_01390_),
    .Q(\fetch.bht.bhtTable_tag[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28378_ (.CLK(clock),
    .D(_01391_),
    .Q(\fetch.bht.bhtTable_tag[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28379_ (.CLK(clock),
    .D(_01392_),
    .Q(\fetch.bht.bhtTable_tag[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28380_ (.CLK(clock),
    .D(_01393_),
    .Q(\fetch.bht.bhtTable_tag[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28381_ (.CLK(clock),
    .D(_01394_),
    .Q(\fetch.bht.bhtTable_tag[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28382_ (.CLK(clock),
    .D(_01395_),
    .Q(\fetch.bht.bhtTable_tag[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28383_ (.CLK(clock),
    .D(_01396_),
    .Q(io_fetch_address[2]));
 sky130_fd_sc_hd__dfxtp_2 _28384_ (.CLK(clock),
    .D(_01397_),
    .Q(io_fetch_address[3]));
 sky130_fd_sc_hd__dfxtp_2 _28385_ (.CLK(clock),
    .D(_01398_),
    .Q(io_fetch_address[4]));
 sky130_fd_sc_hd__dfxtp_2 _28386_ (.CLK(clock),
    .D(_01399_),
    .Q(io_fetch_address[5]));
 sky130_fd_sc_hd__dfxtp_2 _28387_ (.CLK(clock),
    .D(_01400_),
    .Q(io_fetch_address[6]));
 sky130_fd_sc_hd__dfxtp_2 _28388_ (.CLK(clock),
    .D(_01401_),
    .Q(io_fetch_address[7]));
 sky130_fd_sc_hd__dfxtp_2 _28389_ (.CLK(clock),
    .D(_01402_),
    .Q(io_fetch_address[8]));
 sky130_fd_sc_hd__dfxtp_2 _28390_ (.CLK(clock),
    .D(_01403_),
    .Q(io_fetch_address[9]));
 sky130_fd_sc_hd__dfxtp_2 _28391_ (.CLK(clock),
    .D(_01404_),
    .Q(io_fetch_address[10]));
 sky130_fd_sc_hd__dfxtp_2 _28392_ (.CLK(clock),
    .D(_01405_),
    .Q(io_fetch_address[11]));
 sky130_fd_sc_hd__dfxtp_2 _28393_ (.CLK(clock),
    .D(_01406_),
    .Q(io_fetch_address[12]));
 sky130_fd_sc_hd__dfxtp_2 _28394_ (.CLK(clock),
    .D(_01407_),
    .Q(io_fetch_address[13]));
 sky130_fd_sc_hd__dfxtp_2 _28395_ (.CLK(clock),
    .D(_01408_),
    .Q(io_fetch_address[14]));
 sky130_fd_sc_hd__dfxtp_2 _28396_ (.CLK(clock),
    .D(_01409_),
    .Q(io_fetch_address[15]));
 sky130_fd_sc_hd__dfxtp_2 _28397_ (.CLK(clock),
    .D(_01410_),
    .Q(io_fetch_address[16]));
 sky130_fd_sc_hd__dfxtp_2 _28398_ (.CLK(clock),
    .D(_01411_),
    .Q(io_fetch_address[17]));
 sky130_fd_sc_hd__dfxtp_2 _28399_ (.CLK(clock),
    .D(_01412_),
    .Q(io_fetch_address[18]));
 sky130_fd_sc_hd__dfxtp_2 _28400_ (.CLK(clock),
    .D(_01413_),
    .Q(io_fetch_address[19]));
 sky130_fd_sc_hd__dfxtp_2 _28401_ (.CLK(clock),
    .D(_01414_),
    .Q(io_fetch_address[20]));
 sky130_fd_sc_hd__dfxtp_2 _28402_ (.CLK(clock),
    .D(_01415_),
    .Q(io_fetch_address[21]));
 sky130_fd_sc_hd__dfxtp_2 _28403_ (.CLK(clock),
    .D(_01416_),
    .Q(io_fetch_address[22]));
 sky130_fd_sc_hd__dfxtp_2 _28404_ (.CLK(clock),
    .D(_01417_),
    .Q(io_fetch_address[23]));
 sky130_fd_sc_hd__dfxtp_2 _28405_ (.CLK(clock),
    .D(_01418_),
    .Q(io_fetch_address[24]));
 sky130_fd_sc_hd__dfxtp_2 _28406_ (.CLK(clock),
    .D(_01419_),
    .Q(io_fetch_address[25]));
 sky130_fd_sc_hd__dfxtp_2 _28407_ (.CLK(clock),
    .D(_01420_),
    .Q(io_fetch_address[26]));
 sky130_fd_sc_hd__dfxtp_2 _28408_ (.CLK(clock),
    .D(_01421_),
    .Q(io_fetch_address[27]));
 sky130_fd_sc_hd__dfxtp_2 _28409_ (.CLK(clock),
    .D(_01422_),
    .Q(io_fetch_address[28]));
 sky130_fd_sc_hd__dfxtp_2 _28410_ (.CLK(clock),
    .D(_01423_),
    .Q(io_fetch_address[29]));
 sky130_fd_sc_hd__dfxtp_2 _28411_ (.CLK(clock),
    .D(_01424_),
    .Q(io_fetch_address[30]));
 sky130_fd_sc_hd__dfxtp_2 _28412_ (.CLK(clock),
    .D(_01425_),
    .Q(io_fetch_address[31]));
 sky130_fd_sc_hd__dfxtp_2 _28413_ (.CLK(clock),
    .D(_01426_),
    .Q(\decode.control.io_opcode[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28414_ (.CLK(clock),
    .D(_01427_),
    .Q(\decode.control.io_opcode[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28415_ (.CLK(clock),
    .D(_01428_),
    .Q(\decode.control.io_opcode[5] ));
 sky130_fd_sc_hd__dfxtp_2 _28416_ (.CLK(clock),
    .D(_01429_),
    .Q(\decode.control.io_opcode[6] ));
 sky130_fd_sc_hd__dfxtp_2 _28417_ (.CLK(clock),
    .D(_01430_),
    .Q(\decode.immGen._imm_T_10[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28418_ (.CLK(clock),
    .D(_01431_),
    .Q(\decode.immGen._imm_T_10[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28419_ (.CLK(clock),
    .D(_01432_),
    .Q(\decode.immGen._imm_T_10[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28420_ (.CLK(clock),
    .D(_01433_),
    .Q(\decode.immGen._imm_T_10[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28421_ (.CLK(clock),
    .D(_01434_),
    .Q(\decode.immGen._imm_T_10[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28422_ (.CLK(clock),
    .D(_01435_),
    .Q(\decode.control.io_funct3[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28423_ (.CLK(clock),
    .D(_01436_),
    .Q(\decode.control.io_funct3[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28424_ (.CLK(clock),
    .D(_01437_),
    .Q(\decode.control.io_funct3[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28425_ (.CLK(clock),
    .D(_01438_),
    .Q(\decode.immGen._imm_T_24[15] ));
 sky130_fd_sc_hd__dfxtp_2 _28426_ (.CLK(clock),
    .D(_01439_),
    .Q(\decode.immGen._imm_T_24[16] ));
 sky130_fd_sc_hd__dfxtp_2 _28427_ (.CLK(clock),
    .D(_01440_),
    .Q(\decode.immGen._imm_T_24[17] ));
 sky130_fd_sc_hd__dfxtp_2 _28428_ (.CLK(clock),
    .D(_01441_),
    .Q(\decode.immGen._imm_T_24[18] ));
 sky130_fd_sc_hd__dfxtp_2 _28429_ (.CLK(clock),
    .D(_01442_),
    .Q(\decode.immGen._imm_T_24[19] ));
 sky130_fd_sc_hd__dfxtp_2 _28430_ (.CLK(clock),
    .D(_01443_),
    .Q(\decode.immGen._imm_T_24[11] ));
 sky130_fd_sc_hd__dfxtp_2 _28431_ (.CLK(clock),
    .D(_01444_),
    .Q(\decode.immGen._imm_T_24[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28432_ (.CLK(clock),
    .D(_01445_),
    .Q(\decode.immGen._imm_T_24[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28433_ (.CLK(clock),
    .D(_01446_),
    .Q(\decode.immGen._imm_T_24[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28434_ (.CLK(clock),
    .D(_01447_),
    .Q(\decode.immGen._imm_T_24[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28435_ (.CLK(clock),
    .D(_01448_),
    .Q(\decode.control.io_funct7[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28436_ (.CLK(clock),
    .D(_01449_),
    .Q(\decode.control.io_funct7[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28437_ (.CLK(clock),
    .D(_01450_),
    .Q(\decode.control.io_funct7[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28438_ (.CLK(clock),
    .D(_01451_),
    .Q(\decode.control.io_funct7[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28439_ (.CLK(clock),
    .D(_01452_),
    .Q(\decode.control.io_funct7[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28440_ (.CLK(clock),
    .D(_01453_),
    .Q(\decode.control.io_funct7[5] ));
 sky130_fd_sc_hd__dfxtp_2 _28441_ (.CLK(clock),
    .D(_01454_),
    .Q(\decode.control.io_funct7[6] ));
 sky130_fd_sc_hd__dfxtp_2 _28442_ (.CLK(clock),
    .D(_01455_),
    .Q(\decode.io_id_pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _28443_ (.CLK(clock),
    .D(_01456_),
    .Q(\decode.io_id_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _28444_ (.CLK(clock),
    .D(_01457_),
    .Q(\decode.io_id_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _28445_ (.CLK(clock),
    .D(_01458_),
    .Q(\decode.io_id_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _28446_ (.CLK(clock),
    .D(_01459_),
    .Q(\decode.io_id_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _28447_ (.CLK(clock),
    .D(_01460_),
    .Q(\decode.io_id_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _28448_ (.CLK(clock),
    .D(_01461_),
    .Q(\decode.io_id_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _28449_ (.CLK(clock),
    .D(_01462_),
    .Q(\decode.io_id_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _28450_ (.CLK(clock),
    .D(_01463_),
    .Q(\decode.io_id_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _28451_ (.CLK(clock),
    .D(_01464_),
    .Q(\decode.io_id_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _28452_ (.CLK(clock),
    .D(_01465_),
    .Q(\decode.io_id_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _28453_ (.CLK(clock),
    .D(_01466_),
    .Q(\decode.io_id_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _28454_ (.CLK(clock),
    .D(_01467_),
    .Q(\decode.io_id_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _28455_ (.CLK(clock),
    .D(_01468_),
    .Q(\decode.io_id_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _28456_ (.CLK(clock),
    .D(_01469_),
    .Q(\decode.io_id_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _28457_ (.CLK(clock),
    .D(_01470_),
    .Q(\decode.io_id_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _28458_ (.CLK(clock),
    .D(_01471_),
    .Q(\decode.io_id_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _28459_ (.CLK(clock),
    .D(_01472_),
    .Q(\decode.io_id_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _28460_ (.CLK(clock),
    .D(_01473_),
    .Q(\decode.io_id_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _28461_ (.CLK(clock),
    .D(_01474_),
    .Q(\decode.io_id_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _28462_ (.CLK(clock),
    .D(_01475_),
    .Q(\decode.io_id_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _28463_ (.CLK(clock),
    .D(_01476_),
    .Q(\decode.io_id_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _28464_ (.CLK(clock),
    .D(_01477_),
    .Q(\decode.io_id_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _28465_ (.CLK(clock),
    .D(_01478_),
    .Q(\decode.io_id_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _28466_ (.CLK(clock),
    .D(_01479_),
    .Q(\decode.io_id_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _28467_ (.CLK(clock),
    .D(_01480_),
    .Q(\decode.io_id_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _28468_ (.CLK(clock),
    .D(_01481_),
    .Q(\decode.io_id_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _28469_ (.CLK(clock),
    .D(_01482_),
    .Q(\decode.io_id_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _28470_ (.CLK(clock),
    .D(_01483_),
    .Q(\decode.io_id_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _28471_ (.CLK(clock),
    .D(_01484_),
    .Q(\decode.io_id_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _28472_ (.CLK(clock),
    .D(_01485_),
    .Q(\decode.io_id_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _28473_ (.CLK(clock),
    .D(_01486_),
    .Q(\decode.io_id_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _28474_ (.CLK(clock),
    .D(_01487_),
    .Q(\fetch.bht.bhtTable_tag[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28475_ (.CLK(clock),
    .D(_01488_),
    .Q(\fetch.bht.bhtTable_tag[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28476_ (.CLK(clock),
    .D(_01489_),
    .Q(\fetch.bht.bhtTable_tag[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28477_ (.CLK(clock),
    .D(_01490_),
    .Q(\fetch.bht.bhtTable_tag[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28478_ (.CLK(clock),
    .D(_01491_),
    .Q(\fetch.bht.bhtTable_tag[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28479_ (.CLK(clock),
    .D(_01492_),
    .Q(\fetch.bht.bhtTable_tag[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28480_ (.CLK(clock),
    .D(_01493_),
    .Q(\fetch.bht.bhtTable_tag[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28481_ (.CLK(clock),
    .D(_01494_),
    .Q(\fetch.bht.bhtTable_tag[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28482_ (.CLK(clock),
    .D(_01495_),
    .Q(\fetch.bht.bhtTable_tag[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28483_ (.CLK(clock),
    .D(_01496_),
    .Q(\fetch.bht.bhtTable_tag[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28484_ (.CLK(clock),
    .D(_01497_),
    .Q(\fetch.bht.bhtTable_tag[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28485_ (.CLK(clock),
    .D(_01498_),
    .Q(\fetch.bht.bhtTable_tag[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28486_ (.CLK(clock),
    .D(_01499_),
    .Q(\fetch.bht.bhtTable_tag[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28487_ (.CLK(clock),
    .D(_01500_),
    .Q(\fetch.bht.bhtTable_tag[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28488_ (.CLK(clock),
    .D(_01501_),
    .Q(\fetch.bht.bhtTable_tag[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28489_ (.CLK(clock),
    .D(_01502_),
    .Q(\fetch.bht.bhtTable_tag[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28490_ (.CLK(clock),
    .D(_01503_),
    .Q(\fetch.bht.bhtTable_tag[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28491_ (.CLK(clock),
    .D(_01504_),
    .Q(\fetch.bht.bhtTable_tag[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28492_ (.CLK(clock),
    .D(_01505_),
    .Q(\fetch.bht.bhtTable_tag[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28493_ (.CLK(clock),
    .D(_01506_),
    .Q(\fetch.bht.bhtTable_tag[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28494_ (.CLK(clock),
    .D(_01507_),
    .Q(\fetch.bht.bhtTable_tag[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28495_ (.CLK(clock),
    .D(_01508_),
    .Q(\fetch.bht.bhtTable_tag[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28496_ (.CLK(clock),
    .D(_01509_),
    .Q(\fetch.bht.bhtTable_tag[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28497_ (.CLK(clock),
    .D(_01510_),
    .Q(\fetch.bht.bhtTable_tag[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28498_ (.CLK(clock),
    .D(_01511_),
    .Q(\fetch.bht.bhtTable_tag[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28499_ (.CLK(clock),
    .D(_01512_),
    .Q(\fetch.bht.bhtTable_tag[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28500_ (.CLK(clock),
    .D(_01513_),
    .Q(\fetch.bht.bhtTable_tag[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28501_ (.CLK(clock),
    .D(_01514_),
    .Q(\fetch.bht.bhtTable_tag[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28502_ (.CLK(clock),
    .D(_01515_),
    .Q(\fetch.bht.bhtTable_tag[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28503_ (.CLK(clock),
    .D(_01516_),
    .Q(\fetch.bht.bhtTable_tag[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28504_ (.CLK(clock),
    .D(_01517_),
    .Q(\fetch.bht.bhtTable_tag[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28505_ (.CLK(clock),
    .D(_01518_),
    .Q(\fetch.bht.bhtTable_tag[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28506_ (.CLK(clock),
    .D(_01519_),
    .Q(\fetch.bht.bhtTable_tag[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28507_ (.CLK(clock),
    .D(_01520_),
    .Q(\fetch.bht.bhtTable_tag[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28508_ (.CLK(clock),
    .D(_01521_),
    .Q(\fetch.bht.bhtTable_tag[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28509_ (.CLK(clock),
    .D(_01522_),
    .Q(\fetch.bht.bhtTable_tag[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28510_ (.CLK(clock),
    .D(_01523_),
    .Q(\fetch.bht.bhtTable_tag[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28511_ (.CLK(clock),
    .D(_01524_),
    .Q(\fetch.bht.bhtTable_tag[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28512_ (.CLK(clock),
    .D(_01525_),
    .Q(\fetch.bht.bhtTable_tag[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28513_ (.CLK(clock),
    .D(_01526_),
    .Q(\fetch.bht.bhtTable_tag[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28514_ (.CLK(clock),
    .D(_01527_),
    .Q(\fetch.bht.bhtTable_tag[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28515_ (.CLK(clock),
    .D(_01528_),
    .Q(\fetch.bht.bhtTable_tag[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28516_ (.CLK(clock),
    .D(_01529_),
    .Q(\fetch.bht.bhtTable_tag[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28517_ (.CLK(clock),
    .D(_01530_),
    .Q(\fetch.bht.bhtTable_tag[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28518_ (.CLK(clock),
    .D(_01531_),
    .Q(\fetch.bht.bhtTable_tag[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28519_ (.CLK(clock),
    .D(_01532_),
    .Q(\fetch.bht.bhtTable_tag[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28520_ (.CLK(clock),
    .D(_01533_),
    .Q(\fetch.bht.bhtTable_tag[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28521_ (.CLK(clock),
    .D(_01534_),
    .Q(\fetch.bht.bhtTable_tag[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28522_ (.CLK(clock),
    .D(_01535_),
    .Q(\fetch.bht.bhtTable_tag[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28523_ (.CLK(clock),
    .D(_01536_),
    .Q(\fetch.bht.bhtTable_tag[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28524_ (.CLK(clock),
    .D(_01537_),
    .Q(\fetch.bht.bhtTable_tag[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28525_ (.CLK(clock),
    .D(_01538_),
    .Q(\fetch.bht.bhtTable_tag[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28526_ (.CLK(clock),
    .D(_01539_),
    .Q(\fetch.bht.bhtTable_tag[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28527_ (.CLK(clock),
    .D(_01540_),
    .Q(\fetch.bht.bhtTable_tag[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28528_ (.CLK(clock),
    .D(_01541_),
    .Q(\fetch.bht.bhtTable_tag[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28529_ (.CLK(clock),
    .D(_01542_),
    .Q(\fetch.bht.bhtTable_tag[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28530_ (.CLK(clock),
    .D(_01543_),
    .Q(\fetch.bht.bhtTable_tag[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28531_ (.CLK(clock),
    .D(_01544_),
    .Q(\fetch.bht.bhtTable_tag[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28532_ (.CLK(clock),
    .D(_01545_),
    .Q(\fetch.bht.bhtTable_tag[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28533_ (.CLK(clock),
    .D(_01546_),
    .Q(\fetch.bht.bhtTable_tag[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28534_ (.CLK(clock),
    .D(_01547_),
    .Q(\fetch.bht.bhtTable_tag[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28535_ (.CLK(clock),
    .D(_01548_),
    .Q(\fetch.bht.bhtTable_tag[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28536_ (.CLK(clock),
    .D(_01549_),
    .Q(\fetch.bht.bhtTable_tag[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28537_ (.CLK(clock),
    .D(_01550_),
    .Q(\fetch.bht.bhtTable_tag[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28538_ (.CLK(clock),
    .D(_01551_),
    .Q(\fetch.bht.bhtTable_tag[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28539_ (.CLK(clock),
    .D(_01552_),
    .Q(\fetch.bht.bhtTable_tag[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28540_ (.CLK(clock),
    .D(_01553_),
    .Q(\fetch.bht.bhtTable_tag[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28541_ (.CLK(clock),
    .D(_01554_),
    .Q(\fetch.bht.bhtTable_tag[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28542_ (.CLK(clock),
    .D(_01555_),
    .Q(\fetch.bht.bhtTable_tag[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28543_ (.CLK(clock),
    .D(_01556_),
    .Q(\fetch.bht.bhtTable_tag[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28544_ (.CLK(clock),
    .D(_01557_),
    .Q(\fetch.bht.bhtTable_tag[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28545_ (.CLK(clock),
    .D(_01558_),
    .Q(\fetch.bht.bhtTable_tag[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28546_ (.CLK(clock),
    .D(_01559_),
    .Q(\fetch.bht.bhtTable_tag[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28547_ (.CLK(clock),
    .D(_01560_),
    .Q(\fetch.bht.bhtTable_tag[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28548_ (.CLK(clock),
    .D(_01561_),
    .Q(\fetch.bht.bhtTable_tag[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28549_ (.CLK(clock),
    .D(_01562_),
    .Q(\fetch.bht.bhtTable_tag[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28550_ (.CLK(clock),
    .D(_01563_),
    .Q(\fetch.bht.bhtTable_tag[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28551_ (.CLK(clock),
    .D(_01564_),
    .Q(\fetch.bht.bhtTable_tag[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28552_ (.CLK(clock),
    .D(_01565_),
    .Q(\fetch.bht.bhtTable_tag[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28553_ (.CLK(clock),
    .D(_01566_),
    .Q(\fetch.bht.bhtTable_tag[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28554_ (.CLK(clock),
    .D(_01567_),
    .Q(\fetch.bht.bhtTable_tag[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28555_ (.CLK(clock),
    .D(_01568_),
    .Q(\fetch.bht.bhtTable_tag[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28556_ (.CLK(clock),
    .D(_01569_),
    .Q(\fetch.bht.bhtTable_tag[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28557_ (.CLK(clock),
    .D(_01570_),
    .Q(\fetch.bht.bhtTable_tag[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28558_ (.CLK(clock),
    .D(_01571_),
    .Q(\fetch.bht.bhtTable_tag[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28559_ (.CLK(clock),
    .D(_01572_),
    .Q(\fetch.bht.bhtTable_tag[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28560_ (.CLK(clock),
    .D(_01573_),
    .Q(\fetch.bht.bhtTable_tag[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28561_ (.CLK(clock),
    .D(_01574_),
    .Q(\fetch.bht.bhtTable_tag[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28562_ (.CLK(clock),
    .D(_01575_),
    .Q(\fetch.bht.bhtTable_tag[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28563_ (.CLK(clock),
    .D(_01576_),
    .Q(\fetch.bht.bhtTable_tag[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28564_ (.CLK(clock),
    .D(_01577_),
    .Q(\fetch.bht.bhtTable_tag[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28565_ (.CLK(clock),
    .D(_01578_),
    .Q(\fetch.bht.bhtTable_tag[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28566_ (.CLK(clock),
    .D(_01579_),
    .Q(\fetch.bht.bhtTable_tag[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28567_ (.CLK(clock),
    .D(_01580_),
    .Q(\fetch.bht.bhtTable_tag[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28568_ (.CLK(clock),
    .D(_01581_),
    .Q(\fetch.bht.bhtTable_tag[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28569_ (.CLK(clock),
    .D(_01582_),
    .Q(\fetch.bht.bhtTable_tag[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28570_ (.CLK(clock),
    .D(_01583_),
    .Q(\fetch.bht.bhtTable_tag[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28571_ (.CLK(clock),
    .D(_01584_),
    .Q(\fetch.bht.bhtTable_tag[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28572_ (.CLK(clock),
    .D(_01585_),
    .Q(\fetch.bht.bhtTable_tag[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28573_ (.CLK(clock),
    .D(_01586_),
    .Q(\fetch.bht.bhtTable_tag[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28574_ (.CLK(clock),
    .D(_01587_),
    .Q(\fetch.bht.bhtTable_tag[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28575_ (.CLK(clock),
    .D(_01588_),
    .Q(\fetch.bht.bhtTable_tag[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28576_ (.CLK(clock),
    .D(_01589_),
    .Q(\fetch.bht.bhtTable_tag[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28577_ (.CLK(clock),
    .D(_01590_),
    .Q(\fetch.bht.bhtTable_tag[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28578_ (.CLK(clock),
    .D(_01591_),
    .Q(\fetch.bht.bhtTable_target_pc[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28579_ (.CLK(clock),
    .D(_01592_),
    .Q(\fetch.bht.bhtTable_target_pc[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28580_ (.CLK(clock),
    .D(_01593_),
    .Q(\fetch.bht.bhtTable_target_pc[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28581_ (.CLK(clock),
    .D(_01594_),
    .Q(\fetch.bht.bhtTable_target_pc[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28582_ (.CLK(clock),
    .D(_01595_),
    .Q(\fetch.bht.bhtTable_target_pc[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28583_ (.CLK(clock),
    .D(_01596_),
    .Q(\fetch.bht.bhtTable_target_pc[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28584_ (.CLK(clock),
    .D(_01597_),
    .Q(\fetch.bht.bhtTable_target_pc[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28585_ (.CLK(clock),
    .D(_01598_),
    .Q(\fetch.bht.bhtTable_target_pc[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28586_ (.CLK(clock),
    .D(_01599_),
    .Q(\fetch.bht.bhtTable_target_pc[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28587_ (.CLK(clock),
    .D(_01600_),
    .Q(\fetch.bht.bhtTable_target_pc[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28588_ (.CLK(clock),
    .D(_01601_),
    .Q(\fetch.bht.bhtTable_target_pc[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28589_ (.CLK(clock),
    .D(_01602_),
    .Q(\fetch.bht.bhtTable_target_pc[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28590_ (.CLK(clock),
    .D(_01603_),
    .Q(\fetch.bht.bhtTable_target_pc[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28591_ (.CLK(clock),
    .D(_01604_),
    .Q(\fetch.bht.bhtTable_target_pc[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28592_ (.CLK(clock),
    .D(_01605_),
    .Q(\fetch.bht.bhtTable_target_pc[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28593_ (.CLK(clock),
    .D(_01606_),
    .Q(\fetch.bht.bhtTable_target_pc[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28594_ (.CLK(clock),
    .D(_01607_),
    .Q(\fetch.bht.bhtTable_target_pc[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28595_ (.CLK(clock),
    .D(_01608_),
    .Q(\fetch.bht.bhtTable_target_pc[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28596_ (.CLK(clock),
    .D(_01609_),
    .Q(\fetch.bht.bhtTable_target_pc[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28597_ (.CLK(clock),
    .D(_01610_),
    .Q(\fetch.bht.bhtTable_target_pc[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28598_ (.CLK(clock),
    .D(_01611_),
    .Q(\fetch.bht.bhtTable_target_pc[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28599_ (.CLK(clock),
    .D(_01612_),
    .Q(\fetch.bht.bhtTable_target_pc[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28600_ (.CLK(clock),
    .D(_01613_),
    .Q(\fetch.bht.bhtTable_target_pc[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28601_ (.CLK(clock),
    .D(_01614_),
    .Q(\fetch.bht.bhtTable_target_pc[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28602_ (.CLK(clock),
    .D(_01615_),
    .Q(\fetch.bht.bhtTable_target_pc[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28603_ (.CLK(clock),
    .D(_01616_),
    .Q(\fetch.bht.bhtTable_target_pc[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28604_ (.CLK(clock),
    .D(_01617_),
    .Q(\fetch.bht.bhtTable_target_pc[15][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28605_ (.CLK(clock),
    .D(_01618_),
    .Q(\fetch.bht.bhtTable_target_pc[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28606_ (.CLK(clock),
    .D(_01619_),
    .Q(\fetch.bht.bhtTable_target_pc[15][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28607_ (.CLK(clock),
    .D(_01620_),
    .Q(\fetch.bht.bhtTable_target_pc[15][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28608_ (.CLK(clock),
    .D(_01621_),
    .Q(\fetch.bht.bhtTable_target_pc[15][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28609_ (.CLK(clock),
    .D(_01622_),
    .Q(\fetch.bht.bhtTable_target_pc[15][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28610_ (.CLK(clock),
    .D(_01623_),
    .Q(\fetch.bht.bhtTable_target_pc[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28611_ (.CLK(clock),
    .D(_01624_),
    .Q(\fetch.bht.bhtTable_target_pc[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28612_ (.CLK(clock),
    .D(_01625_),
    .Q(\fetch.bht.bhtTable_target_pc[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28613_ (.CLK(clock),
    .D(_01626_),
    .Q(\fetch.bht.bhtTable_target_pc[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28614_ (.CLK(clock),
    .D(_01627_),
    .Q(\fetch.bht.bhtTable_target_pc[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28615_ (.CLK(clock),
    .D(_01628_),
    .Q(\fetch.bht.bhtTable_target_pc[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28616_ (.CLK(clock),
    .D(_01629_),
    .Q(\fetch.bht.bhtTable_target_pc[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28617_ (.CLK(clock),
    .D(_01630_),
    .Q(\fetch.bht.bhtTable_target_pc[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28618_ (.CLK(clock),
    .D(_01631_),
    .Q(\fetch.bht.bhtTable_target_pc[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28619_ (.CLK(clock),
    .D(_01632_),
    .Q(\fetch.bht.bhtTable_target_pc[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28620_ (.CLK(clock),
    .D(_01633_),
    .Q(\fetch.bht.bhtTable_target_pc[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28621_ (.CLK(clock),
    .D(_01634_),
    .Q(\fetch.bht.bhtTable_target_pc[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28622_ (.CLK(clock),
    .D(_01635_),
    .Q(\fetch.bht.bhtTable_target_pc[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28623_ (.CLK(clock),
    .D(_01636_),
    .Q(\fetch.bht.bhtTable_target_pc[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28624_ (.CLK(clock),
    .D(_01637_),
    .Q(\fetch.bht.bhtTable_target_pc[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28625_ (.CLK(clock),
    .D(_01638_),
    .Q(\fetch.bht.bhtTable_target_pc[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28626_ (.CLK(clock),
    .D(_01639_),
    .Q(\fetch.bht.bhtTable_target_pc[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28627_ (.CLK(clock),
    .D(_01640_),
    .Q(\fetch.bht.bhtTable_target_pc[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28628_ (.CLK(clock),
    .D(_01641_),
    .Q(\fetch.bht.bhtTable_target_pc[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28629_ (.CLK(clock),
    .D(_01642_),
    .Q(\fetch.bht.bhtTable_target_pc[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28630_ (.CLK(clock),
    .D(_01643_),
    .Q(\fetch.bht.bhtTable_target_pc[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28631_ (.CLK(clock),
    .D(_01644_),
    .Q(\fetch.bht.bhtTable_target_pc[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28632_ (.CLK(clock),
    .D(_01645_),
    .Q(\fetch.bht.bhtTable_target_pc[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28633_ (.CLK(clock),
    .D(_01646_),
    .Q(\fetch.bht.bhtTable_target_pc[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28634_ (.CLK(clock),
    .D(_01647_),
    .Q(\fetch.bht.bhtTable_target_pc[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28635_ (.CLK(clock),
    .D(_01648_),
    .Q(\fetch.bht.bhtTable_target_pc[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28636_ (.CLK(clock),
    .D(_01649_),
    .Q(\fetch.bht.bhtTable_target_pc[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28637_ (.CLK(clock),
    .D(_01650_),
    .Q(\fetch.bht.bhtTable_target_pc[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28638_ (.CLK(clock),
    .D(_01651_),
    .Q(\fetch.bht.bhtTable_target_pc[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28639_ (.CLK(clock),
    .D(_01652_),
    .Q(\fetch.bht.bhtTable_target_pc[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28640_ (.CLK(clock),
    .D(_01653_),
    .Q(\fetch.bht.bhtTable_target_pc[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28641_ (.CLK(clock),
    .D(_01654_),
    .Q(\fetch.bht.bhtTable_target_pc[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28642_ (.CLK(clock),
    .D(_01655_),
    .Q(\fetch.bht.bhtTable_target_pc[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28643_ (.CLK(clock),
    .D(_01656_),
    .Q(\fetch.bht.bhtTable_target_pc[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28644_ (.CLK(clock),
    .D(_01657_),
    .Q(\fetch.bht.bhtTable_target_pc[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28645_ (.CLK(clock),
    .D(_01658_),
    .Q(\fetch.bht.bhtTable_target_pc[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28646_ (.CLK(clock),
    .D(_01659_),
    .Q(\fetch.bht.bhtTable_target_pc[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28647_ (.CLK(clock),
    .D(_01660_),
    .Q(\fetch.bht.bhtTable_target_pc[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28648_ (.CLK(clock),
    .D(_01661_),
    .Q(\fetch.bht.bhtTable_target_pc[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28649_ (.CLK(clock),
    .D(_01662_),
    .Q(\fetch.bht.bhtTable_target_pc[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28650_ (.CLK(clock),
    .D(_01663_),
    .Q(\fetch.bht.bhtTable_target_pc[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28651_ (.CLK(clock),
    .D(_01664_),
    .Q(\fetch.bht.bhtTable_target_pc[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28652_ (.CLK(clock),
    .D(_01665_),
    .Q(\fetch.bht.bhtTable_target_pc[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28653_ (.CLK(clock),
    .D(_01666_),
    .Q(\fetch.bht.bhtTable_target_pc[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28654_ (.CLK(clock),
    .D(_01667_),
    .Q(\fetch.bht.bhtTable_target_pc[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28655_ (.CLK(clock),
    .D(_01668_),
    .Q(\fetch.bht.bhtTable_target_pc[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28656_ (.CLK(clock),
    .D(_01669_),
    .Q(\fetch.bht.bhtTable_target_pc[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28657_ (.CLK(clock),
    .D(_01670_),
    .Q(\fetch.bht.bhtTable_target_pc[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28658_ (.CLK(clock),
    .D(_01671_),
    .Q(\fetch.bht.bhtTable_target_pc[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28659_ (.CLK(clock),
    .D(_01672_),
    .Q(\fetch.bht.bhtTable_target_pc[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28660_ (.CLK(clock),
    .D(_01673_),
    .Q(\fetch.bht.bhtTable_target_pc[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28661_ (.CLK(clock),
    .D(_01674_),
    .Q(\fetch.bht.bhtTable_target_pc[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28662_ (.CLK(clock),
    .D(_01675_),
    .Q(\fetch.bht.bhtTable_target_pc[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28663_ (.CLK(clock),
    .D(_01676_),
    .Q(\fetch.bht.bhtTable_target_pc[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28664_ (.CLK(clock),
    .D(_01677_),
    .Q(\fetch.bht.bhtTable_target_pc[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28665_ (.CLK(clock),
    .D(_01678_),
    .Q(\fetch.bht.bhtTable_target_pc[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28666_ (.CLK(clock),
    .D(_01679_),
    .Q(\fetch.bht.bhtTable_target_pc[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28667_ (.CLK(clock),
    .D(_01680_),
    .Q(\fetch.bht.bhtTable_target_pc[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28668_ (.CLK(clock),
    .D(_01681_),
    .Q(\fetch.bht.bhtTable_target_pc[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28669_ (.CLK(clock),
    .D(_01682_),
    .Q(\fetch.bht.bhtTable_target_pc[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28670_ (.CLK(clock),
    .D(_01683_),
    .Q(\fetch.bht.bhtTable_target_pc[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28671_ (.CLK(clock),
    .D(_01684_),
    .Q(\fetch.bht.bhtTable_target_pc[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28672_ (.CLK(clock),
    .D(_01685_),
    .Q(\fetch.bht.bhtTable_target_pc[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28673_ (.CLK(clock),
    .D(_01686_),
    .Q(\fetch.bht.bhtTable_target_pc[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28674_ (.CLK(clock),
    .D(_01687_),
    .Q(\fetch.bht.bhtTable_target_pc[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28675_ (.CLK(clock),
    .D(_01688_),
    .Q(\fetch.bht.bhtTable_target_pc[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28676_ (.CLK(clock),
    .D(_01689_),
    .Q(\fetch.bht.bhtTable_target_pc[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28677_ (.CLK(clock),
    .D(_01690_),
    .Q(\fetch.bht.bhtTable_target_pc[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28678_ (.CLK(clock),
    .D(_01691_),
    .Q(\fetch.bht.bhtTable_target_pc[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28679_ (.CLK(clock),
    .D(_01692_),
    .Q(\fetch.bht.bhtTable_target_pc[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28680_ (.CLK(clock),
    .D(_01693_),
    .Q(\fetch.bht.bhtTable_target_pc[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28681_ (.CLK(clock),
    .D(_01694_),
    .Q(\fetch.bht.bhtTable_target_pc[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28682_ (.CLK(clock),
    .D(_01695_),
    .Q(\fetch.bht.bhtTable_target_pc[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28683_ (.CLK(clock),
    .D(_01696_),
    .Q(\fetch.bht.bhtTable_target_pc[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28684_ (.CLK(clock),
    .D(_01697_),
    .Q(\fetch.bht.bhtTable_target_pc[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28685_ (.CLK(clock),
    .D(_01698_),
    .Q(\fetch.bht.bhtTable_target_pc[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28686_ (.CLK(clock),
    .D(_01699_),
    .Q(\fetch.bht.bhtTable_target_pc[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28687_ (.CLK(clock),
    .D(_01700_),
    .Q(\fetch.bht.bhtTable_target_pc[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28688_ (.CLK(clock),
    .D(_01701_),
    .Q(\fetch.bht.bhtTable_target_pc[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28689_ (.CLK(clock),
    .D(_01702_),
    .Q(\fetch.bht.bhtTable_target_pc[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28690_ (.CLK(clock),
    .D(_01703_),
    .Q(\fetch.bht.bhtTable_target_pc[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28691_ (.CLK(clock),
    .D(_01704_),
    .Q(\fetch.bht.bhtTable_target_pc[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28692_ (.CLK(clock),
    .D(_01705_),
    .Q(\fetch.bht.bhtTable_target_pc[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28693_ (.CLK(clock),
    .D(_01706_),
    .Q(\fetch.bht.bhtTable_target_pc[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28694_ (.CLK(clock),
    .D(_01707_),
    .Q(\fetch.bht.bhtTable_target_pc[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28695_ (.CLK(clock),
    .D(_01708_),
    .Q(\fetch.bht.bhtTable_target_pc[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28696_ (.CLK(clock),
    .D(_01709_),
    .Q(\fetch.bht.bhtTable_target_pc[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28697_ (.CLK(clock),
    .D(_01710_),
    .Q(\fetch.bht.bhtTable_target_pc[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28698_ (.CLK(clock),
    .D(_01711_),
    .Q(\fetch.bht.bhtTable_target_pc[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28699_ (.CLK(clock),
    .D(_01712_),
    .Q(\fetch.bht.bhtTable_target_pc[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28700_ (.CLK(clock),
    .D(_01713_),
    .Q(\fetch.bht.bhtTable_target_pc[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28701_ (.CLK(clock),
    .D(_01714_),
    .Q(\fetch.bht.bhtTable_target_pc[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28702_ (.CLK(clock),
    .D(_01715_),
    .Q(\fetch.bht.bhtTable_target_pc[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28703_ (.CLK(clock),
    .D(_01716_),
    .Q(\fetch.bht.bhtTable_target_pc[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28704_ (.CLK(clock),
    .D(_01717_),
    .Q(\fetch.bht.bhtTable_target_pc[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28705_ (.CLK(clock),
    .D(_01718_),
    .Q(\fetch.bht.bhtTable_target_pc[3][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28706_ (.CLK(clock),
    .D(_01719_),
    .Q(\fetch.bht.bhtTable_target_pc[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28707_ (.CLK(clock),
    .D(_01720_),
    .Q(\fetch.bht.bhtTable_target_pc[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28708_ (.CLK(clock),
    .D(_01721_),
    .Q(\fetch.bht.bhtTable_target_pc[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28709_ (.CLK(clock),
    .D(_01722_),
    .Q(\fetch.bht.bhtTable_target_pc[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28710_ (.CLK(clock),
    .D(_01723_),
    .Q(\fetch.bht.bhtTable_target_pc[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28711_ (.CLK(clock),
    .D(_01724_),
    .Q(\fetch.bht.bhtTable_target_pc[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28712_ (.CLK(clock),
    .D(_01725_),
    .Q(\fetch.bht.bhtTable_target_pc[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28713_ (.CLK(clock),
    .D(_01726_),
    .Q(\fetch.bht.bhtTable_target_pc[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28714_ (.CLK(clock),
    .D(_01727_),
    .Q(\fetch.bht.bhtTable_target_pc[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28715_ (.CLK(clock),
    .D(_01728_),
    .Q(\fetch.bht.bhtTable_target_pc[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28716_ (.CLK(clock),
    .D(_01729_),
    .Q(\fetch.bht.bhtTable_target_pc[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28717_ (.CLK(clock),
    .D(_01730_),
    .Q(\fetch.bht.bhtTable_target_pc[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28718_ (.CLK(clock),
    .D(_01731_),
    .Q(\fetch.bht.bhtTable_target_pc[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28719_ (.CLK(clock),
    .D(_01732_),
    .Q(\fetch.bht.bhtTable_target_pc[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28720_ (.CLK(clock),
    .D(_01733_),
    .Q(\fetch.bht.bhtTable_target_pc[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28721_ (.CLK(clock),
    .D(_01734_),
    .Q(\fetch.bht.bhtTable_target_pc[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28722_ (.CLK(clock),
    .D(_01735_),
    .Q(\fetch.bht.bhtTable_target_pc[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28723_ (.CLK(clock),
    .D(_01736_),
    .Q(\fetch.bht.bhtTable_target_pc[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28724_ (.CLK(clock),
    .D(_01737_),
    .Q(\fetch.bht.bhtTable_target_pc[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28725_ (.CLK(clock),
    .D(_01738_),
    .Q(\fetch.bht.bhtTable_target_pc[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28726_ (.CLK(clock),
    .D(_01739_),
    .Q(\fetch.bht.bhtTable_target_pc[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28727_ (.CLK(clock),
    .D(_01740_),
    .Q(\fetch.bht.bhtTable_target_pc[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28728_ (.CLK(clock),
    .D(_01741_),
    .Q(\fetch.bht.bhtTable_target_pc[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28729_ (.CLK(clock),
    .D(_01742_),
    .Q(\fetch.bht.bhtTable_target_pc[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28730_ (.CLK(clock),
    .D(_01743_),
    .Q(\fetch.bht.bhtTable_target_pc[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28731_ (.CLK(clock),
    .D(_01744_),
    .Q(\fetch.bht.bhtTable_target_pc[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28732_ (.CLK(clock),
    .D(_01745_),
    .Q(\fetch.bht.bhtTable_target_pc[4][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28733_ (.CLK(clock),
    .D(_01746_),
    .Q(\fetch.bht.bhtTable_target_pc[4][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28734_ (.CLK(clock),
    .D(_01747_),
    .Q(\fetch.bht.bhtTable_target_pc[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28735_ (.CLK(clock),
    .D(_01748_),
    .Q(\fetch.bht.bhtTable_target_pc[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28736_ (.CLK(clock),
    .D(_01749_),
    .Q(\fetch.bht.bhtTable_target_pc[4][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28737_ (.CLK(clock),
    .D(_01750_),
    .Q(\fetch.bht.bhtTable_target_pc[4][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28738_ (.CLK(clock),
    .D(_01751_),
    .Q(\fetch.bht.bhtTable_target_pc[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28739_ (.CLK(clock),
    .D(_01752_),
    .Q(\fetch.bht.bhtTable_target_pc[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28740_ (.CLK(clock),
    .D(_01753_),
    .Q(\fetch.bht.bhtTable_target_pc[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28741_ (.CLK(clock),
    .D(_01754_),
    .Q(\fetch.bht.bhtTable_target_pc[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28742_ (.CLK(clock),
    .D(_01755_),
    .Q(\fetch.bht.bhtTable_target_pc[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28743_ (.CLK(clock),
    .D(_01756_),
    .Q(\fetch.bht.bhtTable_target_pc[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28744_ (.CLK(clock),
    .D(_01757_),
    .Q(\fetch.bht.bhtTable_target_pc[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28745_ (.CLK(clock),
    .D(_01758_),
    .Q(\fetch.bht.bhtTable_target_pc[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28746_ (.CLK(clock),
    .D(_01759_),
    .Q(\fetch.bht.bhtTable_target_pc[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28747_ (.CLK(clock),
    .D(_01760_),
    .Q(\fetch.bht.bhtTable_target_pc[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28748_ (.CLK(clock),
    .D(_01761_),
    .Q(\fetch.bht.bhtTable_target_pc[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28749_ (.CLK(clock),
    .D(_01762_),
    .Q(\fetch.bht.bhtTable_target_pc[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28750_ (.CLK(clock),
    .D(_01763_),
    .Q(\fetch.bht.bhtTable_target_pc[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28751_ (.CLK(clock),
    .D(_01764_),
    .Q(\fetch.bht.bhtTable_target_pc[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28752_ (.CLK(clock),
    .D(_01765_),
    .Q(\fetch.bht.bhtTable_target_pc[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28753_ (.CLK(clock),
    .D(_01766_),
    .Q(\fetch.bht.bhtTable_target_pc[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28754_ (.CLK(clock),
    .D(_01767_),
    .Q(\fetch.bht.bhtTable_target_pc[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28755_ (.CLK(clock),
    .D(_01768_),
    .Q(\fetch.bht.bhtTable_target_pc[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28756_ (.CLK(clock),
    .D(_01769_),
    .Q(\fetch.bht.bhtTable_target_pc[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28757_ (.CLK(clock),
    .D(_01770_),
    .Q(\fetch.bht.bhtTable_target_pc[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28758_ (.CLK(clock),
    .D(_01771_),
    .Q(\fetch.bht.bhtTable_target_pc[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28759_ (.CLK(clock),
    .D(_01772_),
    .Q(\fetch.bht.bhtTable_target_pc[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28760_ (.CLK(clock),
    .D(_01773_),
    .Q(\fetch.bht.bhtTable_target_pc[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28761_ (.CLK(clock),
    .D(_01774_),
    .Q(\fetch.bht.bhtTable_target_pc[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28762_ (.CLK(clock),
    .D(_01775_),
    .Q(\fetch.bht.bhtTable_target_pc[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28763_ (.CLK(clock),
    .D(_01776_),
    .Q(\fetch.bht.bhtTable_target_pc[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28764_ (.CLK(clock),
    .D(_01777_),
    .Q(\fetch.bht.bhtTable_target_pc[5][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28765_ (.CLK(clock),
    .D(_01778_),
    .Q(\fetch.bht.bhtTable_target_pc[5][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28766_ (.CLK(clock),
    .D(_01779_),
    .Q(\fetch.bht.bhtTable_target_pc[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28767_ (.CLK(clock),
    .D(_01780_),
    .Q(\fetch.bht.bhtTable_target_pc[5][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28768_ (.CLK(clock),
    .D(_01781_),
    .Q(\fetch.bht.bhtTable_target_pc[5][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28769_ (.CLK(clock),
    .D(_01782_),
    .Q(\fetch.bht.bhtTable_target_pc[5][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28770_ (.CLK(clock),
    .D(_01783_),
    .Q(\fetch.bht.bhtTable_target_pc[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28771_ (.CLK(clock),
    .D(_01784_),
    .Q(\fetch.bht.bhtTable_target_pc[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28772_ (.CLK(clock),
    .D(_01785_),
    .Q(\fetch.bht.bhtTable_target_pc[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28773_ (.CLK(clock),
    .D(_01786_),
    .Q(\fetch.bht.bhtTable_target_pc[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28774_ (.CLK(clock),
    .D(_01787_),
    .Q(\fetch.bht.bhtTable_target_pc[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28775_ (.CLK(clock),
    .D(_01788_),
    .Q(\fetch.bht.bhtTable_target_pc[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28776_ (.CLK(clock),
    .D(_01789_),
    .Q(\fetch.bht.bhtTable_target_pc[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28777_ (.CLK(clock),
    .D(_01790_),
    .Q(\fetch.bht.bhtTable_target_pc[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28778_ (.CLK(clock),
    .D(_01791_),
    .Q(\fetch.bht.bhtTable_target_pc[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28779_ (.CLK(clock),
    .D(_01792_),
    .Q(\fetch.bht.bhtTable_target_pc[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28780_ (.CLK(clock),
    .D(_01793_),
    .Q(\fetch.bht.bhtTable_target_pc[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28781_ (.CLK(clock),
    .D(_01794_),
    .Q(\fetch.bht.bhtTable_target_pc[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28782_ (.CLK(clock),
    .D(_01795_),
    .Q(\fetch.bht.bhtTable_target_pc[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28783_ (.CLK(clock),
    .D(_01796_),
    .Q(\fetch.bht.bhtTable_target_pc[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28784_ (.CLK(clock),
    .D(_01797_),
    .Q(\fetch.bht.bhtTable_target_pc[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28785_ (.CLK(clock),
    .D(_01798_),
    .Q(\fetch.bht.bhtTable_target_pc[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28786_ (.CLK(clock),
    .D(_01799_),
    .Q(\fetch.bht.bhtTable_target_pc[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28787_ (.CLK(clock),
    .D(_01800_),
    .Q(\fetch.bht.bhtTable_target_pc[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28788_ (.CLK(clock),
    .D(_01801_),
    .Q(\fetch.bht.bhtTable_target_pc[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28789_ (.CLK(clock),
    .D(_01802_),
    .Q(\fetch.bht.bhtTable_target_pc[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28790_ (.CLK(clock),
    .D(_01803_),
    .Q(\fetch.bht.bhtTable_target_pc[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28791_ (.CLK(clock),
    .D(_01804_),
    .Q(\fetch.bht.bhtTable_target_pc[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28792_ (.CLK(clock),
    .D(_01805_),
    .Q(\fetch.bht.bhtTable_target_pc[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28793_ (.CLK(clock),
    .D(_01806_),
    .Q(\fetch.bht.bhtTable_target_pc[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28794_ (.CLK(clock),
    .D(_01807_),
    .Q(\fetch.bht.bhtTable_target_pc[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28795_ (.CLK(clock),
    .D(_01808_),
    .Q(\fetch.bht.bhtTable_target_pc[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28796_ (.CLK(clock),
    .D(_01809_),
    .Q(\fetch.bht.bhtTable_target_pc[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28797_ (.CLK(clock),
    .D(_01810_),
    .Q(\fetch.bht.bhtTable_target_pc[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28798_ (.CLK(clock),
    .D(_01811_),
    .Q(\fetch.bht.bhtTable_target_pc[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28799_ (.CLK(clock),
    .D(_01812_),
    .Q(\fetch.bht.bhtTable_target_pc[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28800_ (.CLK(clock),
    .D(_01813_),
    .Q(\fetch.bht.bhtTable_target_pc[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28801_ (.CLK(clock),
    .D(_01814_),
    .Q(\fetch.bht.bhtTable_target_pc[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28802_ (.CLK(clock),
    .D(_01815_),
    .Q(\fetch.bht.bhtTable_target_pc[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28803_ (.CLK(clock),
    .D(_01816_),
    .Q(\fetch.bht.bhtTable_target_pc[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28804_ (.CLK(clock),
    .D(_01817_),
    .Q(\fetch.bht.bhtTable_target_pc[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28805_ (.CLK(clock),
    .D(_01818_),
    .Q(\fetch.bht.bhtTable_target_pc[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28806_ (.CLK(clock),
    .D(_01819_),
    .Q(\fetch.bht.bhtTable_target_pc[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28807_ (.CLK(clock),
    .D(_01820_),
    .Q(\fetch.bht.bhtTable_target_pc[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28808_ (.CLK(clock),
    .D(_01821_),
    .Q(\fetch.bht.bhtTable_target_pc[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28809_ (.CLK(clock),
    .D(_01822_),
    .Q(\fetch.bht.bhtTable_target_pc[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28810_ (.CLK(clock),
    .D(_01823_),
    .Q(\fetch.bht.bhtTable_target_pc[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28811_ (.CLK(clock),
    .D(_01824_),
    .Q(\fetch.bht.bhtTable_target_pc[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28812_ (.CLK(clock),
    .D(_01825_),
    .Q(\fetch.bht.bhtTable_target_pc[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28813_ (.CLK(clock),
    .D(_01826_),
    .Q(\fetch.bht.bhtTable_target_pc[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28814_ (.CLK(clock),
    .D(_01827_),
    .Q(\fetch.bht.bhtTable_target_pc[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28815_ (.CLK(clock),
    .D(_01828_),
    .Q(\fetch.bht.bhtTable_target_pc[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28816_ (.CLK(clock),
    .D(_01829_),
    .Q(\fetch.bht.bhtTable_target_pc[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28817_ (.CLK(clock),
    .D(_01830_),
    .Q(\fetch.bht.bhtTable_target_pc[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28818_ (.CLK(clock),
    .D(_01831_),
    .Q(\fetch.bht.bhtTable_target_pc[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28819_ (.CLK(clock),
    .D(_01832_),
    .Q(\fetch.bht.bhtTable_target_pc[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28820_ (.CLK(clock),
    .D(_01833_),
    .Q(\fetch.bht.bhtTable_target_pc[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28821_ (.CLK(clock),
    .D(_01834_),
    .Q(\fetch.bht.bhtTable_target_pc[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28822_ (.CLK(clock),
    .D(_01835_),
    .Q(\fetch.bht.bhtTable_target_pc[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28823_ (.CLK(clock),
    .D(_01836_),
    .Q(\fetch.bht.bhtTable_target_pc[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28824_ (.CLK(clock),
    .D(_01837_),
    .Q(\fetch.bht.bhtTable_target_pc[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28825_ (.CLK(clock),
    .D(_01838_),
    .Q(\fetch.bht.bhtTable_target_pc[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28826_ (.CLK(clock),
    .D(_01839_),
    .Q(\fetch.bht.bhtTable_target_pc[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28827_ (.CLK(clock),
    .D(_01840_),
    .Q(\fetch.bht.bhtTable_target_pc[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28828_ (.CLK(clock),
    .D(_01841_),
    .Q(\fetch.bht.bhtTable_target_pc[7][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28829_ (.CLK(clock),
    .D(_01842_),
    .Q(\fetch.bht.bhtTable_target_pc[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28830_ (.CLK(clock),
    .D(_01843_),
    .Q(\fetch.bht.bhtTable_target_pc[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28831_ (.CLK(clock),
    .D(_01844_),
    .Q(\fetch.bht.bhtTable_target_pc[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28832_ (.CLK(clock),
    .D(_01845_),
    .Q(\fetch.bht.bhtTable_target_pc[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28833_ (.CLK(clock),
    .D(_01846_),
    .Q(\fetch.bht.bhtTable_target_pc[7][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28834_ (.CLK(clock),
    .D(_01847_),
    .Q(\fetch.bht.bhtTable_target_pc[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28835_ (.CLK(clock),
    .D(_01848_),
    .Q(\fetch.bht.bhtTable_target_pc[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28836_ (.CLK(clock),
    .D(_01849_),
    .Q(\fetch.bht.bhtTable_target_pc[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28837_ (.CLK(clock),
    .D(_01850_),
    .Q(\fetch.bht.bhtTable_target_pc[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28838_ (.CLK(clock),
    .D(_01851_),
    .Q(\fetch.bht.bhtTable_target_pc[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28839_ (.CLK(clock),
    .D(_01852_),
    .Q(\fetch.bht.bhtTable_target_pc[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28840_ (.CLK(clock),
    .D(_01853_),
    .Q(\fetch.bht.bhtTable_target_pc[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28841_ (.CLK(clock),
    .D(_01854_),
    .Q(\fetch.bht.bhtTable_target_pc[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28842_ (.CLK(clock),
    .D(_01855_),
    .Q(\fetch.bht.bhtTable_target_pc[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28843_ (.CLK(clock),
    .D(_01856_),
    .Q(\fetch.bht.bhtTable_target_pc[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28844_ (.CLK(clock),
    .D(_01857_),
    .Q(\fetch.bht.bhtTable_target_pc[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28845_ (.CLK(clock),
    .D(_01858_),
    .Q(\fetch.bht.bhtTable_target_pc[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28846_ (.CLK(clock),
    .D(_01859_),
    .Q(\fetch.bht.bhtTable_target_pc[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28847_ (.CLK(clock),
    .D(_01860_),
    .Q(\fetch.bht.bhtTable_target_pc[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28848_ (.CLK(clock),
    .D(_01861_),
    .Q(\fetch.bht.bhtTable_target_pc[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28849_ (.CLK(clock),
    .D(_01862_),
    .Q(\fetch.bht.bhtTable_target_pc[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28850_ (.CLK(clock),
    .D(_01863_),
    .Q(\fetch.bht.bhtTable_target_pc[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28851_ (.CLK(clock),
    .D(_01864_),
    .Q(\fetch.bht.bhtTable_target_pc[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28852_ (.CLK(clock),
    .D(_01865_),
    .Q(\fetch.bht.bhtTable_target_pc[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28853_ (.CLK(clock),
    .D(_01866_),
    .Q(\fetch.bht.bhtTable_target_pc[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28854_ (.CLK(clock),
    .D(_01867_),
    .Q(\fetch.bht.bhtTable_target_pc[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28855_ (.CLK(clock),
    .D(_01868_),
    .Q(\fetch.bht.bhtTable_target_pc[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28856_ (.CLK(clock),
    .D(_01869_),
    .Q(\fetch.bht.bhtTable_target_pc[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28857_ (.CLK(clock),
    .D(_01870_),
    .Q(\fetch.bht.bhtTable_target_pc[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28858_ (.CLK(clock),
    .D(_01871_),
    .Q(\fetch.bht.bhtTable_target_pc[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28859_ (.CLK(clock),
    .D(_01872_),
    .Q(\fetch.bht.bhtTable_target_pc[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28860_ (.CLK(clock),
    .D(_01873_),
    .Q(\fetch.bht.bhtTable_target_pc[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28861_ (.CLK(clock),
    .D(_01874_),
    .Q(\fetch.bht.bhtTable_target_pc[8][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28862_ (.CLK(clock),
    .D(_01875_),
    .Q(\fetch.bht.bhtTable_target_pc[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28863_ (.CLK(clock),
    .D(_01876_),
    .Q(\fetch.bht.bhtTable_target_pc[8][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28864_ (.CLK(clock),
    .D(_01877_),
    .Q(\fetch.bht.bhtTable_target_pc[8][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28865_ (.CLK(clock),
    .D(_01878_),
    .Q(\fetch.bht.bhtTable_target_pc[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28866_ (.CLK(clock),
    .D(_01879_),
    .Q(\fetch.bht.bhtTable_target_pc[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28867_ (.CLK(clock),
    .D(_01880_),
    .Q(\fetch.bht.bhtTable_target_pc[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28868_ (.CLK(clock),
    .D(_01881_),
    .Q(\fetch.bht.bhtTable_target_pc[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28869_ (.CLK(clock),
    .D(_01882_),
    .Q(\fetch.bht.bhtTable_target_pc[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28870_ (.CLK(clock),
    .D(_01883_),
    .Q(\fetch.bht.bhtTable_target_pc[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28871_ (.CLK(clock),
    .D(_01884_),
    .Q(\fetch.bht.bhtTable_target_pc[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28872_ (.CLK(clock),
    .D(_01885_),
    .Q(\fetch.bht.bhtTable_target_pc[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28873_ (.CLK(clock),
    .D(_01886_),
    .Q(\fetch.bht.bhtTable_target_pc[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28874_ (.CLK(clock),
    .D(_01887_),
    .Q(\fetch.bht.bhtTable_target_pc[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28875_ (.CLK(clock),
    .D(_01888_),
    .Q(\fetch.bht.bhtTable_target_pc[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28876_ (.CLK(clock),
    .D(_01889_),
    .Q(\fetch.bht.bhtTable_target_pc[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28877_ (.CLK(clock),
    .D(_01890_),
    .Q(\fetch.bht.bhtTable_target_pc[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28878_ (.CLK(clock),
    .D(_01891_),
    .Q(\fetch.bht.bhtTable_target_pc[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28879_ (.CLK(clock),
    .D(_01892_),
    .Q(\fetch.bht.bhtTable_target_pc[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28880_ (.CLK(clock),
    .D(_01893_),
    .Q(\fetch.bht.bhtTable_target_pc[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28881_ (.CLK(clock),
    .D(_01894_),
    .Q(\fetch.bht.bhtTable_target_pc[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28882_ (.CLK(clock),
    .D(_01895_),
    .Q(\fetch.bht.bhtTable_target_pc[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28883_ (.CLK(clock),
    .D(_01896_),
    .Q(\fetch.bht.bhtTable_target_pc[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28884_ (.CLK(clock),
    .D(_01897_),
    .Q(\fetch.bht.bhtTable_target_pc[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28885_ (.CLK(clock),
    .D(_01898_),
    .Q(\fetch.bht.bhtTable_target_pc[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28886_ (.CLK(clock),
    .D(_01899_),
    .Q(\fetch.bht.bhtTable_target_pc[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28887_ (.CLK(clock),
    .D(_01900_),
    .Q(\fetch.bht.bhtTable_target_pc[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28888_ (.CLK(clock),
    .D(_01901_),
    .Q(\fetch.bht.bhtTable_target_pc[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28889_ (.CLK(clock),
    .D(_01902_),
    .Q(\fetch.bht.bhtTable_target_pc[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28890_ (.CLK(clock),
    .D(_01903_),
    .Q(\fetch.bht.bhtTable_target_pc[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28891_ (.CLK(clock),
    .D(_01904_),
    .Q(\fetch.bht.bhtTable_target_pc[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28892_ (.CLK(clock),
    .D(_01905_),
    .Q(\fetch.bht.bhtTable_target_pc[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28893_ (.CLK(clock),
    .D(_01906_),
    .Q(\fetch.bht.bhtTable_target_pc[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28894_ (.CLK(clock),
    .D(_01907_),
    .Q(\fetch.bht.bhtTable_target_pc[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28895_ (.CLK(clock),
    .D(_01908_),
    .Q(\fetch.bht.bhtTable_target_pc[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28896_ (.CLK(clock),
    .D(_01909_),
    .Q(\fetch.bht.bhtTable_target_pc[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28897_ (.CLK(clock),
    .D(_01910_),
    .Q(\fetch.bht.bhtTable_target_pc[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28898_ (.CLK(clock),
    .D(_01911_),
    .Q(\fetch.bht.bhtTable_target_pc[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28899_ (.CLK(clock),
    .D(_01912_),
    .Q(\fetch.bht.bhtTable_target_pc[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28900_ (.CLK(clock),
    .D(_01913_),
    .Q(\fetch.bht.bhtTable_target_pc[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28901_ (.CLK(clock),
    .D(_01914_),
    .Q(\fetch.bht.bhtTable_target_pc[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28902_ (.CLK(clock),
    .D(_01915_),
    .Q(\fetch.bht.bhtTable_target_pc[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28903_ (.CLK(clock),
    .D(_01916_),
    .Q(\fetch.bht.bhtTable_target_pc[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28904_ (.CLK(clock),
    .D(_01917_),
    .Q(\fetch.bht.bhtTable_target_pc[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28905_ (.CLK(clock),
    .D(_01918_),
    .Q(\fetch.bht.bhtTable_target_pc[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28906_ (.CLK(clock),
    .D(_01919_),
    .Q(\fetch.bht.bhtTable_target_pc[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28907_ (.CLK(clock),
    .D(_01920_),
    .Q(\fetch.bht.bhtTable_target_pc[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28908_ (.CLK(clock),
    .D(_01921_),
    .Q(\fetch.bht.bhtTable_target_pc[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28909_ (.CLK(clock),
    .D(_01922_),
    .Q(\fetch.bht.bhtTable_target_pc[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28910_ (.CLK(clock),
    .D(_01923_),
    .Q(\fetch.bht.bhtTable_target_pc[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28911_ (.CLK(clock),
    .D(_01924_),
    .Q(\fetch.bht.bhtTable_target_pc[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28912_ (.CLK(clock),
    .D(_01925_),
    .Q(\fetch.bht.bhtTable_target_pc[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28913_ (.CLK(clock),
    .D(_01926_),
    .Q(\fetch.bht.bhtTable_target_pc[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28914_ (.CLK(clock),
    .D(_01927_),
    .Q(\fetch.bht.bhtTable_target_pc[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28915_ (.CLK(clock),
    .D(_01928_),
    .Q(\fetch.bht.bhtTable_target_pc[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28916_ (.CLK(clock),
    .D(_01929_),
    .Q(\fetch.bht.bhtTable_target_pc[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28917_ (.CLK(clock),
    .D(_01930_),
    .Q(\fetch.bht.bhtTable_target_pc[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28918_ (.CLK(clock),
    .D(_01931_),
    .Q(\fetch.bht.bhtTable_target_pc[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28919_ (.CLK(clock),
    .D(_01932_),
    .Q(\fetch.bht.bhtTable_target_pc[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28920_ (.CLK(clock),
    .D(_01933_),
    .Q(\fetch.bht.bhtTable_target_pc[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28921_ (.CLK(clock),
    .D(_01934_),
    .Q(\fetch.bht.bhtTable_target_pc[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28922_ (.CLK(clock),
    .D(_01935_),
    .Q(\fetch.bht.bhtTable_target_pc[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28923_ (.CLK(clock),
    .D(_01936_),
    .Q(\fetch.bht.bhtTable_target_pc[10][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28924_ (.CLK(clock),
    .D(_01937_),
    .Q(\fetch.bht.bhtTable_target_pc[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28925_ (.CLK(clock),
    .D(_01938_),
    .Q(\fetch.bht.bhtTable_target_pc[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28926_ (.CLK(clock),
    .D(_01939_),
    .Q(\fetch.bht.bhtTable_target_pc[10][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28927_ (.CLK(clock),
    .D(_01940_),
    .Q(\fetch.bht.bhtTable_target_pc[10][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28928_ (.CLK(clock),
    .D(_01941_),
    .Q(\fetch.bht.bhtTable_target_pc[10][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28929_ (.CLK(clock),
    .D(_01942_),
    .Q(\fetch.bht.bhtTable_target_pc[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28930_ (.CLK(clock),
    .D(_01943_),
    .Q(\fetch.bht.bhtTable_target_pc[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28931_ (.CLK(clock),
    .D(_01944_),
    .Q(\fetch.bht.bhtTable_target_pc[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28932_ (.CLK(clock),
    .D(_01945_),
    .Q(\fetch.bht.bhtTable_target_pc[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28933_ (.CLK(clock),
    .D(_01946_),
    .Q(\fetch.bht.bhtTable_target_pc[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28934_ (.CLK(clock),
    .D(_01947_),
    .Q(\fetch.bht.bhtTable_target_pc[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28935_ (.CLK(clock),
    .D(_01948_),
    .Q(\fetch.bht.bhtTable_target_pc[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28936_ (.CLK(clock),
    .D(_01949_),
    .Q(\fetch.bht.bhtTable_target_pc[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28937_ (.CLK(clock),
    .D(_01950_),
    .Q(\fetch.bht.bhtTable_target_pc[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28938_ (.CLK(clock),
    .D(_01951_),
    .Q(\fetch.bht.bhtTable_target_pc[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28939_ (.CLK(clock),
    .D(_01952_),
    .Q(\fetch.bht.bhtTable_target_pc[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28940_ (.CLK(clock),
    .D(_01953_),
    .Q(\fetch.bht.bhtTable_target_pc[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28941_ (.CLK(clock),
    .D(_01954_),
    .Q(\fetch.bht.bhtTable_target_pc[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28942_ (.CLK(clock),
    .D(_01955_),
    .Q(\fetch.bht.bhtTable_target_pc[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28943_ (.CLK(clock),
    .D(_01956_),
    .Q(\fetch.bht.bhtTable_target_pc[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28944_ (.CLK(clock),
    .D(_01957_),
    .Q(\fetch.bht.bhtTable_target_pc[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28945_ (.CLK(clock),
    .D(_01958_),
    .Q(\fetch.bht.bhtTable_target_pc[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28946_ (.CLK(clock),
    .D(_01959_),
    .Q(\fetch.bht.bhtTable_target_pc[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28947_ (.CLK(clock),
    .D(_01960_),
    .Q(\fetch.bht.bhtTable_target_pc[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28948_ (.CLK(clock),
    .D(_01961_),
    .Q(\fetch.bht.bhtTable_target_pc[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28949_ (.CLK(clock),
    .D(_01962_),
    .Q(\fetch.bht.bhtTable_target_pc[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28950_ (.CLK(clock),
    .D(_01963_),
    .Q(\fetch.bht.bhtTable_target_pc[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28951_ (.CLK(clock),
    .D(_01964_),
    .Q(\fetch.bht.bhtTable_target_pc[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28952_ (.CLK(clock),
    .D(_01965_),
    .Q(\fetch.bht.bhtTable_target_pc[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28953_ (.CLK(clock),
    .D(_01966_),
    .Q(\fetch.bht.bhtTable_target_pc[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28954_ (.CLK(clock),
    .D(_01967_),
    .Q(\fetch.bht.bhtTable_target_pc[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28955_ (.CLK(clock),
    .D(_01968_),
    .Q(\fetch.bht.bhtTable_target_pc[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28956_ (.CLK(clock),
    .D(_01969_),
    .Q(\fetch.bht.bhtTable_target_pc[11][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28957_ (.CLK(clock),
    .D(_01970_),
    .Q(\fetch.bht.bhtTable_target_pc[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28958_ (.CLK(clock),
    .D(_01971_),
    .Q(\fetch.bht.bhtTable_target_pc[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28959_ (.CLK(clock),
    .D(_01972_),
    .Q(\fetch.bht.bhtTable_target_pc[11][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28960_ (.CLK(clock),
    .D(_01973_),
    .Q(\fetch.bht.bhtTable_target_pc[11][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28961_ (.CLK(clock),
    .D(_01974_),
    .Q(\fetch.bht.bhtTable_target_pc[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28962_ (.CLK(clock),
    .D(_01975_),
    .Q(\fetch.bht.bhtTable_target_pc[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28963_ (.CLK(clock),
    .D(_01976_),
    .Q(\fetch.bht.bhtTable_target_pc[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28964_ (.CLK(clock),
    .D(_01977_),
    .Q(\fetch.bht.bhtTable_target_pc[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28965_ (.CLK(clock),
    .D(_01978_),
    .Q(\fetch.bht.bhtTable_target_pc[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28966_ (.CLK(clock),
    .D(_01979_),
    .Q(\fetch.bht.bhtTable_target_pc[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28967_ (.CLK(clock),
    .D(_01980_),
    .Q(\fetch.bht.bhtTable_target_pc[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _28968_ (.CLK(clock),
    .D(_01981_),
    .Q(\fetch.bht.bhtTable_target_pc[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _28969_ (.CLK(clock),
    .D(_01982_),
    .Q(\fetch.bht.bhtTable_target_pc[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _28970_ (.CLK(clock),
    .D(_01983_),
    .Q(\fetch.bht.bhtTable_target_pc[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _28971_ (.CLK(clock),
    .D(_01984_),
    .Q(\fetch.bht.bhtTable_target_pc[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _28972_ (.CLK(clock),
    .D(_01985_),
    .Q(\fetch.bht.bhtTable_target_pc[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _28973_ (.CLK(clock),
    .D(_01986_),
    .Q(\fetch.bht.bhtTable_target_pc[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _28974_ (.CLK(clock),
    .D(_01987_),
    .Q(\fetch.bht.bhtTable_target_pc[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _28975_ (.CLK(clock),
    .D(_01988_),
    .Q(\fetch.bht.bhtTable_target_pc[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _28976_ (.CLK(clock),
    .D(_01989_),
    .Q(\fetch.bht.bhtTable_target_pc[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _28977_ (.CLK(clock),
    .D(_01990_),
    .Q(\fetch.bht.bhtTable_target_pc[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _28978_ (.CLK(clock),
    .D(_01991_),
    .Q(\fetch.bht.bhtTable_target_pc[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _28979_ (.CLK(clock),
    .D(_01992_),
    .Q(\fetch.bht.bhtTable_target_pc[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _28980_ (.CLK(clock),
    .D(_01993_),
    .Q(\fetch.bht.bhtTable_target_pc[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _28981_ (.CLK(clock),
    .D(_01994_),
    .Q(\fetch.bht.bhtTable_target_pc[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _28982_ (.CLK(clock),
    .D(_01995_),
    .Q(\fetch.bht.bhtTable_target_pc[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _28983_ (.CLK(clock),
    .D(_01996_),
    .Q(\fetch.bht.bhtTable_target_pc[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _28984_ (.CLK(clock),
    .D(_01997_),
    .Q(\fetch.bht.bhtTable_target_pc[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _28985_ (.CLK(clock),
    .D(_01998_),
    .Q(\fetch.bht.bhtTable_target_pc[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _28986_ (.CLK(clock),
    .D(_01999_),
    .Q(\fetch.bht.bhtTable_target_pc[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _28987_ (.CLK(clock),
    .D(_02000_),
    .Q(\fetch.bht.bhtTable_target_pc[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 _28988_ (.CLK(clock),
    .D(_02001_),
    .Q(\fetch.bht.bhtTable_target_pc[12][26] ));
 sky130_fd_sc_hd__dfxtp_2 _28989_ (.CLK(clock),
    .D(_02002_),
    .Q(\fetch.bht.bhtTable_target_pc[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 _28990_ (.CLK(clock),
    .D(_02003_),
    .Q(\fetch.bht.bhtTable_target_pc[12][28] ));
 sky130_fd_sc_hd__dfxtp_2 _28991_ (.CLK(clock),
    .D(_02004_),
    .Q(\fetch.bht.bhtTable_target_pc[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 _28992_ (.CLK(clock),
    .D(_02005_),
    .Q(\fetch.bht.bhtTable_target_pc[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 _28993_ (.CLK(clock),
    .D(_02006_),
    .Q(\fetch.bht.bhtTable_target_pc[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 _28994_ (.CLK(clock),
    .D(_02007_),
    .Q(\fetch.bht.bhtTable_target_pc[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _28995_ (.CLK(clock),
    .D(_02008_),
    .Q(\fetch.bht.bhtTable_target_pc[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _28996_ (.CLK(clock),
    .D(_02009_),
    .Q(\fetch.bht.bhtTable_target_pc[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _28997_ (.CLK(clock),
    .D(_02010_),
    .Q(\fetch.bht.bhtTable_target_pc[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _28998_ (.CLK(clock),
    .D(_02011_),
    .Q(\fetch.bht.bhtTable_target_pc[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _28999_ (.CLK(clock),
    .D(_02012_),
    .Q(\fetch.bht.bhtTable_target_pc[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _29000_ (.CLK(clock),
    .D(_02013_),
    .Q(\fetch.bht.bhtTable_target_pc[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _29001_ (.CLK(clock),
    .D(_02014_),
    .Q(\fetch.bht.bhtTable_target_pc[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _29002_ (.CLK(clock),
    .D(_02015_),
    .Q(\fetch.bht.bhtTable_target_pc[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _29003_ (.CLK(clock),
    .D(_02016_),
    .Q(\fetch.bht.bhtTable_target_pc[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _29004_ (.CLK(clock),
    .D(_02017_),
    .Q(\fetch.bht.bhtTable_target_pc[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _29005_ (.CLK(clock),
    .D(_02018_),
    .Q(\fetch.bht.bhtTable_target_pc[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _29006_ (.CLK(clock),
    .D(_02019_),
    .Q(\fetch.bht.bhtTable_target_pc[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _29007_ (.CLK(clock),
    .D(_02020_),
    .Q(\fetch.bht.bhtTable_target_pc[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _29008_ (.CLK(clock),
    .D(_02021_),
    .Q(\fetch.bht.bhtTable_target_pc[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _29009_ (.CLK(clock),
    .D(_02022_),
    .Q(\fetch.bht.bhtTable_target_pc[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _29010_ (.CLK(clock),
    .D(_02023_),
    .Q(\fetch.bht.bhtTable_target_pc[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _29011_ (.CLK(clock),
    .D(_02024_),
    .Q(\fetch.bht.bhtTable_target_pc[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _29012_ (.CLK(clock),
    .D(_02025_),
    .Q(\fetch.bht.bhtTable_target_pc[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _29013_ (.CLK(clock),
    .D(_02026_),
    .Q(\fetch.bht.bhtTable_target_pc[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _29014_ (.CLK(clock),
    .D(_02027_),
    .Q(\fetch.bht.bhtTable_target_pc[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _29015_ (.CLK(clock),
    .D(_02028_),
    .Q(\fetch.bht.bhtTable_target_pc[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _29016_ (.CLK(clock),
    .D(_02029_),
    .Q(\fetch.bht.bhtTable_target_pc[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _29017_ (.CLK(clock),
    .D(_02030_),
    .Q(\fetch.bht.bhtTable_target_pc[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _29018_ (.CLK(clock),
    .D(_02031_),
    .Q(\fetch.bht.bhtTable_target_pc[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _29019_ (.CLK(clock),
    .D(_02032_),
    .Q(\fetch.bht.bhtTable_target_pc[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 _29020_ (.CLK(clock),
    .D(_02033_),
    .Q(\fetch.bht.bhtTable_target_pc[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 _29021_ (.CLK(clock),
    .D(_02034_),
    .Q(\fetch.bht.bhtTable_target_pc[13][27] ));
 sky130_fd_sc_hd__dfxtp_2 _29022_ (.CLK(clock),
    .D(_02035_),
    .Q(\fetch.bht.bhtTable_target_pc[13][28] ));
 sky130_fd_sc_hd__dfxtp_2 _29023_ (.CLK(clock),
    .D(_02036_),
    .Q(\fetch.bht.bhtTable_target_pc[13][29] ));
 sky130_fd_sc_hd__dfxtp_2 _29024_ (.CLK(clock),
    .D(_02037_),
    .Q(\fetch.bht.bhtTable_target_pc[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 _29025_ (.CLK(clock),
    .D(_02038_),
    .Q(\fetch.bht.bhtTable_target_pc[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _29026_ (.CLK(clock),
    .D(_02039_),
    .Q(\fetch.bht.bhtTable_target_pc[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29027_ (.CLK(clock),
    .D(_02040_),
    .Q(\fetch.bht.bhtTable_target_pc[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29028_ (.CLK(clock),
    .D(_02041_),
    .Q(\fetch.bht.bhtTable_target_pc[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _29029_ (.CLK(clock),
    .D(_02042_),
    .Q(\fetch.bht.bhtTable_target_pc[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _29030_ (.CLK(clock),
    .D(_02043_),
    .Q(\fetch.bht.bhtTable_target_pc[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _29031_ (.CLK(clock),
    .D(_02044_),
    .Q(\fetch.bht.bhtTable_target_pc[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _29032_ (.CLK(clock),
    .D(_02045_),
    .Q(\fetch.bht.bhtTable_target_pc[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _29033_ (.CLK(clock),
    .D(_02046_),
    .Q(\fetch.bht.bhtTable_target_pc[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _29034_ (.CLK(clock),
    .D(_02047_),
    .Q(\fetch.bht.bhtTable_target_pc[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _29035_ (.CLK(clock),
    .D(_02048_),
    .Q(\fetch.bht.bhtTable_target_pc[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _29036_ (.CLK(clock),
    .D(_02049_),
    .Q(\fetch.bht.bhtTable_target_pc[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _29037_ (.CLK(clock),
    .D(_02050_),
    .Q(\fetch.bht.bhtTable_target_pc[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _29038_ (.CLK(clock),
    .D(_02051_),
    .Q(\fetch.bht.bhtTable_target_pc[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _29039_ (.CLK(clock),
    .D(_02052_),
    .Q(\fetch.bht.bhtTable_target_pc[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _29040_ (.CLK(clock),
    .D(_02053_),
    .Q(\fetch.bht.bhtTable_target_pc[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _29041_ (.CLK(clock),
    .D(_02054_),
    .Q(\fetch.bht.bhtTable_target_pc[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _29042_ (.CLK(clock),
    .D(_02055_),
    .Q(\fetch.bht.bhtTable_target_pc[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _29043_ (.CLK(clock),
    .D(_02056_),
    .Q(\fetch.bht.bhtTable_target_pc[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _29044_ (.CLK(clock),
    .D(_02057_),
    .Q(\fetch.bht.bhtTable_target_pc[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _29045_ (.CLK(clock),
    .D(_02058_),
    .Q(\fetch.bht.bhtTable_target_pc[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _29046_ (.CLK(clock),
    .D(_02059_),
    .Q(\fetch.bht.bhtTable_target_pc[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _29047_ (.CLK(clock),
    .D(_02060_),
    .Q(\fetch.bht.bhtTable_target_pc[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _29048_ (.CLK(clock),
    .D(_02061_),
    .Q(\fetch.bht.bhtTable_target_pc[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _29049_ (.CLK(clock),
    .D(_02062_),
    .Q(\fetch.bht.bhtTable_target_pc[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _29050_ (.CLK(clock),
    .D(_02063_),
    .Q(\fetch.bht.bhtTable_target_pc[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _29051_ (.CLK(clock),
    .D(_02064_),
    .Q(\fetch.bht.bhtTable_target_pc[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _29052_ (.CLK(clock),
    .D(_02065_),
    .Q(\fetch.bht.bhtTable_target_pc[14][26] ));
 sky130_fd_sc_hd__dfxtp_2 _29053_ (.CLK(clock),
    .D(_02066_),
    .Q(\fetch.bht.bhtTable_target_pc[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 _29054_ (.CLK(clock),
    .D(_02067_),
    .Q(\fetch.bht.bhtTable_target_pc[14][28] ));
 sky130_fd_sc_hd__dfxtp_2 _29055_ (.CLK(clock),
    .D(_02068_),
    .Q(\fetch.bht.bhtTable_target_pc[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 _29056_ (.CLK(clock),
    .D(_02069_),
    .Q(\fetch.bht.bhtTable_target_pc[14][30] ));
 sky130_fd_sc_hd__dfxtp_2 _29057_ (.CLK(clock),
    .D(_02070_),
    .Q(\fetch.bht.bhtTable_target_pc[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 _29058_ (.CLK(clock),
    .D(_02071_),
    .Q(\fetch.bht.bhtTable_tag[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29059_ (.CLK(clock),
    .D(_02072_),
    .Q(\fetch.bht.bhtTable_tag[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29060_ (.CLK(clock),
    .D(_02073_),
    .Q(\fetch.bht.bhtTable_tag[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _29061_ (.CLK(clock),
    .D(_02074_),
    .Q(\fetch.bht.bhtTable_tag[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _29062_ (.CLK(clock),
    .D(_02075_),
    .Q(\fetch.bht.bhtTable_tag[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _29063_ (.CLK(clock),
    .D(_02076_),
    .Q(\fetch.bht.bhtTable_tag[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _29064_ (.CLK(clock),
    .D(_02077_),
    .Q(\fetch.bht.bhtTable_tag[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _29065_ (.CLK(clock),
    .D(_02078_),
    .Q(\fetch.bht.bhtTable_tag[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _29066_ (.CLK(clock),
    .D(_02079_),
    .Q(\fetch.bht.bhtTable_tag[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _29067_ (.CLK(clock),
    .D(_02080_),
    .Q(\fetch.bht.bhtTable_tag[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _29068_ (.CLK(clock),
    .D(_02081_),
    .Q(\fetch.bht.bhtTable_tag[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _29069_ (.CLK(clock),
    .D(_02082_),
    .Q(\fetch.bht.bhtTable_tag[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _29070_ (.CLK(clock),
    .D(_02083_),
    .Q(\fetch.bht.bhtTable_tag[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _29071_ (.CLK(clock),
    .D(_02084_),
    .Q(\fetch.bht.bhtTable_tag[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _29072_ (.CLK(clock),
    .D(_02085_),
    .Q(\fetch.bht.bhtTable_tag[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _29073_ (.CLK(clock),
    .D(_02086_),
    .Q(\fetch.bht.bhtTable_tag[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _29074_ (.CLK(clock),
    .D(_02087_),
    .Q(\fetch.bht.bhtTable_tag[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _29075_ (.CLK(clock),
    .D(_02088_),
    .Q(\fetch.bht.bhtTable_tag[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _29076_ (.CLK(clock),
    .D(_02089_),
    .Q(\fetch.bht.bhtTable_tag[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _29077_ (.CLK(clock),
    .D(_02090_),
    .Q(\fetch.bht.bhtTable_tag[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _29078_ (.CLK(clock),
    .D(_02091_),
    .Q(\fetch.bht.bhtTable_tag[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _29079_ (.CLK(clock),
    .D(_02092_),
    .Q(\fetch.bht.bhtTable_tag[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _29080_ (.CLK(clock),
    .D(_02093_),
    .Q(\fetch.bht.bhtTable_tag[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _29081_ (.CLK(clock),
    .D(_02094_),
    .Q(\fetch.bht.bhtTable_tag[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _29082_ (.CLK(clock),
    .D(_02095_),
    .Q(\fetch.bht.bhtTable_tag[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _29083_ (.CLK(clock),
    .D(_02096_),
    .Q(\fetch.bht.bhtTable_tag[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _29084_ (.CLK(clock),
    .D(_02097_),
    .Q(\csr._mcycle_T_3[32] ));
 sky130_fd_sc_hd__dfxtp_2 _29085_ (.CLK(clock),
    .D(_02098_),
    .Q(\csr._mcycle_T_3[33] ));
 sky130_fd_sc_hd__dfxtp_2 _29086_ (.CLK(clock),
    .D(_02099_),
    .Q(\csr._mcycle_T_3[34] ));
 sky130_fd_sc_hd__dfxtp_2 _29087_ (.CLK(clock),
    .D(_02100_),
    .Q(\csr._mcycle_T_3[35] ));
 sky130_fd_sc_hd__dfxtp_2 _29088_ (.CLK(clock),
    .D(_02101_),
    .Q(\csr._mcycle_T_3[36] ));
 sky130_fd_sc_hd__dfxtp_2 _29089_ (.CLK(clock),
    .D(_02102_),
    .Q(\csr._mcycle_T_3[37] ));
 sky130_fd_sc_hd__dfxtp_2 _29090_ (.CLK(clock),
    .D(_02103_),
    .Q(\csr._mcycle_T_3[38] ));
 sky130_fd_sc_hd__dfxtp_2 _29091_ (.CLK(clock),
    .D(_02104_),
    .Q(\csr._mcycle_T_3[39] ));
 sky130_fd_sc_hd__dfxtp_2 _29092_ (.CLK(clock),
    .D(_02105_),
    .Q(\csr._mcycle_T_3[40] ));
 sky130_fd_sc_hd__dfxtp_2 _29093_ (.CLK(clock),
    .D(_02106_),
    .Q(\csr._mcycle_T_3[41] ));
 sky130_fd_sc_hd__dfxtp_2 _29094_ (.CLK(clock),
    .D(_02107_),
    .Q(\csr._mcycle_T_3[42] ));
 sky130_fd_sc_hd__dfxtp_2 _29095_ (.CLK(clock),
    .D(_02108_),
    .Q(\csr._mcycle_T_3[43] ));
 sky130_fd_sc_hd__dfxtp_2 _29096_ (.CLK(clock),
    .D(_02109_),
    .Q(\csr._mcycle_T_3[44] ));
 sky130_fd_sc_hd__dfxtp_2 _29097_ (.CLK(clock),
    .D(_02110_),
    .Q(\csr._mcycle_T_3[45] ));
 sky130_fd_sc_hd__dfxtp_2 _29098_ (.CLK(clock),
    .D(_02111_),
    .Q(\csr._mcycle_T_3[46] ));
 sky130_fd_sc_hd__dfxtp_2 _29099_ (.CLK(clock),
    .D(_02112_),
    .Q(\csr._mcycle_T_3[47] ));
 sky130_fd_sc_hd__dfxtp_2 _29100_ (.CLK(clock),
    .D(_02113_),
    .Q(\csr._mcycle_T_3[48] ));
 sky130_fd_sc_hd__dfxtp_2 _29101_ (.CLK(clock),
    .D(_02114_),
    .Q(\csr._mcycle_T_3[49] ));
 sky130_fd_sc_hd__dfxtp_2 _29102_ (.CLK(clock),
    .D(_02115_),
    .Q(\csr._mcycle_T_3[50] ));
 sky130_fd_sc_hd__dfxtp_2 _29103_ (.CLK(clock),
    .D(_02116_),
    .Q(\csr._mcycle_T_3[51] ));
 sky130_fd_sc_hd__dfxtp_2 _29104_ (.CLK(clock),
    .D(_02117_),
    .Q(\csr._mcycle_T_3[52] ));
 sky130_fd_sc_hd__dfxtp_2 _29105_ (.CLK(clock),
    .D(_02118_),
    .Q(\csr._mcycle_T_3[53] ));
 sky130_fd_sc_hd__dfxtp_2 _29106_ (.CLK(clock),
    .D(_02119_),
    .Q(\csr._mcycle_T_3[54] ));
 sky130_fd_sc_hd__dfxtp_2 _29107_ (.CLK(clock),
    .D(_02120_),
    .Q(\csr._mcycle_T_3[55] ));
 sky130_fd_sc_hd__dfxtp_2 _29108_ (.CLK(clock),
    .D(_02121_),
    .Q(\csr._mcycle_T_3[56] ));
 sky130_fd_sc_hd__dfxtp_2 _29109_ (.CLK(clock),
    .D(_02122_),
    .Q(\csr._mcycle_T_3[57] ));
 sky130_fd_sc_hd__dfxtp_2 _29110_ (.CLK(clock),
    .D(_02123_),
    .Q(\csr._mcycle_T_3[58] ));
 sky130_fd_sc_hd__dfxtp_2 _29111_ (.CLK(clock),
    .D(_02124_),
    .Q(\csr._mcycle_T_3[59] ));
 sky130_fd_sc_hd__dfxtp_2 _29112_ (.CLK(clock),
    .D(_02125_),
    .Q(\csr._mcycle_T_3[60] ));
 sky130_fd_sc_hd__dfxtp_2 _29113_ (.CLK(clock),
    .D(_02126_),
    .Q(\csr._mcycle_T_3[61] ));
 sky130_fd_sc_hd__dfxtp_2 _29114_ (.CLK(clock),
    .D(_02127_),
    .Q(\csr._mcycle_T_3[62] ));
 sky130_fd_sc_hd__dfxtp_2 _29115_ (.CLK(clock),
    .D(_02128_),
    .Q(\csr._mcycle_T_3[63] ));
 sky130_fd_sc_hd__dfxtp_2 _29116_ (.CLK(clock),
    .D(_02129_),
    .Q(\csr.mcycle[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29117_ (.CLK(clock),
    .D(_02130_),
    .Q(\csr.mcycle[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29118_ (.CLK(clock),
    .D(_02131_),
    .Q(\csr.mcycle[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29119_ (.CLK(clock),
    .D(_02132_),
    .Q(\csr.mcycle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29120_ (.CLK(clock),
    .D(_02133_),
    .Q(\csr.mcycle[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29121_ (.CLK(clock),
    .D(_02134_),
    .Q(\csr.mcycle[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29122_ (.CLK(clock),
    .D(_02135_),
    .Q(\csr.mcycle[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29123_ (.CLK(clock),
    .D(_02136_),
    .Q(\csr.mcycle[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29124_ (.CLK(clock),
    .D(_02137_),
    .Q(\csr.mcycle[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29125_ (.CLK(clock),
    .D(_02138_),
    .Q(\csr.mcycle[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29126_ (.CLK(clock),
    .D(_02139_),
    .Q(\csr.mcycle[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29127_ (.CLK(clock),
    .D(_02140_),
    .Q(\csr.mcycle[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29128_ (.CLK(clock),
    .D(_02141_),
    .Q(\csr.mcycle[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29129_ (.CLK(clock),
    .D(_02142_),
    .Q(\csr.mcycle[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29130_ (.CLK(clock),
    .D(_02143_),
    .Q(\csr.mcycle[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29131_ (.CLK(clock),
    .D(_02144_),
    .Q(\csr.mcycle[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29132_ (.CLK(clock),
    .D(_02145_),
    .Q(\csr.mcycle[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29133_ (.CLK(clock),
    .D(_02146_),
    .Q(\csr.mcycle[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29134_ (.CLK(clock),
    .D(_02147_),
    .Q(\csr.mcycle[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29135_ (.CLK(clock),
    .D(_02148_),
    .Q(\csr.mcycle[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29136_ (.CLK(clock),
    .D(_02149_),
    .Q(\csr.mcycle[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29137_ (.CLK(clock),
    .D(_02150_),
    .Q(\csr.mcycle[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29138_ (.CLK(clock),
    .D(_02151_),
    .Q(\csr.mcycle[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29139_ (.CLK(clock),
    .D(_02152_),
    .Q(\csr.mcycle[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29140_ (.CLK(clock),
    .D(_02153_),
    .Q(\csr.mcycle[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29141_ (.CLK(clock),
    .D(_02154_),
    .Q(\csr.mcycle[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29142_ (.CLK(clock),
    .D(_02155_),
    .Q(\csr.mcycle[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29143_ (.CLK(clock),
    .D(_02156_),
    .Q(\csr.mcycle[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29144_ (.CLK(clock),
    .D(_02157_),
    .Q(\csr.mcycle[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29145_ (.CLK(clock),
    .D(_02158_),
    .Q(\csr.mcycle[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29146_ (.CLK(clock),
    .D(_02159_),
    .Q(\csr.mcycle[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29147_ (.CLK(clock),
    .D(_02160_),
    .Q(\csr.mcycle[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29148_ (.CLK(clock),
    .D(_02161_),
    .Q(\fetch.bht.bhtTable_tag[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29149_ (.CLK(clock),
    .D(_02162_),
    .Q(\fetch.bht.bhtTable_tag[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29150_ (.CLK(clock),
    .D(_02163_),
    .Q(\fetch.bht.bhtTable_tag[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _29151_ (.CLK(clock),
    .D(_02164_),
    .Q(\fetch.bht.bhtTable_tag[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _29152_ (.CLK(clock),
    .D(_02165_),
    .Q(\fetch.bht.bhtTable_tag[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _29153_ (.CLK(clock),
    .D(_02166_),
    .Q(\fetch.bht.bhtTable_tag[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _29154_ (.CLK(clock),
    .D(_02167_),
    .Q(\fetch.bht.bhtTable_tag[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _29155_ (.CLK(clock),
    .D(_02168_),
    .Q(\fetch.bht.bhtTable_tag[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _29156_ (.CLK(clock),
    .D(_02169_),
    .Q(\fetch.bht.bhtTable_tag[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _29157_ (.CLK(clock),
    .D(_02170_),
    .Q(\fetch.bht.bhtTable_tag[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _29158_ (.CLK(clock),
    .D(_02171_),
    .Q(\fetch.bht.bhtTable_tag[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _29159_ (.CLK(clock),
    .D(_02172_),
    .Q(\fetch.bht.bhtTable_tag[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _29160_ (.CLK(clock),
    .D(_02173_),
    .Q(\fetch.bht.bhtTable_tag[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _29161_ (.CLK(clock),
    .D(_02174_),
    .Q(\fetch.bht.bhtTable_tag[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _29162_ (.CLK(clock),
    .D(_02175_),
    .Q(\fetch.bht.bhtTable_tag[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _29163_ (.CLK(clock),
    .D(_02176_),
    .Q(\fetch.bht.bhtTable_tag[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _29164_ (.CLK(clock),
    .D(_02177_),
    .Q(\fetch.bht.bhtTable_tag[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _29165_ (.CLK(clock),
    .D(_02178_),
    .Q(\fetch.bht.bhtTable_tag[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _29166_ (.CLK(clock),
    .D(_02179_),
    .Q(\fetch.bht.bhtTable_tag[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _29167_ (.CLK(clock),
    .D(_02180_),
    .Q(\fetch.bht.bhtTable_tag[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _29168_ (.CLK(clock),
    .D(_02181_),
    .Q(\fetch.bht.bhtTable_tag[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _29169_ (.CLK(clock),
    .D(_02182_),
    .Q(\fetch.bht.bhtTable_tag[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _29170_ (.CLK(clock),
    .D(_02183_),
    .Q(\fetch.bht.bhtTable_tag[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _29171_ (.CLK(clock),
    .D(_02184_),
    .Q(\fetch.bht.bhtTable_tag[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _29172_ (.CLK(clock),
    .D(_02185_),
    .Q(\fetch.bht.bhtTable_tag[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _29173_ (.CLK(clock),
    .D(_02186_),
    .Q(\fetch.bht.bhtTable_tag[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _29174_ (.CLK(clock),
    .D(_02187_),
    .Q(\decode.id_ex_aluop_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29175_ (.CLK(clock),
    .D(_02188_),
    .Q(\decode.id_ex_aluop_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29176_ (.CLK(clock),
    .D(_02189_),
    .Q(_00000_));
 sky130_fd_sc_hd__dfxtp_2 _29177_ (.CLK(clock),
    .D(_02190_),
    .Q(_00001_));
 sky130_fd_sc_hd__dfxtp_2 _29178_ (.CLK(clock),
    .D(_02191_),
    .Q(_00002_));
 sky130_fd_sc_hd__dfxtp_2 _29179_ (.CLK(clock),
    .D(_02192_),
    .Q(_00003_));
 sky130_fd_sc_hd__dfxtp_2 _29180_ (.CLK(clock),
    .D(_02193_),
    .Q(\fetch.btb.btbTable[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29181_ (.CLK(clock),
    .D(_02194_),
    .Q(\fetch.btb.btbTable[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29182_ (.CLK(clock),
    .D(_02195_),
    .Q(\fetch.btb.btbTable[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29183_ (.CLK(clock),
    .D(_02196_),
    .Q(\fetch.btb.btbTable[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29184_ (.CLK(clock),
    .D(_02197_),
    .Q(\fetch.btb.btbTable[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29185_ (.CLK(clock),
    .D(_02198_),
    .Q(\fetch.btb.btbTable[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29186_ (.CLK(clock),
    .D(_02199_),
    .Q(\fetch.btb.btbTable[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29187_ (.CLK(clock),
    .D(_02200_),
    .Q(\fetch.btb.btbTable[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29188_ (.CLK(clock),
    .D(_02201_),
    .Q(\fetch.btb.btbTable[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29189_ (.CLK(clock),
    .D(_02202_),
    .Q(\fetch.btb.btbTable[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29190_ (.CLK(clock),
    .D(_02203_),
    .Q(\fetch.btb.btbTable[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29191_ (.CLK(clock),
    .D(_02204_),
    .Q(\fetch.btb.btbTable[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29192_ (.CLK(clock),
    .D(_02205_),
    .Q(\fetch.btb.btbTable[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29193_ (.CLK(clock),
    .D(_02206_),
    .Q(\fetch.btb.btbTable[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29194_ (.CLK(clock),
    .D(_02207_),
    .Q(\fetch.btb.btbTable[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29195_ (.CLK(clock),
    .D(_02208_),
    .Q(\fetch.btb.btbTable[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29196_ (.CLK(clock),
    .D(_02209_),
    .Q(\fetch.btb.btbTable[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29197_ (.CLK(clock),
    .D(_02210_),
    .Q(\fetch.btb.btbTable[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29198_ (.CLK(clock),
    .D(_02211_),
    .Q(\fetch.btb.btbTable[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29199_ (.CLK(clock),
    .D(_02212_),
    .Q(\fetch.btb.btbTable[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29200_ (.CLK(clock),
    .D(_02213_),
    .Q(\fetch.btb.btbTable[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29201_ (.CLK(clock),
    .D(_02214_),
    .Q(\fetch.btb.btbTable[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29202_ (.CLK(clock),
    .D(_02215_),
    .Q(\fetch.btb.btbTable[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29203_ (.CLK(clock),
    .D(_02216_),
    .Q(\fetch.btb.btbTable[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29204_ (.CLK(clock),
    .D(_02217_),
    .Q(\fetch.btb.btbTable[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29205_ (.CLK(clock),
    .D(_02218_),
    .Q(\fetch.btb.btbTable[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29206_ (.CLK(clock),
    .D(_02219_),
    .Q(\fetch.btb.btbTable[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29207_ (.CLK(clock),
    .D(_02220_),
    .Q(\fetch.btb.btbTable[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29208_ (.CLK(clock),
    .D(_02221_),
    .Q(\fetch.btb.btbTable[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29209_ (.CLK(clock),
    .D(_02222_),
    .Q(\fetch.btb.btbTable[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29210_ (.CLK(clock),
    .D(_02223_),
    .Q(\fetch.bht.bhtTable_target_pc[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _29211_ (.CLK(clock),
    .D(_02224_),
    .Q(\fetch.bht.bhtTable_target_pc[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _29212_ (.CLK(clock),
    .D(_02225_),
    .Q(\fetch.bht.bhtTable_target_pc[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _29213_ (.CLK(clock),
    .D(_02226_),
    .Q(\fetch.bht.bhtTable_target_pc[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _29214_ (.CLK(clock),
    .D(_02227_),
    .Q(\fetch.bht.bhtTable_target_pc[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _29215_ (.CLK(clock),
    .D(_02228_),
    .Q(\fetch.bht.bhtTable_target_pc[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _29216_ (.CLK(clock),
    .D(_02229_),
    .Q(\fetch.bht.bhtTable_target_pc[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _29217_ (.CLK(clock),
    .D(_02230_),
    .Q(\fetch.bht.bhtTable_target_pc[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _29218_ (.CLK(clock),
    .D(_02231_),
    .Q(\fetch.bht.bhtTable_target_pc[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _29219_ (.CLK(clock),
    .D(_02232_),
    .Q(\fetch.bht.bhtTable_target_pc[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _29220_ (.CLK(clock),
    .D(_02233_),
    .Q(\fetch.bht.bhtTable_target_pc[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _29221_ (.CLK(clock),
    .D(_02234_),
    .Q(\fetch.bht.bhtTable_target_pc[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _29222_ (.CLK(clock),
    .D(_02235_),
    .Q(\fetch.bht.bhtTable_target_pc[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _29223_ (.CLK(clock),
    .D(_02236_),
    .Q(\fetch.bht.bhtTable_target_pc[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _29224_ (.CLK(clock),
    .D(_02237_),
    .Q(\fetch.bht.bhtTable_target_pc[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _29225_ (.CLK(clock),
    .D(_02238_),
    .Q(\fetch.bht.bhtTable_target_pc[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _29226_ (.CLK(clock),
    .D(_02239_),
    .Q(\fetch.bht.bhtTable_target_pc[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _29227_ (.CLK(clock),
    .D(_02240_),
    .Q(\fetch.bht.bhtTable_target_pc[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _29228_ (.CLK(clock),
    .D(_02241_),
    .Q(\fetch.bht.bhtTable_target_pc[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _29229_ (.CLK(clock),
    .D(_02242_),
    .Q(\fetch.bht.bhtTable_target_pc[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _29230_ (.CLK(clock),
    .D(_02243_),
    .Q(\fetch.bht.bhtTable_target_pc[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _29231_ (.CLK(clock),
    .D(_02244_),
    .Q(\fetch.bht.bhtTable_target_pc[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _29232_ (.CLK(clock),
    .D(_02245_),
    .Q(\fetch.bht.bhtTable_target_pc[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _29233_ (.CLK(clock),
    .D(_02246_),
    .Q(\fetch.bht.bhtTable_target_pc[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _29234_ (.CLK(clock),
    .D(_02247_),
    .Q(\fetch.bht.bhtTable_target_pc[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _29235_ (.CLK(clock),
    .D(_02248_),
    .Q(\fetch.bht.bhtTable_target_pc[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 _29236_ (.CLK(clock),
    .D(_02249_),
    .Q(\fetch.bht.bhtTable_target_pc[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 _29237_ (.CLK(clock),
    .D(_02250_),
    .Q(\fetch.bht.bhtTable_target_pc[9][27] ));
 sky130_fd_sc_hd__dfxtp_2 _29238_ (.CLK(clock),
    .D(_02251_),
    .Q(\fetch.bht.bhtTable_target_pc[9][28] ));
 sky130_fd_sc_hd__dfxtp_2 _29239_ (.CLK(clock),
    .D(_02252_),
    .Q(\fetch.bht.bhtTable_target_pc[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 _29240_ (.CLK(clock),
    .D(_02253_),
    .Q(\fetch.bht.bhtTable_target_pc[9][30] ));
 sky130_fd_sc_hd__dfxtp_2 _29241_ (.CLK(clock),
    .D(_02254_),
    .Q(\fetch.bht.bhtTable_target_pc[9][31] ));
 sky130_fd_sc_hd__dfxtp_2 _29242_ (.CLK(clock),
    .D(_02255_),
    .Q(\decode.regfile.registers_0[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29243_ (.CLK(clock),
    .D(_02256_),
    .Q(\decode.regfile.registers_0[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29244_ (.CLK(clock),
    .D(_02257_),
    .Q(\decode.regfile.registers_0[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29245_ (.CLK(clock),
    .D(_02258_),
    .Q(\decode.regfile.registers_0[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29246_ (.CLK(clock),
    .D(_02259_),
    .Q(\decode.regfile.registers_0[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29247_ (.CLK(clock),
    .D(_02260_),
    .Q(\decode.regfile.registers_0[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29248_ (.CLK(clock),
    .D(_02261_),
    .Q(\decode.regfile.registers_0[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29249_ (.CLK(clock),
    .D(_02262_),
    .Q(\decode.regfile.registers_0[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29250_ (.CLK(clock),
    .D(_02263_),
    .Q(\decode.regfile.registers_0[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29251_ (.CLK(clock),
    .D(_02264_),
    .Q(\decode.regfile.registers_0[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29252_ (.CLK(clock),
    .D(_02265_),
    .Q(\decode.regfile.registers_0[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29253_ (.CLK(clock),
    .D(_02266_),
    .Q(\decode.regfile.registers_0[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29254_ (.CLK(clock),
    .D(_02267_),
    .Q(\decode.regfile.registers_0[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29255_ (.CLK(clock),
    .D(_02268_),
    .Q(\decode.regfile.registers_0[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29256_ (.CLK(clock),
    .D(_02269_),
    .Q(\decode.regfile.registers_0[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29257_ (.CLK(clock),
    .D(_02270_),
    .Q(\decode.regfile.registers_0[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29258_ (.CLK(clock),
    .D(_02271_),
    .Q(\decode.regfile.registers_0[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29259_ (.CLK(clock),
    .D(_02272_),
    .Q(\decode.regfile.registers_0[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29260_ (.CLK(clock),
    .D(_02273_),
    .Q(\decode.regfile.registers_0[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29261_ (.CLK(clock),
    .D(_02274_),
    .Q(\decode.regfile.registers_0[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29262_ (.CLK(clock),
    .D(_02275_),
    .Q(\decode.regfile.registers_0[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29263_ (.CLK(clock),
    .D(_02276_),
    .Q(\decode.regfile.registers_0[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29264_ (.CLK(clock),
    .D(_02277_),
    .Q(\decode.regfile.registers_0[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29265_ (.CLK(clock),
    .D(_02278_),
    .Q(\decode.regfile.registers_0[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29266_ (.CLK(clock),
    .D(_02279_),
    .Q(\decode.regfile.registers_0[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29267_ (.CLK(clock),
    .D(_02280_),
    .Q(\decode.regfile.registers_0[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29268_ (.CLK(clock),
    .D(_02281_),
    .Q(\decode.regfile.registers_0[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29269_ (.CLK(clock),
    .D(_02282_),
    .Q(\decode.regfile.registers_0[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29270_ (.CLK(clock),
    .D(_02283_),
    .Q(\decode.regfile.registers_0[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29271_ (.CLK(clock),
    .D(_02284_),
    .Q(\decode.regfile.registers_0[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29272_ (.CLK(clock),
    .D(_02285_),
    .Q(\decode.regfile.registers_0[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29273_ (.CLK(clock),
    .D(_02286_),
    .Q(\decode.regfile.registers_0[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29274_ (.CLK(clock),
    .D(_02287_),
    .Q(\decode.regfile.registers_1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29275_ (.CLK(clock),
    .D(_02288_),
    .Q(\decode.regfile.registers_1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29276_ (.CLK(clock),
    .D(_02289_),
    .Q(\decode.regfile.registers_1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29277_ (.CLK(clock),
    .D(_02290_),
    .Q(\decode.regfile.registers_1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29278_ (.CLK(clock),
    .D(_02291_),
    .Q(\decode.regfile.registers_1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29279_ (.CLK(clock),
    .D(_02292_),
    .Q(\decode.regfile.registers_1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29280_ (.CLK(clock),
    .D(_02293_),
    .Q(\decode.regfile.registers_1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29281_ (.CLK(clock),
    .D(_02294_),
    .Q(\decode.regfile.registers_1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29282_ (.CLK(clock),
    .D(_02295_),
    .Q(\decode.regfile.registers_1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29283_ (.CLK(clock),
    .D(_02296_),
    .Q(\decode.regfile.registers_1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29284_ (.CLK(clock),
    .D(_02297_),
    .Q(\decode.regfile.registers_1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29285_ (.CLK(clock),
    .D(_02298_),
    .Q(\decode.regfile.registers_1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29286_ (.CLK(clock),
    .D(_02299_),
    .Q(\decode.regfile.registers_1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29287_ (.CLK(clock),
    .D(_02300_),
    .Q(\decode.regfile.registers_1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29288_ (.CLK(clock),
    .D(_02301_),
    .Q(\decode.regfile.registers_1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29289_ (.CLK(clock),
    .D(_02302_),
    .Q(\decode.regfile.registers_1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29290_ (.CLK(clock),
    .D(_02303_),
    .Q(\decode.regfile.registers_1[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29291_ (.CLK(clock),
    .D(_02304_),
    .Q(\decode.regfile.registers_1[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29292_ (.CLK(clock),
    .D(_02305_),
    .Q(\decode.regfile.registers_1[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29293_ (.CLK(clock),
    .D(_02306_),
    .Q(\decode.regfile.registers_1[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29294_ (.CLK(clock),
    .D(_02307_),
    .Q(\decode.regfile.registers_1[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29295_ (.CLK(clock),
    .D(_02308_),
    .Q(\decode.regfile.registers_1[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29296_ (.CLK(clock),
    .D(_02309_),
    .Q(\decode.regfile.registers_1[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29297_ (.CLK(clock),
    .D(_02310_),
    .Q(\decode.regfile.registers_1[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29298_ (.CLK(clock),
    .D(_02311_),
    .Q(\decode.regfile.registers_1[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29299_ (.CLK(clock),
    .D(_02312_),
    .Q(\decode.regfile.registers_1[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29300_ (.CLK(clock),
    .D(_02313_),
    .Q(\decode.regfile.registers_1[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29301_ (.CLK(clock),
    .D(_02314_),
    .Q(\decode.regfile.registers_1[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29302_ (.CLK(clock),
    .D(_02315_),
    .Q(\decode.regfile.registers_1[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29303_ (.CLK(clock),
    .D(_02316_),
    .Q(\decode.regfile.registers_1[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29304_ (.CLK(clock),
    .D(_02317_),
    .Q(\decode.regfile.registers_1[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29305_ (.CLK(clock),
    .D(_02318_),
    .Q(\decode.regfile.registers_1[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29306_ (.CLK(clock),
    .D(_02319_),
    .Q(\decode.regfile.registers_2[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29307_ (.CLK(clock),
    .D(_02320_),
    .Q(\decode.regfile.registers_2[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29308_ (.CLK(clock),
    .D(_02321_),
    .Q(\decode.regfile.registers_2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29309_ (.CLK(clock),
    .D(_02322_),
    .Q(\decode.regfile.registers_2[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29310_ (.CLK(clock),
    .D(_02323_),
    .Q(\decode.regfile.registers_2[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29311_ (.CLK(clock),
    .D(_02324_),
    .Q(\decode.regfile.registers_2[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29312_ (.CLK(clock),
    .D(_02325_),
    .Q(\decode.regfile.registers_2[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29313_ (.CLK(clock),
    .D(_02326_),
    .Q(\decode.regfile.registers_2[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29314_ (.CLK(clock),
    .D(_02327_),
    .Q(\decode.regfile.registers_2[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29315_ (.CLK(clock),
    .D(_02328_),
    .Q(\decode.regfile.registers_2[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29316_ (.CLK(clock),
    .D(_02329_),
    .Q(\decode.regfile.registers_2[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29317_ (.CLK(clock),
    .D(_02330_),
    .Q(\decode.regfile.registers_2[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29318_ (.CLK(clock),
    .D(_02331_),
    .Q(\decode.regfile.registers_2[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29319_ (.CLK(clock),
    .D(_02332_),
    .Q(\decode.regfile.registers_2[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29320_ (.CLK(clock),
    .D(_02333_),
    .Q(\decode.regfile.registers_2[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29321_ (.CLK(clock),
    .D(_02334_),
    .Q(\decode.regfile.registers_2[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29322_ (.CLK(clock),
    .D(_02335_),
    .Q(\decode.regfile.registers_2[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29323_ (.CLK(clock),
    .D(_02336_),
    .Q(\decode.regfile.registers_2[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29324_ (.CLK(clock),
    .D(_02337_),
    .Q(\decode.regfile.registers_2[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29325_ (.CLK(clock),
    .D(_02338_),
    .Q(\decode.regfile.registers_2[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29326_ (.CLK(clock),
    .D(_02339_),
    .Q(\decode.regfile.registers_2[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29327_ (.CLK(clock),
    .D(_02340_),
    .Q(\decode.regfile.registers_2[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29328_ (.CLK(clock),
    .D(_02341_),
    .Q(\decode.regfile.registers_2[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29329_ (.CLK(clock),
    .D(_02342_),
    .Q(\decode.regfile.registers_2[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29330_ (.CLK(clock),
    .D(_02343_),
    .Q(\decode.regfile.registers_2[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29331_ (.CLK(clock),
    .D(_02344_),
    .Q(\decode.regfile.registers_2[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29332_ (.CLK(clock),
    .D(_02345_),
    .Q(\decode.regfile.registers_2[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29333_ (.CLK(clock),
    .D(_02346_),
    .Q(\decode.regfile.registers_2[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29334_ (.CLK(clock),
    .D(_02347_),
    .Q(\decode.regfile.registers_2[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29335_ (.CLK(clock),
    .D(_02348_),
    .Q(\decode.regfile.registers_2[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29336_ (.CLK(clock),
    .D(_02349_),
    .Q(\decode.regfile.registers_2[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29337_ (.CLK(clock),
    .D(_02350_),
    .Q(\decode.regfile.registers_2[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29338_ (.CLK(clock),
    .D(_02351_),
    .Q(\decode.regfile.registers_3[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29339_ (.CLK(clock),
    .D(_02352_),
    .Q(\decode.regfile.registers_3[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29340_ (.CLK(clock),
    .D(_02353_),
    .Q(\decode.regfile.registers_3[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29341_ (.CLK(clock),
    .D(_02354_),
    .Q(\decode.regfile.registers_3[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29342_ (.CLK(clock),
    .D(_02355_),
    .Q(\decode.regfile.registers_3[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29343_ (.CLK(clock),
    .D(_02356_),
    .Q(\decode.regfile.registers_3[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29344_ (.CLK(clock),
    .D(_02357_),
    .Q(\decode.regfile.registers_3[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29345_ (.CLK(clock),
    .D(_02358_),
    .Q(\decode.regfile.registers_3[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29346_ (.CLK(clock),
    .D(_02359_),
    .Q(\decode.regfile.registers_3[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29347_ (.CLK(clock),
    .D(_02360_),
    .Q(\decode.regfile.registers_3[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29348_ (.CLK(clock),
    .D(_02361_),
    .Q(\decode.regfile.registers_3[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29349_ (.CLK(clock),
    .D(_02362_),
    .Q(\decode.regfile.registers_3[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29350_ (.CLK(clock),
    .D(_02363_),
    .Q(\decode.regfile.registers_3[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29351_ (.CLK(clock),
    .D(_02364_),
    .Q(\decode.regfile.registers_3[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29352_ (.CLK(clock),
    .D(_02365_),
    .Q(\decode.regfile.registers_3[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29353_ (.CLK(clock),
    .D(_02366_),
    .Q(\decode.regfile.registers_3[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29354_ (.CLK(clock),
    .D(_02367_),
    .Q(\decode.regfile.registers_3[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29355_ (.CLK(clock),
    .D(_02368_),
    .Q(\decode.regfile.registers_3[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29356_ (.CLK(clock),
    .D(_02369_),
    .Q(\decode.regfile.registers_3[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29357_ (.CLK(clock),
    .D(_02370_),
    .Q(\decode.regfile.registers_3[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29358_ (.CLK(clock),
    .D(_02371_),
    .Q(\decode.regfile.registers_3[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29359_ (.CLK(clock),
    .D(_02372_),
    .Q(\decode.regfile.registers_3[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29360_ (.CLK(clock),
    .D(_02373_),
    .Q(\decode.regfile.registers_3[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29361_ (.CLK(clock),
    .D(_02374_),
    .Q(\decode.regfile.registers_3[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29362_ (.CLK(clock),
    .D(_02375_),
    .Q(\decode.regfile.registers_3[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29363_ (.CLK(clock),
    .D(_02376_),
    .Q(\decode.regfile.registers_3[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29364_ (.CLK(clock),
    .D(_02377_),
    .Q(\decode.regfile.registers_3[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29365_ (.CLK(clock),
    .D(_02378_),
    .Q(\decode.regfile.registers_3[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29366_ (.CLK(clock),
    .D(_02379_),
    .Q(\decode.regfile.registers_3[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29367_ (.CLK(clock),
    .D(_02380_),
    .Q(\decode.regfile.registers_3[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29368_ (.CLK(clock),
    .D(_02381_),
    .Q(\decode.regfile.registers_3[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29369_ (.CLK(clock),
    .D(_02382_),
    .Q(\decode.regfile.registers_3[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29370_ (.CLK(clock),
    .D(_02383_),
    .Q(\decode.regfile.registers_4[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29371_ (.CLK(clock),
    .D(_02384_),
    .Q(\decode.regfile.registers_4[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29372_ (.CLK(clock),
    .D(_02385_),
    .Q(\decode.regfile.registers_4[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29373_ (.CLK(clock),
    .D(_02386_),
    .Q(\decode.regfile.registers_4[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29374_ (.CLK(clock),
    .D(_02387_),
    .Q(\decode.regfile.registers_4[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29375_ (.CLK(clock),
    .D(_02388_),
    .Q(\decode.regfile.registers_4[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29376_ (.CLK(clock),
    .D(_02389_),
    .Q(\decode.regfile.registers_4[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29377_ (.CLK(clock),
    .D(_02390_),
    .Q(\decode.regfile.registers_4[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29378_ (.CLK(clock),
    .D(_02391_),
    .Q(\decode.regfile.registers_4[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29379_ (.CLK(clock),
    .D(_02392_),
    .Q(\decode.regfile.registers_4[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29380_ (.CLK(clock),
    .D(_02393_),
    .Q(\decode.regfile.registers_4[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29381_ (.CLK(clock),
    .D(_02394_),
    .Q(\decode.regfile.registers_4[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29382_ (.CLK(clock),
    .D(_02395_),
    .Q(\decode.regfile.registers_4[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29383_ (.CLK(clock),
    .D(_02396_),
    .Q(\decode.regfile.registers_4[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29384_ (.CLK(clock),
    .D(_02397_),
    .Q(\decode.regfile.registers_4[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29385_ (.CLK(clock),
    .D(_02398_),
    .Q(\decode.regfile.registers_4[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29386_ (.CLK(clock),
    .D(_02399_),
    .Q(\decode.regfile.registers_4[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29387_ (.CLK(clock),
    .D(_02400_),
    .Q(\decode.regfile.registers_4[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29388_ (.CLK(clock),
    .D(_02401_),
    .Q(\decode.regfile.registers_4[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29389_ (.CLK(clock),
    .D(_02402_),
    .Q(\decode.regfile.registers_4[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29390_ (.CLK(clock),
    .D(_02403_),
    .Q(\decode.regfile.registers_4[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29391_ (.CLK(clock),
    .D(_02404_),
    .Q(\decode.regfile.registers_4[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29392_ (.CLK(clock),
    .D(_02405_),
    .Q(\decode.regfile.registers_4[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29393_ (.CLK(clock),
    .D(_02406_),
    .Q(\decode.regfile.registers_4[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29394_ (.CLK(clock),
    .D(_02407_),
    .Q(\decode.regfile.registers_4[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29395_ (.CLK(clock),
    .D(_02408_),
    .Q(\decode.regfile.registers_4[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29396_ (.CLK(clock),
    .D(_02409_),
    .Q(\decode.regfile.registers_4[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29397_ (.CLK(clock),
    .D(_02410_),
    .Q(\decode.regfile.registers_4[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29398_ (.CLK(clock),
    .D(_02411_),
    .Q(\decode.regfile.registers_4[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29399_ (.CLK(clock),
    .D(_02412_),
    .Q(\decode.regfile.registers_4[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29400_ (.CLK(clock),
    .D(_02413_),
    .Q(\decode.regfile.registers_4[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29401_ (.CLK(clock),
    .D(_02414_),
    .Q(\decode.regfile.registers_4[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29402_ (.CLK(clock),
    .D(_02415_),
    .Q(\decode.regfile.registers_5[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29403_ (.CLK(clock),
    .D(_02416_),
    .Q(\decode.regfile.registers_5[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29404_ (.CLK(clock),
    .D(_02417_),
    .Q(\decode.regfile.registers_5[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29405_ (.CLK(clock),
    .D(_02418_),
    .Q(\decode.regfile.registers_5[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29406_ (.CLK(clock),
    .D(_02419_),
    .Q(\decode.regfile.registers_5[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29407_ (.CLK(clock),
    .D(_02420_),
    .Q(\decode.regfile.registers_5[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29408_ (.CLK(clock),
    .D(_02421_),
    .Q(\decode.regfile.registers_5[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29409_ (.CLK(clock),
    .D(_02422_),
    .Q(\decode.regfile.registers_5[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29410_ (.CLK(clock),
    .D(_02423_),
    .Q(\decode.regfile.registers_5[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29411_ (.CLK(clock),
    .D(_02424_),
    .Q(\decode.regfile.registers_5[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29412_ (.CLK(clock),
    .D(_02425_),
    .Q(\decode.regfile.registers_5[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29413_ (.CLK(clock),
    .D(_02426_),
    .Q(\decode.regfile.registers_5[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29414_ (.CLK(clock),
    .D(_02427_),
    .Q(\decode.regfile.registers_5[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29415_ (.CLK(clock),
    .D(_02428_),
    .Q(\decode.regfile.registers_5[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29416_ (.CLK(clock),
    .D(_02429_),
    .Q(\decode.regfile.registers_5[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29417_ (.CLK(clock),
    .D(_02430_),
    .Q(\decode.regfile.registers_5[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29418_ (.CLK(clock),
    .D(_02431_),
    .Q(\decode.regfile.registers_5[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29419_ (.CLK(clock),
    .D(_02432_),
    .Q(\decode.regfile.registers_5[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29420_ (.CLK(clock),
    .D(_02433_),
    .Q(\decode.regfile.registers_5[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29421_ (.CLK(clock),
    .D(_02434_),
    .Q(\decode.regfile.registers_5[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29422_ (.CLK(clock),
    .D(_02435_),
    .Q(\decode.regfile.registers_5[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29423_ (.CLK(clock),
    .D(_02436_),
    .Q(\decode.regfile.registers_5[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29424_ (.CLK(clock),
    .D(_02437_),
    .Q(\decode.regfile.registers_5[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29425_ (.CLK(clock),
    .D(_02438_),
    .Q(\decode.regfile.registers_5[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29426_ (.CLK(clock),
    .D(_02439_),
    .Q(\decode.regfile.registers_5[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29427_ (.CLK(clock),
    .D(_02440_),
    .Q(\decode.regfile.registers_5[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29428_ (.CLK(clock),
    .D(_02441_),
    .Q(\decode.regfile.registers_5[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29429_ (.CLK(clock),
    .D(_02442_),
    .Q(\decode.regfile.registers_5[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29430_ (.CLK(clock),
    .D(_02443_),
    .Q(\decode.regfile.registers_5[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29431_ (.CLK(clock),
    .D(_02444_),
    .Q(\decode.regfile.registers_5[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29432_ (.CLK(clock),
    .D(_02445_),
    .Q(\decode.regfile.registers_5[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29433_ (.CLK(clock),
    .D(_02446_),
    .Q(\decode.regfile.registers_5[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29434_ (.CLK(clock),
    .D(_02447_),
    .Q(\decode.regfile.registers_6[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29435_ (.CLK(clock),
    .D(_02448_),
    .Q(\decode.regfile.registers_6[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29436_ (.CLK(clock),
    .D(_02449_),
    .Q(\decode.regfile.registers_6[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29437_ (.CLK(clock),
    .D(_02450_),
    .Q(\decode.regfile.registers_6[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29438_ (.CLK(clock),
    .D(_02451_),
    .Q(\decode.regfile.registers_6[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29439_ (.CLK(clock),
    .D(_02452_),
    .Q(\decode.regfile.registers_6[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29440_ (.CLK(clock),
    .D(_02453_),
    .Q(\decode.regfile.registers_6[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29441_ (.CLK(clock),
    .D(_02454_),
    .Q(\decode.regfile.registers_6[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29442_ (.CLK(clock),
    .D(_02455_),
    .Q(\decode.regfile.registers_6[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29443_ (.CLK(clock),
    .D(_02456_),
    .Q(\decode.regfile.registers_6[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29444_ (.CLK(clock),
    .D(_02457_),
    .Q(\decode.regfile.registers_6[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29445_ (.CLK(clock),
    .D(_02458_),
    .Q(\decode.regfile.registers_6[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29446_ (.CLK(clock),
    .D(_02459_),
    .Q(\decode.regfile.registers_6[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29447_ (.CLK(clock),
    .D(_02460_),
    .Q(\decode.regfile.registers_6[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29448_ (.CLK(clock),
    .D(_02461_),
    .Q(\decode.regfile.registers_6[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29449_ (.CLK(clock),
    .D(_02462_),
    .Q(\decode.regfile.registers_6[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29450_ (.CLK(clock),
    .D(_02463_),
    .Q(\decode.regfile.registers_6[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29451_ (.CLK(clock),
    .D(_02464_),
    .Q(\decode.regfile.registers_6[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29452_ (.CLK(clock),
    .D(_02465_),
    .Q(\decode.regfile.registers_6[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29453_ (.CLK(clock),
    .D(_02466_),
    .Q(\decode.regfile.registers_6[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29454_ (.CLK(clock),
    .D(_02467_),
    .Q(\decode.regfile.registers_6[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29455_ (.CLK(clock),
    .D(_02468_),
    .Q(\decode.regfile.registers_6[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29456_ (.CLK(clock),
    .D(_02469_),
    .Q(\decode.regfile.registers_6[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29457_ (.CLK(clock),
    .D(_02470_),
    .Q(\decode.regfile.registers_6[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29458_ (.CLK(clock),
    .D(_02471_),
    .Q(\decode.regfile.registers_6[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29459_ (.CLK(clock),
    .D(_02472_),
    .Q(\decode.regfile.registers_6[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29460_ (.CLK(clock),
    .D(_02473_),
    .Q(\decode.regfile.registers_6[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29461_ (.CLK(clock),
    .D(_02474_),
    .Q(\decode.regfile.registers_6[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29462_ (.CLK(clock),
    .D(_02475_),
    .Q(\decode.regfile.registers_6[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29463_ (.CLK(clock),
    .D(_02476_),
    .Q(\decode.regfile.registers_6[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29464_ (.CLK(clock),
    .D(_02477_),
    .Q(\decode.regfile.registers_6[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29465_ (.CLK(clock),
    .D(_02478_),
    .Q(\decode.regfile.registers_6[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29466_ (.CLK(clock),
    .D(_02479_),
    .Q(\decode.regfile.registers_7[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29467_ (.CLK(clock),
    .D(_02480_),
    .Q(\decode.regfile.registers_7[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29468_ (.CLK(clock),
    .D(_02481_),
    .Q(\decode.regfile.registers_7[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29469_ (.CLK(clock),
    .D(_02482_),
    .Q(\decode.regfile.registers_7[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29470_ (.CLK(clock),
    .D(_02483_),
    .Q(\decode.regfile.registers_7[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29471_ (.CLK(clock),
    .D(_02484_),
    .Q(\decode.regfile.registers_7[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29472_ (.CLK(clock),
    .D(_02485_),
    .Q(\decode.regfile.registers_7[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29473_ (.CLK(clock),
    .D(_02486_),
    .Q(\decode.regfile.registers_7[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29474_ (.CLK(clock),
    .D(_02487_),
    .Q(\decode.regfile.registers_7[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29475_ (.CLK(clock),
    .D(_02488_),
    .Q(\decode.regfile.registers_7[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29476_ (.CLK(clock),
    .D(_02489_),
    .Q(\decode.regfile.registers_7[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29477_ (.CLK(clock),
    .D(_02490_),
    .Q(\decode.regfile.registers_7[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29478_ (.CLK(clock),
    .D(_02491_),
    .Q(\decode.regfile.registers_7[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29479_ (.CLK(clock),
    .D(_02492_),
    .Q(\decode.regfile.registers_7[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29480_ (.CLK(clock),
    .D(_02493_),
    .Q(\decode.regfile.registers_7[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29481_ (.CLK(clock),
    .D(_02494_),
    .Q(\decode.regfile.registers_7[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29482_ (.CLK(clock),
    .D(_02495_),
    .Q(\decode.regfile.registers_7[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29483_ (.CLK(clock),
    .D(_02496_),
    .Q(\decode.regfile.registers_7[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29484_ (.CLK(clock),
    .D(_02497_),
    .Q(\decode.regfile.registers_7[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29485_ (.CLK(clock),
    .D(_02498_),
    .Q(\decode.regfile.registers_7[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29486_ (.CLK(clock),
    .D(_02499_),
    .Q(\decode.regfile.registers_7[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29487_ (.CLK(clock),
    .D(_02500_),
    .Q(\decode.regfile.registers_7[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29488_ (.CLK(clock),
    .D(_02501_),
    .Q(\decode.regfile.registers_7[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29489_ (.CLK(clock),
    .D(_02502_),
    .Q(\decode.regfile.registers_7[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29490_ (.CLK(clock),
    .D(_02503_),
    .Q(\decode.regfile.registers_7[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29491_ (.CLK(clock),
    .D(_02504_),
    .Q(\decode.regfile.registers_7[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29492_ (.CLK(clock),
    .D(_02505_),
    .Q(\decode.regfile.registers_7[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29493_ (.CLK(clock),
    .D(_02506_),
    .Q(\decode.regfile.registers_7[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29494_ (.CLK(clock),
    .D(_02507_),
    .Q(\decode.regfile.registers_7[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29495_ (.CLK(clock),
    .D(_02508_),
    .Q(\decode.regfile.registers_7[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29496_ (.CLK(clock),
    .D(_02509_),
    .Q(\decode.regfile.registers_7[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29497_ (.CLK(clock),
    .D(_02510_),
    .Q(\decode.regfile.registers_7[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29498_ (.CLK(clock),
    .D(_02511_),
    .Q(\decode.regfile.registers_8[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29499_ (.CLK(clock),
    .D(_02512_),
    .Q(\decode.regfile.registers_8[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29500_ (.CLK(clock),
    .D(_02513_),
    .Q(\decode.regfile.registers_8[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29501_ (.CLK(clock),
    .D(_02514_),
    .Q(\decode.regfile.registers_8[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29502_ (.CLK(clock),
    .D(_02515_),
    .Q(\decode.regfile.registers_8[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29503_ (.CLK(clock),
    .D(_02516_),
    .Q(\decode.regfile.registers_8[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29504_ (.CLK(clock),
    .D(_02517_),
    .Q(\decode.regfile.registers_8[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29505_ (.CLK(clock),
    .D(_02518_),
    .Q(\decode.regfile.registers_8[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29506_ (.CLK(clock),
    .D(_02519_),
    .Q(\decode.regfile.registers_8[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29507_ (.CLK(clock),
    .D(_02520_),
    .Q(\decode.regfile.registers_8[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29508_ (.CLK(clock),
    .D(_02521_),
    .Q(\decode.regfile.registers_8[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29509_ (.CLK(clock),
    .D(_02522_),
    .Q(\decode.regfile.registers_8[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29510_ (.CLK(clock),
    .D(_02523_),
    .Q(\decode.regfile.registers_8[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29511_ (.CLK(clock),
    .D(_02524_),
    .Q(\decode.regfile.registers_8[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29512_ (.CLK(clock),
    .D(_02525_),
    .Q(\decode.regfile.registers_8[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29513_ (.CLK(clock),
    .D(_02526_),
    .Q(\decode.regfile.registers_8[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29514_ (.CLK(clock),
    .D(_02527_),
    .Q(\decode.regfile.registers_8[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29515_ (.CLK(clock),
    .D(_02528_),
    .Q(\decode.regfile.registers_8[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29516_ (.CLK(clock),
    .D(_02529_),
    .Q(\decode.regfile.registers_8[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29517_ (.CLK(clock),
    .D(_02530_),
    .Q(\decode.regfile.registers_8[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29518_ (.CLK(clock),
    .D(_02531_),
    .Q(\decode.regfile.registers_8[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29519_ (.CLK(clock),
    .D(_02532_),
    .Q(\decode.regfile.registers_8[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29520_ (.CLK(clock),
    .D(_02533_),
    .Q(\decode.regfile.registers_8[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29521_ (.CLK(clock),
    .D(_02534_),
    .Q(\decode.regfile.registers_8[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29522_ (.CLK(clock),
    .D(_02535_),
    .Q(\decode.regfile.registers_8[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29523_ (.CLK(clock),
    .D(_02536_),
    .Q(\decode.regfile.registers_8[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29524_ (.CLK(clock),
    .D(_02537_),
    .Q(\decode.regfile.registers_8[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29525_ (.CLK(clock),
    .D(_02538_),
    .Q(\decode.regfile.registers_8[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29526_ (.CLK(clock),
    .D(_02539_),
    .Q(\decode.regfile.registers_8[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29527_ (.CLK(clock),
    .D(_02540_),
    .Q(\decode.regfile.registers_8[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29528_ (.CLK(clock),
    .D(_02541_),
    .Q(\decode.regfile.registers_8[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29529_ (.CLK(clock),
    .D(_02542_),
    .Q(\decode.regfile.registers_8[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29530_ (.CLK(clock),
    .D(_02543_),
    .Q(\decode.regfile.registers_9[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29531_ (.CLK(clock),
    .D(_02544_),
    .Q(\decode.regfile.registers_9[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29532_ (.CLK(clock),
    .D(_02545_),
    .Q(\decode.regfile.registers_9[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29533_ (.CLK(clock),
    .D(_02546_),
    .Q(\decode.regfile.registers_9[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29534_ (.CLK(clock),
    .D(_02547_),
    .Q(\decode.regfile.registers_9[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29535_ (.CLK(clock),
    .D(_02548_),
    .Q(\decode.regfile.registers_9[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29536_ (.CLK(clock),
    .D(_02549_),
    .Q(\decode.regfile.registers_9[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29537_ (.CLK(clock),
    .D(_02550_),
    .Q(\decode.regfile.registers_9[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29538_ (.CLK(clock),
    .D(_02551_),
    .Q(\decode.regfile.registers_9[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29539_ (.CLK(clock),
    .D(_02552_),
    .Q(\decode.regfile.registers_9[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29540_ (.CLK(clock),
    .D(_02553_),
    .Q(\decode.regfile.registers_9[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29541_ (.CLK(clock),
    .D(_02554_),
    .Q(\decode.regfile.registers_9[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29542_ (.CLK(clock),
    .D(_02555_),
    .Q(\decode.regfile.registers_9[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29543_ (.CLK(clock),
    .D(_02556_),
    .Q(\decode.regfile.registers_9[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29544_ (.CLK(clock),
    .D(_02557_),
    .Q(\decode.regfile.registers_9[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29545_ (.CLK(clock),
    .D(_02558_),
    .Q(\decode.regfile.registers_9[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29546_ (.CLK(clock),
    .D(_02559_),
    .Q(\decode.regfile.registers_9[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29547_ (.CLK(clock),
    .D(_02560_),
    .Q(\decode.regfile.registers_9[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29548_ (.CLK(clock),
    .D(_02561_),
    .Q(\decode.regfile.registers_9[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29549_ (.CLK(clock),
    .D(_02562_),
    .Q(\decode.regfile.registers_9[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29550_ (.CLK(clock),
    .D(_02563_),
    .Q(\decode.regfile.registers_9[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29551_ (.CLK(clock),
    .D(_02564_),
    .Q(\decode.regfile.registers_9[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29552_ (.CLK(clock),
    .D(_02565_),
    .Q(\decode.regfile.registers_9[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29553_ (.CLK(clock),
    .D(_02566_),
    .Q(\decode.regfile.registers_9[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29554_ (.CLK(clock),
    .D(_02567_),
    .Q(\decode.regfile.registers_9[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29555_ (.CLK(clock),
    .D(_02568_),
    .Q(\decode.regfile.registers_9[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29556_ (.CLK(clock),
    .D(_02569_),
    .Q(\decode.regfile.registers_9[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29557_ (.CLK(clock),
    .D(_02570_),
    .Q(\decode.regfile.registers_9[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29558_ (.CLK(clock),
    .D(_02571_),
    .Q(\decode.regfile.registers_9[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29559_ (.CLK(clock),
    .D(_02572_),
    .Q(\decode.regfile.registers_9[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29560_ (.CLK(clock),
    .D(_02573_),
    .Q(\decode.regfile.registers_9[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29561_ (.CLK(clock),
    .D(_02574_),
    .Q(\decode.regfile.registers_9[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29562_ (.CLK(clock),
    .D(_02575_),
    .Q(\decode.regfile.registers_10[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29563_ (.CLK(clock),
    .D(_02576_),
    .Q(\decode.regfile.registers_10[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29564_ (.CLK(clock),
    .D(_02577_),
    .Q(\decode.regfile.registers_10[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29565_ (.CLK(clock),
    .D(_02578_),
    .Q(\decode.regfile.registers_10[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29566_ (.CLK(clock),
    .D(_02579_),
    .Q(\decode.regfile.registers_10[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29567_ (.CLK(clock),
    .D(_02580_),
    .Q(\decode.regfile.registers_10[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29568_ (.CLK(clock),
    .D(_02581_),
    .Q(\decode.regfile.registers_10[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29569_ (.CLK(clock),
    .D(_02582_),
    .Q(\decode.regfile.registers_10[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29570_ (.CLK(clock),
    .D(_02583_),
    .Q(\decode.regfile.registers_10[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29571_ (.CLK(clock),
    .D(_02584_),
    .Q(\decode.regfile.registers_10[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29572_ (.CLK(clock),
    .D(_02585_),
    .Q(\decode.regfile.registers_10[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29573_ (.CLK(clock),
    .D(_02586_),
    .Q(\decode.regfile.registers_10[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29574_ (.CLK(clock),
    .D(_02587_),
    .Q(\decode.regfile.registers_10[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29575_ (.CLK(clock),
    .D(_02588_),
    .Q(\decode.regfile.registers_10[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29576_ (.CLK(clock),
    .D(_02589_),
    .Q(\decode.regfile.registers_10[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29577_ (.CLK(clock),
    .D(_02590_),
    .Q(\decode.regfile.registers_10[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29578_ (.CLK(clock),
    .D(_02591_),
    .Q(\decode.regfile.registers_10[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29579_ (.CLK(clock),
    .D(_02592_),
    .Q(\decode.regfile.registers_10[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29580_ (.CLK(clock),
    .D(_02593_),
    .Q(\decode.regfile.registers_10[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29581_ (.CLK(clock),
    .D(_02594_),
    .Q(\decode.regfile.registers_10[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29582_ (.CLK(clock),
    .D(_02595_),
    .Q(\decode.regfile.registers_10[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29583_ (.CLK(clock),
    .D(_02596_),
    .Q(\decode.regfile.registers_10[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29584_ (.CLK(clock),
    .D(_02597_),
    .Q(\decode.regfile.registers_10[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29585_ (.CLK(clock),
    .D(_02598_),
    .Q(\decode.regfile.registers_10[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29586_ (.CLK(clock),
    .D(_02599_),
    .Q(\decode.regfile.registers_10[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29587_ (.CLK(clock),
    .D(_02600_),
    .Q(\decode.regfile.registers_10[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29588_ (.CLK(clock),
    .D(_02601_),
    .Q(\decode.regfile.registers_10[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29589_ (.CLK(clock),
    .D(_02602_),
    .Q(\decode.regfile.registers_10[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29590_ (.CLK(clock),
    .D(_02603_),
    .Q(\decode.regfile.registers_10[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29591_ (.CLK(clock),
    .D(_02604_),
    .Q(\decode.regfile.registers_10[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29592_ (.CLK(clock),
    .D(_02605_),
    .Q(\decode.regfile.registers_10[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29593_ (.CLK(clock),
    .D(_02606_),
    .Q(\decode.regfile.registers_10[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29594_ (.CLK(clock),
    .D(_02607_),
    .Q(\decode.regfile.registers_11[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29595_ (.CLK(clock),
    .D(_02608_),
    .Q(\decode.regfile.registers_11[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29596_ (.CLK(clock),
    .D(_02609_),
    .Q(\decode.regfile.registers_11[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29597_ (.CLK(clock),
    .D(_02610_),
    .Q(\decode.regfile.registers_11[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29598_ (.CLK(clock),
    .D(_02611_),
    .Q(\decode.regfile.registers_11[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29599_ (.CLK(clock),
    .D(_02612_),
    .Q(\decode.regfile.registers_11[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29600_ (.CLK(clock),
    .D(_02613_),
    .Q(\decode.regfile.registers_11[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29601_ (.CLK(clock),
    .D(_02614_),
    .Q(\decode.regfile.registers_11[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29602_ (.CLK(clock),
    .D(_02615_),
    .Q(\decode.regfile.registers_11[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29603_ (.CLK(clock),
    .D(_02616_),
    .Q(\decode.regfile.registers_11[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29604_ (.CLK(clock),
    .D(_02617_),
    .Q(\decode.regfile.registers_11[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29605_ (.CLK(clock),
    .D(_02618_),
    .Q(\decode.regfile.registers_11[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29606_ (.CLK(clock),
    .D(_02619_),
    .Q(\decode.regfile.registers_11[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29607_ (.CLK(clock),
    .D(_02620_),
    .Q(\decode.regfile.registers_11[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29608_ (.CLK(clock),
    .D(_02621_),
    .Q(\decode.regfile.registers_11[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29609_ (.CLK(clock),
    .D(_02622_),
    .Q(\decode.regfile.registers_11[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29610_ (.CLK(clock),
    .D(_02623_),
    .Q(\decode.regfile.registers_11[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29611_ (.CLK(clock),
    .D(_02624_),
    .Q(\decode.regfile.registers_11[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29612_ (.CLK(clock),
    .D(_02625_),
    .Q(\decode.regfile.registers_11[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29613_ (.CLK(clock),
    .D(_02626_),
    .Q(\decode.regfile.registers_11[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29614_ (.CLK(clock),
    .D(_02627_),
    .Q(\decode.regfile.registers_11[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29615_ (.CLK(clock),
    .D(_02628_),
    .Q(\decode.regfile.registers_11[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29616_ (.CLK(clock),
    .D(_02629_),
    .Q(\decode.regfile.registers_11[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29617_ (.CLK(clock),
    .D(_02630_),
    .Q(\decode.regfile.registers_11[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29618_ (.CLK(clock),
    .D(_02631_),
    .Q(\decode.regfile.registers_11[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29619_ (.CLK(clock),
    .D(_02632_),
    .Q(\decode.regfile.registers_11[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29620_ (.CLK(clock),
    .D(_02633_),
    .Q(\decode.regfile.registers_11[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29621_ (.CLK(clock),
    .D(_02634_),
    .Q(\decode.regfile.registers_11[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29622_ (.CLK(clock),
    .D(_02635_),
    .Q(\decode.regfile.registers_11[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29623_ (.CLK(clock),
    .D(_02636_),
    .Q(\decode.regfile.registers_11[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29624_ (.CLK(clock),
    .D(_02637_),
    .Q(\decode.regfile.registers_11[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29625_ (.CLK(clock),
    .D(_02638_),
    .Q(\decode.regfile.registers_11[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29626_ (.CLK(clock),
    .D(_02639_),
    .Q(\decode.regfile.registers_12[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29627_ (.CLK(clock),
    .D(_02640_),
    .Q(\decode.regfile.registers_12[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29628_ (.CLK(clock),
    .D(_02641_),
    .Q(\decode.regfile.registers_12[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29629_ (.CLK(clock),
    .D(_02642_),
    .Q(\decode.regfile.registers_12[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29630_ (.CLK(clock),
    .D(_02643_),
    .Q(\decode.regfile.registers_12[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29631_ (.CLK(clock),
    .D(_02644_),
    .Q(\decode.regfile.registers_12[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29632_ (.CLK(clock),
    .D(_02645_),
    .Q(\decode.regfile.registers_12[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29633_ (.CLK(clock),
    .D(_02646_),
    .Q(\decode.regfile.registers_12[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29634_ (.CLK(clock),
    .D(_02647_),
    .Q(\decode.regfile.registers_12[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29635_ (.CLK(clock),
    .D(_02648_),
    .Q(\decode.regfile.registers_12[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29636_ (.CLK(clock),
    .D(_02649_),
    .Q(\decode.regfile.registers_12[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29637_ (.CLK(clock),
    .D(_02650_),
    .Q(\decode.regfile.registers_12[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29638_ (.CLK(clock),
    .D(_02651_),
    .Q(\decode.regfile.registers_12[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29639_ (.CLK(clock),
    .D(_02652_),
    .Q(\decode.regfile.registers_12[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29640_ (.CLK(clock),
    .D(_02653_),
    .Q(\decode.regfile.registers_12[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29641_ (.CLK(clock),
    .D(_02654_),
    .Q(\decode.regfile.registers_12[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29642_ (.CLK(clock),
    .D(_02655_),
    .Q(\decode.regfile.registers_12[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29643_ (.CLK(clock),
    .D(_02656_),
    .Q(\decode.regfile.registers_12[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29644_ (.CLK(clock),
    .D(_02657_),
    .Q(\decode.regfile.registers_12[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29645_ (.CLK(clock),
    .D(_02658_),
    .Q(\decode.regfile.registers_12[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29646_ (.CLK(clock),
    .D(_02659_),
    .Q(\decode.regfile.registers_12[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29647_ (.CLK(clock),
    .D(_02660_),
    .Q(\decode.regfile.registers_12[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29648_ (.CLK(clock),
    .D(_02661_),
    .Q(\decode.regfile.registers_12[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29649_ (.CLK(clock),
    .D(_02662_),
    .Q(\decode.regfile.registers_12[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29650_ (.CLK(clock),
    .D(_02663_),
    .Q(\decode.regfile.registers_12[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29651_ (.CLK(clock),
    .D(_02664_),
    .Q(\decode.regfile.registers_12[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29652_ (.CLK(clock),
    .D(_02665_),
    .Q(\decode.regfile.registers_12[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29653_ (.CLK(clock),
    .D(_02666_),
    .Q(\decode.regfile.registers_12[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29654_ (.CLK(clock),
    .D(_02667_),
    .Q(\decode.regfile.registers_12[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29655_ (.CLK(clock),
    .D(_02668_),
    .Q(\decode.regfile.registers_12[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29656_ (.CLK(clock),
    .D(_02669_),
    .Q(\decode.regfile.registers_12[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29657_ (.CLK(clock),
    .D(_02670_),
    .Q(\decode.regfile.registers_12[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29658_ (.CLK(clock),
    .D(_02671_),
    .Q(\decode.regfile.registers_13[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29659_ (.CLK(clock),
    .D(_02672_),
    .Q(\decode.regfile.registers_13[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29660_ (.CLK(clock),
    .D(_02673_),
    .Q(\decode.regfile.registers_13[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29661_ (.CLK(clock),
    .D(_02674_),
    .Q(\decode.regfile.registers_13[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29662_ (.CLK(clock),
    .D(_02675_),
    .Q(\decode.regfile.registers_13[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29663_ (.CLK(clock),
    .D(_02676_),
    .Q(\decode.regfile.registers_13[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29664_ (.CLK(clock),
    .D(_02677_),
    .Q(\decode.regfile.registers_13[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29665_ (.CLK(clock),
    .D(_02678_),
    .Q(\decode.regfile.registers_13[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29666_ (.CLK(clock),
    .D(_02679_),
    .Q(\decode.regfile.registers_13[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29667_ (.CLK(clock),
    .D(_02680_),
    .Q(\decode.regfile.registers_13[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29668_ (.CLK(clock),
    .D(_02681_),
    .Q(\decode.regfile.registers_13[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29669_ (.CLK(clock),
    .D(_02682_),
    .Q(\decode.regfile.registers_13[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29670_ (.CLK(clock),
    .D(_02683_),
    .Q(\decode.regfile.registers_13[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29671_ (.CLK(clock),
    .D(_02684_),
    .Q(\decode.regfile.registers_13[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29672_ (.CLK(clock),
    .D(_02685_),
    .Q(\decode.regfile.registers_13[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29673_ (.CLK(clock),
    .D(_02686_),
    .Q(\decode.regfile.registers_13[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29674_ (.CLK(clock),
    .D(_02687_),
    .Q(\decode.regfile.registers_13[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29675_ (.CLK(clock),
    .D(_02688_),
    .Q(\decode.regfile.registers_13[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29676_ (.CLK(clock),
    .D(_02689_),
    .Q(\decode.regfile.registers_13[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29677_ (.CLK(clock),
    .D(_02690_),
    .Q(\decode.regfile.registers_13[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29678_ (.CLK(clock),
    .D(_02691_),
    .Q(\decode.regfile.registers_13[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29679_ (.CLK(clock),
    .D(_02692_),
    .Q(\decode.regfile.registers_13[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29680_ (.CLK(clock),
    .D(_02693_),
    .Q(\decode.regfile.registers_13[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29681_ (.CLK(clock),
    .D(_02694_),
    .Q(\decode.regfile.registers_13[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29682_ (.CLK(clock),
    .D(_02695_),
    .Q(\decode.regfile.registers_13[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29683_ (.CLK(clock),
    .D(_02696_),
    .Q(\decode.regfile.registers_13[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29684_ (.CLK(clock),
    .D(_02697_),
    .Q(\decode.regfile.registers_13[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29685_ (.CLK(clock),
    .D(_02698_),
    .Q(\decode.regfile.registers_13[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29686_ (.CLK(clock),
    .D(_02699_),
    .Q(\decode.regfile.registers_13[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29687_ (.CLK(clock),
    .D(_02700_),
    .Q(\decode.regfile.registers_13[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29688_ (.CLK(clock),
    .D(_02701_),
    .Q(\decode.regfile.registers_13[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29689_ (.CLK(clock),
    .D(_02702_),
    .Q(\decode.regfile.registers_13[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29690_ (.CLK(clock),
    .D(_02703_),
    .Q(\decode.regfile.registers_14[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29691_ (.CLK(clock),
    .D(_02704_),
    .Q(\decode.regfile.registers_14[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29692_ (.CLK(clock),
    .D(_02705_),
    .Q(\decode.regfile.registers_14[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29693_ (.CLK(clock),
    .D(_02706_),
    .Q(\decode.regfile.registers_14[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29694_ (.CLK(clock),
    .D(_02707_),
    .Q(\decode.regfile.registers_14[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29695_ (.CLK(clock),
    .D(_02708_),
    .Q(\decode.regfile.registers_14[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29696_ (.CLK(clock),
    .D(_02709_),
    .Q(\decode.regfile.registers_14[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29697_ (.CLK(clock),
    .D(_02710_),
    .Q(\decode.regfile.registers_14[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29698_ (.CLK(clock),
    .D(_02711_),
    .Q(\decode.regfile.registers_14[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29699_ (.CLK(clock),
    .D(_02712_),
    .Q(\decode.regfile.registers_14[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29700_ (.CLK(clock),
    .D(_02713_),
    .Q(\decode.regfile.registers_14[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29701_ (.CLK(clock),
    .D(_02714_),
    .Q(\decode.regfile.registers_14[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29702_ (.CLK(clock),
    .D(_02715_),
    .Q(\decode.regfile.registers_14[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29703_ (.CLK(clock),
    .D(_02716_),
    .Q(\decode.regfile.registers_14[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29704_ (.CLK(clock),
    .D(_02717_),
    .Q(\decode.regfile.registers_14[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29705_ (.CLK(clock),
    .D(_02718_),
    .Q(\decode.regfile.registers_14[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29706_ (.CLK(clock),
    .D(_02719_),
    .Q(\decode.regfile.registers_14[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29707_ (.CLK(clock),
    .D(_02720_),
    .Q(\decode.regfile.registers_14[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29708_ (.CLK(clock),
    .D(_02721_),
    .Q(\decode.regfile.registers_14[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29709_ (.CLK(clock),
    .D(_02722_),
    .Q(\decode.regfile.registers_14[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29710_ (.CLK(clock),
    .D(_02723_),
    .Q(\decode.regfile.registers_14[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29711_ (.CLK(clock),
    .D(_02724_),
    .Q(\decode.regfile.registers_14[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29712_ (.CLK(clock),
    .D(_02725_),
    .Q(\decode.regfile.registers_14[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29713_ (.CLK(clock),
    .D(_02726_),
    .Q(\decode.regfile.registers_14[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29714_ (.CLK(clock),
    .D(_02727_),
    .Q(\decode.regfile.registers_14[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29715_ (.CLK(clock),
    .D(_02728_),
    .Q(\decode.regfile.registers_14[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29716_ (.CLK(clock),
    .D(_02729_),
    .Q(\decode.regfile.registers_14[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29717_ (.CLK(clock),
    .D(_02730_),
    .Q(\decode.regfile.registers_14[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29718_ (.CLK(clock),
    .D(_02731_),
    .Q(\decode.regfile.registers_14[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29719_ (.CLK(clock),
    .D(_02732_),
    .Q(\decode.regfile.registers_14[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29720_ (.CLK(clock),
    .D(_02733_),
    .Q(\decode.regfile.registers_14[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29721_ (.CLK(clock),
    .D(_02734_),
    .Q(\decode.regfile.registers_14[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29722_ (.CLK(clock),
    .D(_02735_),
    .Q(\decode.regfile.registers_15[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29723_ (.CLK(clock),
    .D(_02736_),
    .Q(\decode.regfile.registers_15[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29724_ (.CLK(clock),
    .D(_02737_),
    .Q(\decode.regfile.registers_15[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29725_ (.CLK(clock),
    .D(_02738_),
    .Q(\decode.regfile.registers_15[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29726_ (.CLK(clock),
    .D(_02739_),
    .Q(\decode.regfile.registers_15[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29727_ (.CLK(clock),
    .D(_02740_),
    .Q(\decode.regfile.registers_15[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29728_ (.CLK(clock),
    .D(_02741_),
    .Q(\decode.regfile.registers_15[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29729_ (.CLK(clock),
    .D(_02742_),
    .Q(\decode.regfile.registers_15[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29730_ (.CLK(clock),
    .D(_02743_),
    .Q(\decode.regfile.registers_15[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29731_ (.CLK(clock),
    .D(_02744_),
    .Q(\decode.regfile.registers_15[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29732_ (.CLK(clock),
    .D(_02745_),
    .Q(\decode.regfile.registers_15[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29733_ (.CLK(clock),
    .D(_02746_),
    .Q(\decode.regfile.registers_15[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29734_ (.CLK(clock),
    .D(_02747_),
    .Q(\decode.regfile.registers_15[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29735_ (.CLK(clock),
    .D(_02748_),
    .Q(\decode.regfile.registers_15[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29736_ (.CLK(clock),
    .D(_02749_),
    .Q(\decode.regfile.registers_15[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29737_ (.CLK(clock),
    .D(_02750_),
    .Q(\decode.regfile.registers_15[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29738_ (.CLK(clock),
    .D(_02751_),
    .Q(\decode.regfile.registers_15[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29739_ (.CLK(clock),
    .D(_02752_),
    .Q(\decode.regfile.registers_15[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29740_ (.CLK(clock),
    .D(_02753_),
    .Q(\decode.regfile.registers_15[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29741_ (.CLK(clock),
    .D(_02754_),
    .Q(\decode.regfile.registers_15[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29742_ (.CLK(clock),
    .D(_02755_),
    .Q(\decode.regfile.registers_15[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29743_ (.CLK(clock),
    .D(_02756_),
    .Q(\decode.regfile.registers_15[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29744_ (.CLK(clock),
    .D(_02757_),
    .Q(\decode.regfile.registers_15[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29745_ (.CLK(clock),
    .D(_02758_),
    .Q(\decode.regfile.registers_15[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29746_ (.CLK(clock),
    .D(_02759_),
    .Q(\decode.regfile.registers_15[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29747_ (.CLK(clock),
    .D(_02760_),
    .Q(\decode.regfile.registers_15[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29748_ (.CLK(clock),
    .D(_02761_),
    .Q(\decode.regfile.registers_15[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29749_ (.CLK(clock),
    .D(_02762_),
    .Q(\decode.regfile.registers_15[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29750_ (.CLK(clock),
    .D(_02763_),
    .Q(\decode.regfile.registers_15[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29751_ (.CLK(clock),
    .D(_02764_),
    .Q(\decode.regfile.registers_15[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29752_ (.CLK(clock),
    .D(_02765_),
    .Q(\decode.regfile.registers_15[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29753_ (.CLK(clock),
    .D(_02766_),
    .Q(\decode.regfile.registers_15[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29754_ (.CLK(clock),
    .D(_02767_),
    .Q(\decode.regfile.registers_16[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29755_ (.CLK(clock),
    .D(_02768_),
    .Q(\decode.regfile.registers_16[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29756_ (.CLK(clock),
    .D(_02769_),
    .Q(\decode.regfile.registers_16[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29757_ (.CLK(clock),
    .D(_02770_),
    .Q(\decode.regfile.registers_16[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29758_ (.CLK(clock),
    .D(_02771_),
    .Q(\decode.regfile.registers_16[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29759_ (.CLK(clock),
    .D(_02772_),
    .Q(\decode.regfile.registers_16[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29760_ (.CLK(clock),
    .D(_02773_),
    .Q(\decode.regfile.registers_16[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29761_ (.CLK(clock),
    .D(_02774_),
    .Q(\decode.regfile.registers_16[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29762_ (.CLK(clock),
    .D(_02775_),
    .Q(\decode.regfile.registers_16[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29763_ (.CLK(clock),
    .D(_02776_),
    .Q(\decode.regfile.registers_16[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29764_ (.CLK(clock),
    .D(_02777_),
    .Q(\decode.regfile.registers_16[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29765_ (.CLK(clock),
    .D(_02778_),
    .Q(\decode.regfile.registers_16[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29766_ (.CLK(clock),
    .D(_02779_),
    .Q(\decode.regfile.registers_16[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29767_ (.CLK(clock),
    .D(_02780_),
    .Q(\decode.regfile.registers_16[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29768_ (.CLK(clock),
    .D(_02781_),
    .Q(\decode.regfile.registers_16[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29769_ (.CLK(clock),
    .D(_02782_),
    .Q(\decode.regfile.registers_16[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29770_ (.CLK(clock),
    .D(_02783_),
    .Q(\decode.regfile.registers_16[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29771_ (.CLK(clock),
    .D(_02784_),
    .Q(\decode.regfile.registers_16[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29772_ (.CLK(clock),
    .D(_02785_),
    .Q(\decode.regfile.registers_16[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29773_ (.CLK(clock),
    .D(_02786_),
    .Q(\decode.regfile.registers_16[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29774_ (.CLK(clock),
    .D(_02787_),
    .Q(\decode.regfile.registers_16[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29775_ (.CLK(clock),
    .D(_02788_),
    .Q(\decode.regfile.registers_16[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29776_ (.CLK(clock),
    .D(_02789_),
    .Q(\decode.regfile.registers_16[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29777_ (.CLK(clock),
    .D(_02790_),
    .Q(\decode.regfile.registers_16[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29778_ (.CLK(clock),
    .D(_02791_),
    .Q(\decode.regfile.registers_16[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29779_ (.CLK(clock),
    .D(_02792_),
    .Q(\decode.regfile.registers_16[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29780_ (.CLK(clock),
    .D(_02793_),
    .Q(\decode.regfile.registers_16[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29781_ (.CLK(clock),
    .D(_02794_),
    .Q(\decode.regfile.registers_16[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29782_ (.CLK(clock),
    .D(_02795_),
    .Q(\decode.regfile.registers_16[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29783_ (.CLK(clock),
    .D(_02796_),
    .Q(\decode.regfile.registers_16[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29784_ (.CLK(clock),
    .D(_02797_),
    .Q(\decode.regfile.registers_16[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29785_ (.CLK(clock),
    .D(_02798_),
    .Q(\decode.regfile.registers_16[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29786_ (.CLK(clock),
    .D(_02799_),
    .Q(\decode.regfile.registers_17[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29787_ (.CLK(clock),
    .D(_02800_),
    .Q(\decode.regfile.registers_17[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29788_ (.CLK(clock),
    .D(_02801_),
    .Q(\decode.regfile.registers_17[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29789_ (.CLK(clock),
    .D(_02802_),
    .Q(\decode.regfile.registers_17[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29790_ (.CLK(clock),
    .D(_02803_),
    .Q(\decode.regfile.registers_17[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29791_ (.CLK(clock),
    .D(_02804_),
    .Q(\decode.regfile.registers_17[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29792_ (.CLK(clock),
    .D(_02805_),
    .Q(\decode.regfile.registers_17[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29793_ (.CLK(clock),
    .D(_02806_),
    .Q(\decode.regfile.registers_17[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29794_ (.CLK(clock),
    .D(_02807_),
    .Q(\decode.regfile.registers_17[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29795_ (.CLK(clock),
    .D(_02808_),
    .Q(\decode.regfile.registers_17[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29796_ (.CLK(clock),
    .D(_02809_),
    .Q(\decode.regfile.registers_17[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29797_ (.CLK(clock),
    .D(_02810_),
    .Q(\decode.regfile.registers_17[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29798_ (.CLK(clock),
    .D(_02811_),
    .Q(\decode.regfile.registers_17[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29799_ (.CLK(clock),
    .D(_02812_),
    .Q(\decode.regfile.registers_17[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29800_ (.CLK(clock),
    .D(_02813_),
    .Q(\decode.regfile.registers_17[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29801_ (.CLK(clock),
    .D(_02814_),
    .Q(\decode.regfile.registers_17[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29802_ (.CLK(clock),
    .D(_02815_),
    .Q(\decode.regfile.registers_17[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29803_ (.CLK(clock),
    .D(_02816_),
    .Q(\decode.regfile.registers_17[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29804_ (.CLK(clock),
    .D(_02817_),
    .Q(\decode.regfile.registers_17[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29805_ (.CLK(clock),
    .D(_02818_),
    .Q(\decode.regfile.registers_17[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29806_ (.CLK(clock),
    .D(_02819_),
    .Q(\decode.regfile.registers_17[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29807_ (.CLK(clock),
    .D(_02820_),
    .Q(\decode.regfile.registers_17[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29808_ (.CLK(clock),
    .D(_02821_),
    .Q(\decode.regfile.registers_17[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29809_ (.CLK(clock),
    .D(_02822_),
    .Q(\decode.regfile.registers_17[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29810_ (.CLK(clock),
    .D(_02823_),
    .Q(\decode.regfile.registers_17[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29811_ (.CLK(clock),
    .D(_02824_),
    .Q(\decode.regfile.registers_17[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29812_ (.CLK(clock),
    .D(_02825_),
    .Q(\decode.regfile.registers_17[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29813_ (.CLK(clock),
    .D(_02826_),
    .Q(\decode.regfile.registers_17[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29814_ (.CLK(clock),
    .D(_02827_),
    .Q(\decode.regfile.registers_17[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29815_ (.CLK(clock),
    .D(_02828_),
    .Q(\decode.regfile.registers_17[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29816_ (.CLK(clock),
    .D(_02829_),
    .Q(\decode.regfile.registers_17[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29817_ (.CLK(clock),
    .D(_02830_),
    .Q(\decode.regfile.registers_17[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29818_ (.CLK(clock),
    .D(_02831_),
    .Q(\decode.regfile.registers_18[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29819_ (.CLK(clock),
    .D(_02832_),
    .Q(\decode.regfile.registers_18[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29820_ (.CLK(clock),
    .D(_02833_),
    .Q(\decode.regfile.registers_18[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29821_ (.CLK(clock),
    .D(_02834_),
    .Q(\decode.regfile.registers_18[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29822_ (.CLK(clock),
    .D(_02835_),
    .Q(\decode.regfile.registers_18[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29823_ (.CLK(clock),
    .D(_02836_),
    .Q(\decode.regfile.registers_18[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29824_ (.CLK(clock),
    .D(_02837_),
    .Q(\decode.regfile.registers_18[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29825_ (.CLK(clock),
    .D(_02838_),
    .Q(\decode.regfile.registers_18[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29826_ (.CLK(clock),
    .D(_02839_),
    .Q(\decode.regfile.registers_18[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29827_ (.CLK(clock),
    .D(_02840_),
    .Q(\decode.regfile.registers_18[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29828_ (.CLK(clock),
    .D(_02841_),
    .Q(\decode.regfile.registers_18[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29829_ (.CLK(clock),
    .D(_02842_),
    .Q(\decode.regfile.registers_18[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29830_ (.CLK(clock),
    .D(_02843_),
    .Q(\decode.regfile.registers_18[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29831_ (.CLK(clock),
    .D(_02844_),
    .Q(\decode.regfile.registers_18[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29832_ (.CLK(clock),
    .D(_02845_),
    .Q(\decode.regfile.registers_18[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29833_ (.CLK(clock),
    .D(_02846_),
    .Q(\decode.regfile.registers_18[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29834_ (.CLK(clock),
    .D(_02847_),
    .Q(\decode.regfile.registers_18[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29835_ (.CLK(clock),
    .D(_02848_),
    .Q(\decode.regfile.registers_18[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29836_ (.CLK(clock),
    .D(_02849_),
    .Q(\decode.regfile.registers_18[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29837_ (.CLK(clock),
    .D(_02850_),
    .Q(\decode.regfile.registers_18[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29838_ (.CLK(clock),
    .D(_02851_),
    .Q(\decode.regfile.registers_18[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29839_ (.CLK(clock),
    .D(_02852_),
    .Q(\decode.regfile.registers_18[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29840_ (.CLK(clock),
    .D(_02853_),
    .Q(\decode.regfile.registers_18[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29841_ (.CLK(clock),
    .D(_02854_),
    .Q(\decode.regfile.registers_18[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29842_ (.CLK(clock),
    .D(_02855_),
    .Q(\decode.regfile.registers_18[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29843_ (.CLK(clock),
    .D(_02856_),
    .Q(\decode.regfile.registers_18[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29844_ (.CLK(clock),
    .D(_02857_),
    .Q(\decode.regfile.registers_18[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29845_ (.CLK(clock),
    .D(_02858_),
    .Q(\decode.regfile.registers_18[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29846_ (.CLK(clock),
    .D(_02859_),
    .Q(\decode.regfile.registers_18[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29847_ (.CLK(clock),
    .D(_02860_),
    .Q(\decode.regfile.registers_18[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29848_ (.CLK(clock),
    .D(_02861_),
    .Q(\decode.regfile.registers_18[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29849_ (.CLK(clock),
    .D(_02862_),
    .Q(\decode.regfile.registers_18[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29850_ (.CLK(clock),
    .D(_02863_),
    .Q(\decode.regfile.registers_19[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29851_ (.CLK(clock),
    .D(_02864_),
    .Q(\decode.regfile.registers_19[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29852_ (.CLK(clock),
    .D(_02865_),
    .Q(\decode.regfile.registers_19[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29853_ (.CLK(clock),
    .D(_02866_),
    .Q(\decode.regfile.registers_19[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29854_ (.CLK(clock),
    .D(_02867_),
    .Q(\decode.regfile.registers_19[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29855_ (.CLK(clock),
    .D(_02868_),
    .Q(\decode.regfile.registers_19[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29856_ (.CLK(clock),
    .D(_02869_),
    .Q(\decode.regfile.registers_19[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29857_ (.CLK(clock),
    .D(_02870_),
    .Q(\decode.regfile.registers_19[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29858_ (.CLK(clock),
    .D(_02871_),
    .Q(\decode.regfile.registers_19[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29859_ (.CLK(clock),
    .D(_02872_),
    .Q(\decode.regfile.registers_19[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29860_ (.CLK(clock),
    .D(_02873_),
    .Q(\decode.regfile.registers_19[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29861_ (.CLK(clock),
    .D(_02874_),
    .Q(\decode.regfile.registers_19[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29862_ (.CLK(clock),
    .D(_02875_),
    .Q(\decode.regfile.registers_19[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29863_ (.CLK(clock),
    .D(_02876_),
    .Q(\decode.regfile.registers_19[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29864_ (.CLK(clock),
    .D(_02877_),
    .Q(\decode.regfile.registers_19[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29865_ (.CLK(clock),
    .D(_02878_),
    .Q(\decode.regfile.registers_19[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29866_ (.CLK(clock),
    .D(_02879_),
    .Q(\decode.regfile.registers_19[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29867_ (.CLK(clock),
    .D(_02880_),
    .Q(\decode.regfile.registers_19[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29868_ (.CLK(clock),
    .D(_02881_),
    .Q(\decode.regfile.registers_19[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29869_ (.CLK(clock),
    .D(_02882_),
    .Q(\decode.regfile.registers_19[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29870_ (.CLK(clock),
    .D(_02883_),
    .Q(\decode.regfile.registers_19[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29871_ (.CLK(clock),
    .D(_02884_),
    .Q(\decode.regfile.registers_19[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29872_ (.CLK(clock),
    .D(_02885_),
    .Q(\decode.regfile.registers_19[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29873_ (.CLK(clock),
    .D(_02886_),
    .Q(\decode.regfile.registers_19[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29874_ (.CLK(clock),
    .D(_02887_),
    .Q(\decode.regfile.registers_19[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29875_ (.CLK(clock),
    .D(_02888_),
    .Q(\decode.regfile.registers_19[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29876_ (.CLK(clock),
    .D(_02889_),
    .Q(\decode.regfile.registers_19[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29877_ (.CLK(clock),
    .D(_02890_),
    .Q(\decode.regfile.registers_19[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29878_ (.CLK(clock),
    .D(_02891_),
    .Q(\decode.regfile.registers_19[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29879_ (.CLK(clock),
    .D(_02892_),
    .Q(\decode.regfile.registers_19[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29880_ (.CLK(clock),
    .D(_02893_),
    .Q(\decode.regfile.registers_19[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29881_ (.CLK(clock),
    .D(_02894_),
    .Q(\decode.regfile.registers_19[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29882_ (.CLK(clock),
    .D(_02895_),
    .Q(\decode.regfile.registers_20[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29883_ (.CLK(clock),
    .D(_02896_),
    .Q(\decode.regfile.registers_20[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29884_ (.CLK(clock),
    .D(_02897_),
    .Q(\decode.regfile.registers_20[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29885_ (.CLK(clock),
    .D(_02898_),
    .Q(\decode.regfile.registers_20[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29886_ (.CLK(clock),
    .D(_02899_),
    .Q(\decode.regfile.registers_20[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29887_ (.CLK(clock),
    .D(_02900_),
    .Q(\decode.regfile.registers_20[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29888_ (.CLK(clock),
    .D(_02901_),
    .Q(\decode.regfile.registers_20[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29889_ (.CLK(clock),
    .D(_02902_),
    .Q(\decode.regfile.registers_20[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29890_ (.CLK(clock),
    .D(_02903_),
    .Q(\decode.regfile.registers_20[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29891_ (.CLK(clock),
    .D(_02904_),
    .Q(\decode.regfile.registers_20[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29892_ (.CLK(clock),
    .D(_02905_),
    .Q(\decode.regfile.registers_20[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29893_ (.CLK(clock),
    .D(_02906_),
    .Q(\decode.regfile.registers_20[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29894_ (.CLK(clock),
    .D(_02907_),
    .Q(\decode.regfile.registers_20[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29895_ (.CLK(clock),
    .D(_02908_),
    .Q(\decode.regfile.registers_20[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29896_ (.CLK(clock),
    .D(_02909_),
    .Q(\decode.regfile.registers_20[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29897_ (.CLK(clock),
    .D(_02910_),
    .Q(\decode.regfile.registers_20[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29898_ (.CLK(clock),
    .D(_02911_),
    .Q(\decode.regfile.registers_20[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29899_ (.CLK(clock),
    .D(_02912_),
    .Q(\decode.regfile.registers_20[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29900_ (.CLK(clock),
    .D(_02913_),
    .Q(\decode.regfile.registers_20[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29901_ (.CLK(clock),
    .D(_02914_),
    .Q(\decode.regfile.registers_20[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29902_ (.CLK(clock),
    .D(_02915_),
    .Q(\decode.regfile.registers_20[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29903_ (.CLK(clock),
    .D(_02916_),
    .Q(\decode.regfile.registers_20[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29904_ (.CLK(clock),
    .D(_02917_),
    .Q(\decode.regfile.registers_20[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29905_ (.CLK(clock),
    .D(_02918_),
    .Q(\decode.regfile.registers_20[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29906_ (.CLK(clock),
    .D(_02919_),
    .Q(\decode.regfile.registers_20[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29907_ (.CLK(clock),
    .D(_02920_),
    .Q(\decode.regfile.registers_20[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29908_ (.CLK(clock),
    .D(_02921_),
    .Q(\decode.regfile.registers_20[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29909_ (.CLK(clock),
    .D(_02922_),
    .Q(\decode.regfile.registers_20[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29910_ (.CLK(clock),
    .D(_02923_),
    .Q(\decode.regfile.registers_20[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29911_ (.CLK(clock),
    .D(_02924_),
    .Q(\decode.regfile.registers_20[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29912_ (.CLK(clock),
    .D(_02925_),
    .Q(\decode.regfile.registers_20[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29913_ (.CLK(clock),
    .D(_02926_),
    .Q(\decode.regfile.registers_20[31] ));
 sky130_fd_sc_hd__dfxtp_2 _29914_ (.CLK(clock),
    .D(_02927_),
    .Q(\decode.regfile.registers_21[0] ));
 sky130_fd_sc_hd__dfxtp_2 _29915_ (.CLK(clock),
    .D(_02928_),
    .Q(\decode.regfile.registers_21[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29916_ (.CLK(clock),
    .D(_02929_),
    .Q(\decode.regfile.registers_21[2] ));
 sky130_fd_sc_hd__dfxtp_2 _29917_ (.CLK(clock),
    .D(_02930_),
    .Q(\decode.regfile.registers_21[3] ));
 sky130_fd_sc_hd__dfxtp_2 _29918_ (.CLK(clock),
    .D(_02931_),
    .Q(\decode.regfile.registers_21[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29919_ (.CLK(clock),
    .D(_02932_),
    .Q(\decode.regfile.registers_21[5] ));
 sky130_fd_sc_hd__dfxtp_2 _29920_ (.CLK(clock),
    .D(_02933_),
    .Q(\decode.regfile.registers_21[6] ));
 sky130_fd_sc_hd__dfxtp_2 _29921_ (.CLK(clock),
    .D(_02934_),
    .Q(\decode.regfile.registers_21[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29922_ (.CLK(clock),
    .D(_02935_),
    .Q(\decode.regfile.registers_21[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29923_ (.CLK(clock),
    .D(_02936_),
    .Q(\decode.regfile.registers_21[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29924_ (.CLK(clock),
    .D(_02937_),
    .Q(\decode.regfile.registers_21[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29925_ (.CLK(clock),
    .D(_02938_),
    .Q(\decode.regfile.registers_21[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29926_ (.CLK(clock),
    .D(_02939_),
    .Q(\decode.regfile.registers_21[12] ));
 sky130_fd_sc_hd__dfxtp_2 _29927_ (.CLK(clock),
    .D(_02940_),
    .Q(\decode.regfile.registers_21[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29928_ (.CLK(clock),
    .D(_02941_),
    .Q(\decode.regfile.registers_21[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29929_ (.CLK(clock),
    .D(_02942_),
    .Q(\decode.regfile.registers_21[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29930_ (.CLK(clock),
    .D(_02943_),
    .Q(\decode.regfile.registers_21[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29931_ (.CLK(clock),
    .D(_02944_),
    .Q(\decode.regfile.registers_21[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29932_ (.CLK(clock),
    .D(_02945_),
    .Q(\decode.regfile.registers_21[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29933_ (.CLK(clock),
    .D(_02946_),
    .Q(\decode.regfile.registers_21[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29934_ (.CLK(clock),
    .D(_02947_),
    .Q(\decode.regfile.registers_21[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29935_ (.CLK(clock),
    .D(_02948_),
    .Q(\decode.regfile.registers_21[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29936_ (.CLK(clock),
    .D(_02949_),
    .Q(\decode.regfile.registers_21[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29937_ (.CLK(clock),
    .D(_02950_),
    .Q(\decode.regfile.registers_21[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29938_ (.CLK(clock),
    .D(_02951_),
    .Q(\decode.regfile.registers_21[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29939_ (.CLK(clock),
    .D(_02952_),
    .Q(\decode.regfile.registers_21[25] ));
 sky130_fd_sc_hd__dfxtp_2 _29940_ (.CLK(clock),
    .D(_02953_),
    .Q(\decode.regfile.registers_21[26] ));
 sky130_fd_sc_hd__dfxtp_2 _29941_ (.CLK(clock),
    .D(_02954_),
    .Q(\decode.regfile.registers_21[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29942_ (.CLK(clock),
    .D(_02955_),
    .Q(\decode.regfile.registers_21[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29943_ (.CLK(clock),
    .D(_02956_),
    .Q(\decode.regfile.registers_21[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29944_ (.CLK(clock),
    .D(_02957_),
    .Q(\decode.regfile.registers_21[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29945_ (.CLK(clock),
    .D(_02958_),
    .Q(\decode.regfile.registers_21[31] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Right_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Right_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Right_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Right_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Right_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Right_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Right_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Right_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Right_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Right_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Right_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Right_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Right_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Right_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Right_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_Right_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Right_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Right_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Left_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Left_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Left_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Left_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Left_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Left_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Left_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Left_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Left_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Left_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Left_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Left_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Left_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_Left_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Left_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Left_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6027 ();
endmodule
