magic
tech sky130A
magscale 1 2
timestamp 1713182377
<< obsli1 >>
rect 1104 2159 126408 127313
<< obsm1 >>
rect 750 2048 126468 127560
<< metal2 >>
rect 43810 128921 43866 129721
rect 44454 128921 44510 129721
rect 45098 128921 45154 129721
rect 45742 128921 45798 129721
rect 68282 128921 68338 129721
rect 68926 128921 68982 129721
rect 69570 128921 69626 129721
rect 70214 128921 70270 129721
rect 70858 128921 70914 129721
rect 71502 128921 71558 129721
rect 72146 128921 72202 129721
rect 72790 128921 72846 129721
rect 73434 128921 73490 129721
rect 74078 128921 74134 129721
rect 74722 128921 74778 129721
rect 75366 128921 75422 129721
rect 76010 128921 76066 129721
rect 76654 128921 76710 129721
rect 77298 128921 77354 129721
rect 77942 128921 77998 129721
rect 78586 128921 78642 129721
rect 79230 128921 79286 129721
rect 79874 128921 79930 129721
rect 80518 128921 80574 129721
rect 81162 128921 81218 129721
rect 81806 128921 81862 129721
rect 82450 128921 82506 129721
rect 83094 128921 83150 129721
rect 83738 128921 83794 129721
rect 86958 128921 87014 129721
rect 90178 128921 90234 129721
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
<< obsm2 >>
rect 754 128865 43754 129010
rect 43922 128865 44398 129010
rect 44566 128865 45042 129010
rect 45210 128865 45686 129010
rect 45854 128865 68226 129010
rect 68394 128865 68870 129010
rect 69038 128865 69514 129010
rect 69682 128865 70158 129010
rect 70326 128865 70802 129010
rect 70970 128865 71446 129010
rect 71614 128865 72090 129010
rect 72258 128865 72734 129010
rect 72902 128865 73378 129010
rect 73546 128865 74022 129010
rect 74190 128865 74666 129010
rect 74834 128865 75310 129010
rect 75478 128865 75954 129010
rect 76122 128865 76598 129010
rect 76766 128865 77242 129010
rect 77410 128865 77886 129010
rect 78054 128865 78530 129010
rect 78698 128865 79174 129010
rect 79342 128865 79818 129010
rect 79986 128865 80462 129010
rect 80630 128865 81106 129010
rect 81274 128865 81750 129010
rect 81918 128865 82394 129010
rect 82562 128865 83038 129010
rect 83206 128865 83682 129010
rect 83850 128865 86902 129010
rect 87070 128865 90122 129010
rect 90290 128865 126112 129010
rect 754 856 126112 128865
rect 754 734 38602 856
rect 38770 734 39246 856
rect 39414 734 39890 856
rect 40058 734 40534 856
rect 40702 734 41178 856
rect 41346 734 41822 856
rect 41990 734 42466 856
rect 42634 734 43754 856
rect 43922 734 44398 856
rect 44566 734 45042 856
rect 45210 734 45686 856
rect 45854 734 46330 856
rect 46498 734 46974 856
rect 47142 734 47618 856
rect 47786 734 48262 856
rect 48430 734 48906 856
rect 49074 734 49550 856
rect 49718 734 50194 856
rect 50362 734 50838 856
rect 51006 734 51482 856
rect 51650 734 52126 856
rect 52294 734 52770 856
rect 52938 734 53414 856
rect 53582 734 54058 856
rect 54226 734 54702 856
rect 54870 734 55346 856
rect 55514 734 55990 856
rect 56158 734 56634 856
rect 56802 734 57278 856
rect 57446 734 57922 856
rect 58090 734 58566 856
rect 58734 734 59210 856
rect 59378 734 59854 856
rect 60022 734 60498 856
rect 60666 734 61142 856
rect 61310 734 61786 856
rect 61954 734 62430 856
rect 62598 734 63074 856
rect 63242 734 63718 856
rect 63886 734 64362 856
rect 64530 734 65006 856
rect 65174 734 65650 856
rect 65818 734 66294 856
rect 66462 734 66938 856
rect 67106 734 67582 856
rect 67750 734 68226 856
rect 68394 734 68870 856
rect 69038 734 69514 856
rect 69682 734 70158 856
rect 70326 734 70802 856
rect 70970 734 71446 856
rect 71614 734 72090 856
rect 72258 734 126112 856
<< metal3 >>
rect 0 126488 800 126608
rect 0 84328 800 84448
rect 0 83648 800 83768
rect 0 82968 800 83088
rect 0 82288 800 82408
rect 0 81608 800 81728
rect 0 80928 800 81048
rect 0 80248 800 80368
rect 0 79568 800 79688
rect 0 78888 800 79008
rect 0 78208 800 78328
rect 0 77528 800 77648
rect 0 76848 800 76968
rect 0 76168 800 76288
rect 0 75488 800 75608
rect 0 74808 800 74928
rect 0 74128 800 74248
rect 0 73448 800 73568
rect 0 72768 800 72888
rect 0 72088 800 72208
rect 0 71408 800 71528
rect 0 70728 800 70848
rect 0 70048 800 70168
rect 0 69368 800 69488
rect 0 68688 800 68808
rect 0 68008 800 68128
rect 0 67328 800 67448
rect 0 66648 800 66768
rect 0 65968 800 66088
rect 0 65288 800 65408
rect 0 64608 800 64728
rect 0 63928 800 64048
rect 0 63248 800 63368
rect 0 62568 800 62688
rect 0 61888 800 62008
rect 0 61208 800 61328
rect 0 60528 800 60648
rect 0 59848 800 59968
rect 0 59168 800 59288
rect 0 58488 800 58608
rect 0 57808 800 57928
rect 0 57128 800 57248
rect 0 56448 800 56568
rect 0 55768 800 55888
rect 0 55088 800 55208
rect 0 54408 800 54528
rect 0 53728 800 53848
rect 0 53048 800 53168
rect 0 52368 800 52488
rect 0 51688 800 51808
rect 0 51008 800 51128
rect 0 50328 800 50448
rect 0 49648 800 49768
rect 0 48968 800 49088
rect 0 48288 800 48408
rect 0 47608 800 47728
rect 0 46928 800 47048
rect 0 46248 800 46368
rect 0 45568 800 45688
rect 0 44888 800 45008
rect 0 44208 800 44328
rect 0 43528 800 43648
rect 0 42848 800 42968
rect 0 42168 800 42288
rect 0 41488 800 41608
rect 0 40808 800 40928
rect 0 40128 800 40248
rect 0 39448 800 39568
rect 0 38768 800 38888
rect 0 38088 800 38208
rect 0 37408 800 37528
rect 0 36728 800 36848
rect 0 36048 800 36168
rect 0 35368 800 35488
rect 0 34688 800 34808
rect 0 34008 800 34128
rect 0 33328 800 33448
rect 0 32648 800 32768
rect 0 31968 800 32088
rect 0 31288 800 31408
rect 0 30608 800 30728
rect 0 29928 800 30048
rect 0 29248 800 29368
rect 0 28568 800 28688
rect 0 27888 800 28008
<< obsm3 >>
rect 749 126688 126027 127941
rect 880 126408 126027 126688
rect 749 84528 126027 126408
rect 880 84248 126027 84528
rect 749 83848 126027 84248
rect 880 83568 126027 83848
rect 749 83168 126027 83568
rect 880 82888 126027 83168
rect 749 82488 126027 82888
rect 880 82208 126027 82488
rect 749 81808 126027 82208
rect 880 81528 126027 81808
rect 749 81128 126027 81528
rect 880 80848 126027 81128
rect 749 80448 126027 80848
rect 880 80168 126027 80448
rect 749 79768 126027 80168
rect 880 79488 126027 79768
rect 749 79088 126027 79488
rect 880 78808 126027 79088
rect 749 78408 126027 78808
rect 880 78128 126027 78408
rect 749 77728 126027 78128
rect 880 77448 126027 77728
rect 749 77048 126027 77448
rect 880 76768 126027 77048
rect 749 76368 126027 76768
rect 880 76088 126027 76368
rect 749 75688 126027 76088
rect 880 75408 126027 75688
rect 749 75008 126027 75408
rect 880 74728 126027 75008
rect 749 74328 126027 74728
rect 880 74048 126027 74328
rect 749 73648 126027 74048
rect 880 73368 126027 73648
rect 749 72968 126027 73368
rect 880 72688 126027 72968
rect 749 72288 126027 72688
rect 880 72008 126027 72288
rect 749 71608 126027 72008
rect 880 71328 126027 71608
rect 749 70928 126027 71328
rect 880 70648 126027 70928
rect 749 70248 126027 70648
rect 880 69968 126027 70248
rect 749 69568 126027 69968
rect 880 69288 126027 69568
rect 749 68888 126027 69288
rect 880 68608 126027 68888
rect 749 68208 126027 68608
rect 880 67928 126027 68208
rect 749 67528 126027 67928
rect 880 67248 126027 67528
rect 749 66848 126027 67248
rect 880 66568 126027 66848
rect 749 66168 126027 66568
rect 880 65888 126027 66168
rect 749 65488 126027 65888
rect 880 65208 126027 65488
rect 749 64808 126027 65208
rect 880 64528 126027 64808
rect 749 64128 126027 64528
rect 880 63848 126027 64128
rect 749 63448 126027 63848
rect 880 63168 126027 63448
rect 749 62768 126027 63168
rect 880 62488 126027 62768
rect 749 62088 126027 62488
rect 880 61808 126027 62088
rect 749 61408 126027 61808
rect 880 61128 126027 61408
rect 749 60728 126027 61128
rect 880 60448 126027 60728
rect 749 60048 126027 60448
rect 880 59768 126027 60048
rect 749 59368 126027 59768
rect 880 59088 126027 59368
rect 749 58688 126027 59088
rect 880 58408 126027 58688
rect 749 58008 126027 58408
rect 880 57728 126027 58008
rect 749 57328 126027 57728
rect 880 57048 126027 57328
rect 749 56648 126027 57048
rect 880 56368 126027 56648
rect 749 55968 126027 56368
rect 880 55688 126027 55968
rect 749 55288 126027 55688
rect 880 55008 126027 55288
rect 749 54608 126027 55008
rect 880 54328 126027 54608
rect 749 53928 126027 54328
rect 880 53648 126027 53928
rect 749 53248 126027 53648
rect 880 52968 126027 53248
rect 749 52568 126027 52968
rect 880 52288 126027 52568
rect 749 51888 126027 52288
rect 880 51608 126027 51888
rect 749 51208 126027 51608
rect 880 50928 126027 51208
rect 749 50528 126027 50928
rect 880 50248 126027 50528
rect 749 49848 126027 50248
rect 880 49568 126027 49848
rect 749 49168 126027 49568
rect 880 48888 126027 49168
rect 749 48488 126027 48888
rect 880 48208 126027 48488
rect 749 47808 126027 48208
rect 880 47528 126027 47808
rect 749 47128 126027 47528
rect 880 46848 126027 47128
rect 749 46448 126027 46848
rect 880 46168 126027 46448
rect 749 45768 126027 46168
rect 880 45488 126027 45768
rect 749 45088 126027 45488
rect 880 44808 126027 45088
rect 749 44408 126027 44808
rect 880 44128 126027 44408
rect 749 43728 126027 44128
rect 880 43448 126027 43728
rect 749 43048 126027 43448
rect 880 42768 126027 43048
rect 749 42368 126027 42768
rect 880 42088 126027 42368
rect 749 41688 126027 42088
rect 880 41408 126027 41688
rect 749 41008 126027 41408
rect 880 40728 126027 41008
rect 749 40328 126027 40728
rect 880 40048 126027 40328
rect 749 39648 126027 40048
rect 880 39368 126027 39648
rect 749 38968 126027 39368
rect 880 38688 126027 38968
rect 749 38288 126027 38688
rect 880 38008 126027 38288
rect 749 37608 126027 38008
rect 880 37328 126027 37608
rect 749 36928 126027 37328
rect 880 36648 126027 36928
rect 749 36248 126027 36648
rect 880 35968 126027 36248
rect 749 35568 126027 35968
rect 880 35288 126027 35568
rect 749 34888 126027 35288
rect 880 34608 126027 34888
rect 749 34208 126027 34608
rect 880 33928 126027 34208
rect 749 33528 126027 33928
rect 880 33248 126027 33528
rect 749 32848 126027 33248
rect 880 32568 126027 32848
rect 749 32168 126027 32568
rect 880 31888 126027 32168
rect 749 31488 126027 31888
rect 880 31208 126027 31488
rect 749 30808 126027 31208
rect 880 30528 126027 30808
rect 749 30128 126027 30528
rect 880 29848 126027 30128
rect 749 29448 126027 29848
rect 880 29168 126027 29448
rect 749 28768 126027 29168
rect 880 28488 126027 28768
rect 749 28088 126027 28488
rect 880 27808 126027 28088
rect 749 2143 126027 27808
<< metal4 >>
rect 4208 2128 4528 127344
rect 4868 2128 5188 127344
rect 34928 2128 35248 127344
rect 35588 2128 35908 127344
rect 65648 2128 65968 127344
rect 66308 2128 66628 127344
rect 96368 2128 96688 127344
rect 97028 2128 97348 127344
<< obsm4 >>
rect 795 127424 124141 127941
rect 795 2211 4128 127424
rect 4608 2211 4788 127424
rect 5268 2211 34848 127424
rect 35328 2211 35508 127424
rect 35988 2211 65568 127424
rect 66048 2211 66228 127424
rect 66708 2211 96288 127424
rect 96768 2211 96948 127424
rect 97428 2211 124141 127424
<< metal5 >>
rect 1056 97914 126456 98234
rect 1056 97254 126456 97574
rect 1056 67278 126456 67598
rect 1056 66618 126456 66938
rect 1056 36642 126456 36962
rect 1056 35982 126456 36302
rect 1056 6006 126456 6326
rect 1056 5346 126456 5666
<< obsm5 >>
rect 13548 67918 122244 69180
rect 13548 37282 122244 66298
rect 13548 13100 122244 35662
<< labels >>
rlabel metal4 s 4868 2128 5188 127344 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 127344 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 127344 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97028 2128 97348 127344 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 126456 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 126456 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67278 126456 67598 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 97914 126456 98234 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 127344 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 127344 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 127344 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 127344 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 126456 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 126456 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 126456 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97254 126456 97574 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 126488 800 126608 6 clock
port 3 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 io_fetch_address[0]
port 4 nsew signal output
rlabel metal2 s 81806 128921 81862 129721 6 io_fetch_address[10]
port 5 nsew signal output
rlabel metal2 s 83738 128921 83794 129721 6 io_fetch_address[11]
port 6 nsew signal output
rlabel metal2 s 81162 128921 81218 129721 6 io_fetch_address[12]
port 7 nsew signal output
rlabel metal2 s 79230 128921 79286 129721 6 io_fetch_address[13]
port 8 nsew signal output
rlabel metal2 s 76010 128921 76066 129721 6 io_fetch_address[14]
port 9 nsew signal output
rlabel metal2 s 82450 128921 82506 129721 6 io_fetch_address[15]
port 10 nsew signal output
rlabel metal2 s 75366 128921 75422 129721 6 io_fetch_address[16]
port 11 nsew signal output
rlabel metal2 s 80518 128921 80574 129721 6 io_fetch_address[17]
port 12 nsew signal output
rlabel metal2 s 68282 128921 68338 129721 6 io_fetch_address[18]
port 13 nsew signal output
rlabel metal2 s 73434 128921 73490 129721 6 io_fetch_address[19]
port 14 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 io_fetch_address[1]
port 15 nsew signal output
rlabel metal2 s 74722 128921 74778 129721 6 io_fetch_address[20]
port 16 nsew signal output
rlabel metal2 s 76654 128921 76710 129721 6 io_fetch_address[21]
port 17 nsew signal output
rlabel metal2 s 77298 128921 77354 129721 6 io_fetch_address[22]
port 18 nsew signal output
rlabel metal2 s 83094 128921 83150 129721 6 io_fetch_address[23]
port 19 nsew signal output
rlabel metal2 s 77942 128921 77998 129721 6 io_fetch_address[24]
port 20 nsew signal output
rlabel metal2 s 90178 128921 90234 129721 6 io_fetch_address[25]
port 21 nsew signal output
rlabel metal2 s 79874 128921 79930 129721 6 io_fetch_address[26]
port 22 nsew signal output
rlabel metal2 s 68926 128921 68982 129721 6 io_fetch_address[27]
port 23 nsew signal output
rlabel metal2 s 78586 128921 78642 129721 6 io_fetch_address[28]
port 24 nsew signal output
rlabel metal2 s 72790 128921 72846 129721 6 io_fetch_address[29]
port 25 nsew signal output
rlabel metal2 s 45098 128921 45154 129721 6 io_fetch_address[2]
port 26 nsew signal output
rlabel metal2 s 72146 128921 72202 129721 6 io_fetch_address[30]
port 27 nsew signal output
rlabel metal2 s 71502 128921 71558 129721 6 io_fetch_address[31]
port 28 nsew signal output
rlabel metal2 s 44454 128921 44510 129721 6 io_fetch_address[3]
port 29 nsew signal output
rlabel metal2 s 43810 128921 43866 129721 6 io_fetch_address[4]
port 30 nsew signal output
rlabel metal2 s 45742 128921 45798 129721 6 io_fetch_address[5]
port 31 nsew signal output
rlabel metal2 s 86958 128921 87014 129721 6 io_fetch_address[6]
port 32 nsew signal output
rlabel metal2 s 70858 128921 70914 129721 6 io_fetch_address[7]
port 33 nsew signal output
rlabel metal2 s 70214 128921 70270 129721 6 io_fetch_address[8]
port 34 nsew signal output
rlabel metal2 s 69570 128921 69626 129721 6 io_fetch_address[9]
port 35 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 io_fetch_data[0]
port 36 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 io_fetch_data[10]
port 37 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 io_fetch_data[11]
port 38 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 io_fetch_data[12]
port 39 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 io_fetch_data[13]
port 40 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 io_fetch_data[14]
port 41 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 io_fetch_data[15]
port 42 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 io_fetch_data[16]
port 43 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 io_fetch_data[17]
port 44 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 io_fetch_data[18]
port 45 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 io_fetch_data[19]
port 46 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 io_fetch_data[1]
port 47 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 io_fetch_data[20]
port 48 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 io_fetch_data[21]
port 49 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 io_fetch_data[22]
port 50 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 io_fetch_data[23]
port 51 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 io_fetch_data[24]
port 52 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 io_fetch_data[25]
port 53 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 io_fetch_data[26]
port 54 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 io_fetch_data[27]
port 55 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 io_fetch_data[28]
port 56 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 io_fetch_data[29]
port 57 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 io_fetch_data[2]
port 58 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 io_fetch_data[30]
port 59 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 io_fetch_data[31]
port 60 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 io_fetch_data[3]
port 61 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 io_fetch_data[4]
port 62 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 io_fetch_data[5]
port 63 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 io_fetch_data[6]
port 64 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 io_fetch_data[7]
port 65 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 io_fetch_data[8]
port 66 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 io_fetch_data[9]
port 67 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 io_load_store_unsigned
port 68 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 io_meip
port 69 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 io_memory_address[0]
port 70 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 io_memory_address[10]
port 71 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 io_memory_address[11]
port 72 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 io_memory_address[12]
port 73 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 io_memory_address[13]
port 74 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 io_memory_address[14]
port 75 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 io_memory_address[15]
port 76 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 io_memory_address[16]
port 77 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 io_memory_address[17]
port 78 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 io_memory_address[18]
port 79 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 io_memory_address[19]
port 80 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 io_memory_address[1]
port 81 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 io_memory_address[20]
port 82 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 io_memory_address[21]
port 83 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 io_memory_address[22]
port 84 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 io_memory_address[23]
port 85 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 io_memory_address[24]
port 86 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 io_memory_address[25]
port 87 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_memory_address[26]
port 88 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 io_memory_address[27]
port 89 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 io_memory_address[28]
port 90 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 io_memory_address[29]
port 91 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 io_memory_address[2]
port 92 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 io_memory_address[30]
port 93 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 io_memory_address[31]
port 94 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 io_memory_address[3]
port 95 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 io_memory_address[4]
port 96 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 io_memory_address[5]
port 97 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 io_memory_address[6]
port 98 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 io_memory_address[7]
port 99 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 io_memory_address[8]
port 100 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 io_memory_address[9]
port 101 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 io_memory_read
port 102 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 io_memory_read_data[0]
port 103 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 io_memory_read_data[10]
port 104 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 io_memory_read_data[11]
port 105 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 io_memory_read_data[12]
port 106 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 io_memory_read_data[13]
port 107 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 io_memory_read_data[14]
port 108 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 io_memory_read_data[15]
port 109 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 io_memory_read_data[16]
port 110 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 io_memory_read_data[17]
port 111 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 io_memory_read_data[18]
port 112 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 io_memory_read_data[19]
port 113 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 io_memory_read_data[1]
port 114 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 io_memory_read_data[20]
port 115 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 io_memory_read_data[21]
port 116 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 io_memory_read_data[22]
port 117 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 io_memory_read_data[23]
port 118 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 io_memory_read_data[24]
port 119 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 io_memory_read_data[25]
port 120 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 io_memory_read_data[26]
port 121 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 io_memory_read_data[27]
port 122 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 io_memory_read_data[28]
port 123 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 io_memory_read_data[29]
port 124 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 io_memory_read_data[2]
port 125 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 io_memory_read_data[30]
port 126 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 io_memory_read_data[31]
port 127 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 io_memory_read_data[3]
port 128 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 io_memory_read_data[4]
port 129 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 io_memory_read_data[5]
port 130 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 io_memory_read_data[6]
port 131 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 io_memory_read_data[7]
port 132 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 io_memory_read_data[8]
port 133 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 io_memory_read_data[9]
port 134 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 io_memory_size[0]
port 135 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 io_memory_size[1]
port 136 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 io_memory_write
port 137 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 io_memory_write_data[0]
port 138 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 io_memory_write_data[10]
port 139 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 io_memory_write_data[11]
port 140 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 io_memory_write_data[12]
port 141 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 io_memory_write_data[13]
port 142 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 io_memory_write_data[14]
port 143 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 io_memory_write_data[15]
port 144 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 io_memory_write_data[16]
port 145 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 io_memory_write_data[17]
port 146 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 io_memory_write_data[18]
port 147 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 io_memory_write_data[19]
port 148 nsew signal output
rlabel metal2 s 74078 128921 74134 129721 6 io_memory_write_data[1]
port 149 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 io_memory_write_data[20]
port 150 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_memory_write_data[21]
port 151 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 io_memory_write_data[22]
port 152 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 io_memory_write_data[23]
port 153 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 io_memory_write_data[24]
port 154 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 io_memory_write_data[25]
port 155 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 io_memory_write_data[26]
port 156 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 io_memory_write_data[27]
port 157 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 io_memory_write_data[28]
port 158 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 io_memory_write_data[29]
port 159 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_memory_write_data[2]
port 160 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 io_memory_write_data[30]
port 161 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 io_memory_write_data[31]
port 162 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 io_memory_write_data[3]
port 163 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 io_memory_write_data[4]
port 164 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 io_memory_write_data[5]
port 165 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 io_memory_write_data[6]
port 166 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 io_memory_write_data[7]
port 167 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 io_memory_write_data[8]
port 168 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 io_memory_write_data[9]
port 169 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 reset
port 170 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 127577 129721
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 54278544
string GDS_FILE /openlane/designs/core/runs/core/results/signoff/core.magic.gds
string GDS_START 1698900
<< end >>

