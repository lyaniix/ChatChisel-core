* NGSPICE file created from core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

.subckt core VGND VPWR clock io_fetch_address[0] io_fetch_address[10] io_fetch_address[11]
+ io_fetch_address[12] io_fetch_address[13] io_fetch_address[14] io_fetch_address[15]
+ io_fetch_address[16] io_fetch_address[17] io_fetch_address[18] io_fetch_address[19]
+ io_fetch_address[1] io_fetch_address[20] io_fetch_address[21] io_fetch_address[22]
+ io_fetch_address[23] io_fetch_address[24] io_fetch_address[25] io_fetch_address[26]
+ io_fetch_address[27] io_fetch_address[28] io_fetch_address[29] io_fetch_address[2]
+ io_fetch_address[30] io_fetch_address[31] io_fetch_address[3] io_fetch_address[4]
+ io_fetch_address[5] io_fetch_address[6] io_fetch_address[7] io_fetch_address[8]
+ io_fetch_address[9] io_fetch_data[0] io_fetch_data[10] io_fetch_data[11] io_fetch_data[12]
+ io_fetch_data[13] io_fetch_data[14] io_fetch_data[15] io_fetch_data[16] io_fetch_data[17]
+ io_fetch_data[18] io_fetch_data[19] io_fetch_data[1] io_fetch_data[20] io_fetch_data[21]
+ io_fetch_data[22] io_fetch_data[23] io_fetch_data[24] io_fetch_data[25] io_fetch_data[26]
+ io_fetch_data[27] io_fetch_data[28] io_fetch_data[29] io_fetch_data[2] io_fetch_data[30]
+ io_fetch_data[31] io_fetch_data[3] io_fetch_data[4] io_fetch_data[5] io_fetch_data[6]
+ io_fetch_data[7] io_fetch_data[8] io_fetch_data[9] io_load_store_unsigned io_meip
+ io_memory_address[0] io_memory_address[10] io_memory_address[11] io_memory_address[12]
+ io_memory_address[13] io_memory_address[14] io_memory_address[15] io_memory_address[16]
+ io_memory_address[17] io_memory_address[18] io_memory_address[19] io_memory_address[1]
+ io_memory_address[20] io_memory_address[21] io_memory_address[22] io_memory_address[23]
+ io_memory_address[24] io_memory_address[25] io_memory_address[26] io_memory_address[27]
+ io_memory_address[28] io_memory_address[29] io_memory_address[2] io_memory_address[30]
+ io_memory_address[31] io_memory_address[3] io_memory_address[4] io_memory_address[5]
+ io_memory_address[6] io_memory_address[7] io_memory_address[8] io_memory_address[9]
+ io_memory_read io_memory_read_data[0] io_memory_read_data[10] io_memory_read_data[11]
+ io_memory_read_data[12] io_memory_read_data[13] io_memory_read_data[14] io_memory_read_data[15]
+ io_memory_read_data[16] io_memory_read_data[17] io_memory_read_data[18] io_memory_read_data[19]
+ io_memory_read_data[1] io_memory_read_data[20] io_memory_read_data[21] io_memory_read_data[22]
+ io_memory_read_data[23] io_memory_read_data[24] io_memory_read_data[25] io_memory_read_data[26]
+ io_memory_read_data[27] io_memory_read_data[28] io_memory_read_data[29] io_memory_read_data[2]
+ io_memory_read_data[30] io_memory_read_data[31] io_memory_read_data[3] io_memory_read_data[4]
+ io_memory_read_data[5] io_memory_read_data[6] io_memory_read_data[7] io_memory_read_data[8]
+ io_memory_read_data[9] io_memory_size[0] io_memory_size[1] io_memory_write io_memory_write_data[0]
+ io_memory_write_data[10] io_memory_write_data[11] io_memory_write_data[12] io_memory_write_data[13]
+ io_memory_write_data[14] io_memory_write_data[15] io_memory_write_data[16] io_memory_write_data[17]
+ io_memory_write_data[18] io_memory_write_data[19] io_memory_write_data[1] io_memory_write_data[20]
+ io_memory_write_data[21] io_memory_write_data[22] io_memory_write_data[23] io_memory_write_data[24]
+ io_memory_write_data[25] io_memory_write_data[26] io_memory_write_data[27] io_memory_write_data[28]
+ io_memory_write_data[29] io_memory_write_data[2] io_memory_write_data[30] io_memory_write_data[31]
+ io_memory_write_data[3] io_memory_write_data[4] io_memory_write_data[5] io_memory_write_data[6]
+ io_memory_write_data[7] io_memory_write_data[8] io_memory_write_data[9] reset
XFILLER_0_193_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18869_ _04167_ _04165_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__nand2_2
XFILLER_0_222_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20900_ _05929_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21880_ _06525_ _06519_ _06520_ _06526_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20831_ net102 _05891_ _05887_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23550_ net223 _07917_ _07919_ _07907_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__o211a_1
X_20762_ _03452_ _05425_ csr.io_csr_address\[8\] VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__and3b_1
XFILLER_0_65_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22501_ net67 _07065_ _07093_ _07095_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23481_ net18 _07875_ _07878_ _07879_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20693_ _03728_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25220_ _08839_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__clkbuf_1
X_22432_ fetch.bht.bhtTable_tag\[12\]\[12\] fetch.bht.bhtTable_tag\[13\]\[12\] _06616_
+ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_350_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_350_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25151_ _08803_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__clkbuf_1
X_22363_ fetch.bht.bhtTable_tag\[4\]\[2\] fetch.bht.bhtTable_tag\[5\]\[2\] fetch.bht.bhtTable_tag\[6\]\[2\]
+ fetch.bht.bhtTable_tag\[7\]\[2\] _06679_ _06620_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__mux4_2
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24102_ net829 execute.io_target_pc\[6\] _08221_ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__mux2_1
X_21314_ net1284 _10807_ _06157_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25082_ net2800 _08712_ _08646_ csr.mcycle\[31\] VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__a211oi_1
X_22294_ net69 _06794_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24033_ _08188_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__clkbuf_1
X_28910_ clknet_leaf_87_clock _01923_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_1168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21245_ net1056 _06122_ _06120_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__mux2_1
Xhold340 csr.minstret\[19\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29890_ clknet_leaf_304_clock _02903_ VGND VGND VPWR VPWR decode.regfile.registers_20\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold351 _06317_ VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold362 decode.regfile.registers_22\[12\] VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold373 decode.regfile.registers_31\[21\] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__buf_1
XFILLER_0_102_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28841_ clknet_leaf_88_clock _01854_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold384 decode.regfile.registers_16\[15\] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__dlygate4sd3_1
X_21176_ _06074_ _06082_ net2657 VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__and3_1
Xhold395 decode.regfile.registers_3\[6\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_225_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20127_ _05320_ _05335_ _05327_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__nand3_1
X_28772_ clknet_leaf_131_clock _01785_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25984_ _09287_ _09949_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__nand2_1
X_27723_ clknet_leaf_23_clock _00752_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20058_ _05275_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__xor2_1
X_24935_ csr._mcycle_T_3\[46\] csr._mcycle_T_3\[45\] csr._mcycle_T_3\[44\] _08665_
+ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1040 fetch.bht.bhtTable_tag\[0\]\[0\] VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1051 fetch.bht.bhtTable_target_pc\[6\]\[0\] VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1062 fetch.bht.bhtTable_tag\[5\]\[9\] VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27654_ clknet_leaf_48_clock _00683_ VGND VGND VPWR VPWR execute.io_reg_pc\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_24866_ _06145_ net1407 _08388_ VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1073 decode.regfile.registers_3\[7\] VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 fetch.bht.bhtTable_target_pc\[15\]\[9\] VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 fetch.bht.bhtTable_target_pc\[3\]\[16\] VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26605_ net2518 _09649_ _09657_ _09648_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__o211a_1
X_23817_ _08065_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_303_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_303_clock
+ sky130_fd_sc_hd__clkbuf_8
X_27585_ clknet_leaf_136_clock _00614_ VGND VGND VPWR VPWR csr.io_mem_pc\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24797_ _08561_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_155_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29324_ clknet_leaf_226_clock _02337_ VGND VGND VPWR VPWR decode.regfile.registers_2\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14550_ _10592_ VGND VGND VPWR VPWR _10593_ sky130_fd_sc_hd__clkbuf_4
X_26536_ net1271 _09579_ _09617_ _09608_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23748_ _08025_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_81_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13501_ _09882_ VGND VGND VPWR VPWR _09883_ sky130_fd_sc_hd__buf_2
XFILLER_0_138_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29255_ clknet_leaf_233_clock _02268_ VGND VGND VPWR VPWR decode.regfile.registers_0\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26467_ _09577_ VGND VGND VPWR VPWR _09579_ sky130_fd_sc_hd__buf_2
X_14481_ net600 _10533_ _10536_ _10535_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__o211a_1
X_23679_ _07988_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28206_ clknet_leaf_63_clock net1734 VGND VGND VPWR VPWR csr.mscratch\[8\] sky130_fd_sc_hd__dfxtp_1
X_16220_ decode.regfile.registers_20\[23\] _11103_ _11222_ _12193_ VGND VGND VPWR
+ VPWR _12194_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25418_ net193 VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_318_clock clknet_5_18__leaf_clock VGND VGND VPWR VPWR clknet_leaf_318_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_192_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29186_ clknet_leaf_239_clock _02199_ VGND VGND VPWR VPWR fetch.btb.btbTable\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_26398_ _09379_ _09535_ VGND VGND VPWR VPWR _09539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28137_ clknet_leaf_212_clock _01159_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16151_ decode.regfile.registers_25\[21\] _11483_ _11484_ decode.regfile.registers_24\[21\]
+ VGND VGND VPWR VPWR _12127_ sky130_fd_sc_hd__o22a_1
XFILLER_0_148_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25349_ net792 _08906_ _08908_ _07247_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_114_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer7 net232 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15102_ _11098_ VGND VGND VPWR VPWR _11099_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_79_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28068_ clknet_leaf_183_clock _01090_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_16082_ _11117_ _11057_ _11109_ decode.regfile.registers_0\[20\] VGND VGND VPWR VPWR
+ _12059_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_185_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15033_ net677 _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__a31o_1
X_27019_ clknet_leaf_338_clock _00048_ VGND VGND VPWR VPWR decode.regfile.registers_22\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19910_ _05178_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19841_ _03705_ _04305_ _04751_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19772_ _05026_ _03851_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__nand2_1
X_16984_ _12931_ _12943_ _12607_ VGND VGND VPWR VPWR _12944_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_88_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15935_ _11154_ decode.regfile.registers_0\[16\] _11156_ _11915_ VGND VGND VPWR VPWR
+ _11916_ sky130_fd_sc_hd__a211o_1
X_18723_ _04014_ _04021_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__nor2_2
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18654_ decode.id_ex_rs2_data_reg\[20\] _03746_ _03949_ _03952_ VGND VGND VPWR VPWR
+ _03953_ sky130_fd_sc_hd__o211ai_4
X_15866_ _11841_ _11848_ _11136_ VGND VGND VPWR VPWR _11849_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_189_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14817_ _10770_ _10859_ VGND VGND VPWR VPWR _10860_ sky130_fd_sc_hd__nand2_1
X_17605_ decode.regfile.registers_11\[20\] _12594_ _03010_ _03011_ _12794_ VGND VGND
+ VPWR VPWR _03012_ sky130_fd_sc_hd__a221o_1
X_18585_ _03659_ execute.csr_read_data_out_reg\[22\] execute.io_reg_pc\[22\] _03777_
+ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15797_ _11199_ _11780_ _11781_ VGND VGND VPWR VPWR _11782_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17536_ _13407_ decode.regfile.registers_25\[18\] _13482_ _13294_ VGND VGND VPWR
+ VPWR _13483_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14748_ csr.io_mem_pc\[24\] _10768_ csr.io_mem_pc\[25\] VGND VGND VPWR VPWR _10791_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_103_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17467_ _13055_ net1324 _13097_ VGND VGND VPWR VPWR _13415_ sky130_fd_sc_hd__o21a_1
X_14679_ _10721_ execute.io_target_pc\[10\] _10720_ execute.io_target_pc\[26\] VGND
+ VGND VPWR VPWR _10722_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_11_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19206_ _04494_ _04496_ _04445_ _04501_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__a211o_1
X_16418_ decode.regfile.registers_3\[29\] _11110_ _11141_ _11146_ VGND VGND VPWR VPWR
+ _12386_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17398_ decode.regfile.registers_6\[15\] _12880_ _13342_ _13347_ VGND VGND VPWR VPWR
+ _13348_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_55_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19137_ _04255_ _04070_ _04251_ _04252_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16349_ decode.regfile.registers_4\[27\] _10636_ _11410_ _12314_ _12318_ VGND VGND
+ VPWR VPWR _12319_ sky130_fd_sc_hd__o32a_1
XFILLER_0_15_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19068_ _03772_ net194 _03775_ _03780_ _03988_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_140_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18019_ decode.regfile.registers_2\[31\] _12882_ _12729_ VGND VGND VPWR VPWR _03415_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21030_ execute.csr_read_data_out_reg\[5\] _05989_ _05998_ VGND VGND VPWR VPWR _06000_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_11_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22981_ _07367_ _07427_ _07428_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__or3b_1
X_24720_ _08544_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__clkbuf_1
X_21932_ _06561_ _06543_ _06544_ _06562_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24651_ net995 execute.io_target_pc\[14\] _08508_ VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__mux2_1
X_21863_ net1733 _06497_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__or2_1
X_23602_ _06132_ net1538 _07941_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27370_ clknet_leaf_29_clock _00399_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_20814_ _05882_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24582_ _09896_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__buf_4
XFILLER_0_166_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21794_ _06457_ net217 _06458_ _06459_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__and4b_1
XFILLER_0_92_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26321_ _09377_ _09492_ VGND VGND VPWR VPWR _09495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23533_ net73 _07903_ _07909_ _07907_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20745_ _05831_ _05813_ decode.id_ex_rs1_data_reg\[29\] _05843_ _00514_ VGND VGND
+ VPWR VPWR _00748_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29040_ clknet_leaf_105_clock _02053_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_189_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26252_ _09383_ _09448_ VGND VGND VPWR VPWR _09455_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_189_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23464_ _11027_ _07862_ _07859_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__or3b_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20676_ _00689_ _05800_ _05801_ _05799_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25203_ net424 _08830_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__xnor2_1
X_22415_ _07008_ _07009_ _06790_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__mux2_1
X_26183_ net1138 _09395_ _09407_ _09394_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__o211a_1
X_23395_ net88 _07706_ _07707_ _07818_ _07705_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__o311a_1
XFILLER_0_33_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25134_ _08795_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22346_ _06940_ _06650_ _06686_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_227_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_227_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_227_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25065_ csr.mcycle\[24\] csr.mcycle\[23\] _08756_ VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__and3_1
X_22277_ fetch.bht.bhtTable_tag\[4\]\[6\] fetch.bht.bhtTable_tag\[5\]\[6\] _06617_
+ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29942_ clknet_leaf_341_clock _02955_ VGND VGND VPWR VPWR decode.regfile.registers_21\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_148_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24016_ _08179_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__clkbuf_1
X_21228_ _10812_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__buf_2
XFILLER_0_218_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold170 io_fetch_data[6] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold181 _10732_ VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29873_ clknet_leaf_299_clock _02886_ VGND VGND VPWR VPWR decode.regfile.registers_19\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_180_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold192 fetch.btb.btbTable\[11\]\[0\] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28824_ clknet_leaf_121_clock _01837_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21159_ _06073_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28755_ clknet_leaf_140_clock _01768_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_13981_ _09970_ _10244_ VGND VGND VPWR VPWR _10248_ sky130_fd_sc_hd__nand2_1
X_25967_ net2525 _09270_ _09276_ _09277_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15720_ decode.regfile.registers_15\[10\] _11037_ _11205_ _11208_ decode.regfile.registers_14\[10\]
+ VGND VGND VPWR VPWR _11707_ sky130_fd_sc_hd__a32o_1
X_27706_ clknet_leaf_22_clock _00735_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_24918_ _07199_ net525 _08659_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_107_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28686_ clknet_leaf_112_clock _01699_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_242_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_242_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25898_ _08970_ _09198_ VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27637_ clknet_leaf_156_clock _00666_ VGND VGND VPWR VPWR execute.io_reg_pc\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ decode.regfile.registers_25\[8\] _11483_ _11484_ decode.regfile.registers_24\[8\]
+ VGND VGND VPWR VPWR _11640_ sky130_fd_sc_hd__o22a_1
X_24849_ _08612_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_178_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_60 _10101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_71 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14602_ decode.immGen._imm_T_24\[4\] VGND VGND VPWR VPWR _10645_ sky130_fd_sc_hd__buf_2
XINSDIODE1_82 _10588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_93 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18370_ decode.id_ex_islui_reg VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__inv_2
X_27568_ clknet_leaf_158_clock _00597_ VGND VGND VPWR VPWR csr.io_mem_pc\[9\] sky130_fd_sc_hd__dfxtp_1
X_15582_ _11571_ net2785 _11039_ _11032_ _11033_ VGND VGND VPWR VPWR _11572_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_84_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29307_ clknet_leaf_244_clock _02320_ VGND VGND VPWR VPWR decode.regfile.registers_2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_17321_ _13268_ _13271_ _13272_ VGND VGND VPWR VPWR _13273_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_51_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14533_ _10575_ VGND VGND VPWR VPWR _10576_ sky130_fd_sc_hd__buf_4
X_26519_ _09424_ _09602_ VGND VGND VPWR VPWR _09609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_257_clock clknet_5_22__leaf_clock VGND VGND VPWR VPWR clknet_leaf_257_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_166_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27499_ clknet_leaf_33_clock _00528_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29238_ clknet_leaf_177_clock _02251_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_17252_ decode.regfile.registers_21\[11\] _12822_ _13184_ _13205_ _12806_ VGND VGND
+ VPWR VPWR _13206_ sky130_fd_sc_hd__o221a_1
X_14464_ net431 _10520_ _10526_ _10522_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_137_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ _11154_ decode.regfile.registers_0\[23\] _11156_ _12176_ VGND VGND VPWR VPWR
+ _12177_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29169_ clknet_leaf_191_clock _02182_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17183_ _13055_ decode.regfile.registers_30\[10\] _13097_ VGND VGND VPWR VPWR _13138_
+ sky130_fd_sc_hd__o21a_1
X_14395_ net1324 _10477_ _10486_ _10481_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_77_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16134_ decode.regfile.registers_7\[21\] _11378_ _11170_ decode.regfile.registers_6\[21\]
+ _11166_ VGND VGND VPWR VPWR _12110_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_148_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16065_ decode.regfile.registers_20\[19\] _11102_ _12041_ _12042_ _11327_ VGND VGND
+ VPWR VPWR _12043_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15016_ _11025_ VGND VGND VPWR VPWR _11026_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19824_ _04618_ _04589_ _05090_ _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_36_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1809 fetch.bht.bhtTable_tag\[6\]\[19\] VGND VGND VPWR VPWR net2036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19755_ _03847_ _04442_ _04444_ _03851_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16967_ _12533_ VGND VGND VPWR VPWR _12927_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18706_ _09963_ net230 net232 VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__nand3_2
XFILLER_0_194_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15918_ decode.regfile.registers_18\[15\] _11455_ _11898_ _11899_ _11456_ VGND VGND
+ VPWR VPWR _11900_ sky130_fd_sc_hd__a221o_1
X_16898_ decode.regfile.registers_22\[3\] _12528_ _12859_ _12687_ VGND VGND VPWR VPWR
+ _12860_ sky130_fd_sc_hd__a211o_1
X_19686_ _03944_ net190 _04253_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__mux2_1
X_15849_ _11761_ net409 _11796_ _11832_ _11760_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__o221a_1
X_18637_ _03929_ _03933_ _03934_ _03935_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_204_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18568_ _03791_ _03803_ _03830_ _03866_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17519_ decode.regfile.registers_10\[18\] _12654_ _12878_ _13465_ VGND VGND VPWR
+ VPWR _13466_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18499_ net239 _03797_ net191 VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__or3b_1
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20530_ csr.mcycle\[12\] _05552_ _05676_ _05677_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20461_ _03718_ _05516_ _05528_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__and3_2
XFILLER_0_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22200_ net87 VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__buf_4
XFILLER_0_171_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23180_ execute.io_target_pc\[16\] _05864_ _07091_ _07616_ _07347_ VGND VGND VPWR
+ VPWR _07617_ sky130_fd_sc_hd__a311o_1
XFILLER_0_144_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20392_ _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_207_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22131_ fetch.bht.bhtTable_tag\[12\]\[4\] fetch.bht.bhtTable_tag\[13\]\[4\] _06706_
+ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22062_ fetch.bht.bhtTable_tag\[0\]\[18\] fetch.bht.bhtTable_tag\[1\]\[18\] fetch.bht.bhtTable_tag\[2\]\[18\]
+ fetch.bht.bhtTable_tag\[3\]\[18\] _06646_ _06652_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__mux4_1
XFILLER_0_218_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21013_ execute.io_reg_pc\[30\] _05989_ _05985_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_222_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26870_ _09398_ _09806_ VGND VGND VPWR VPWR _09811_ sky130_fd_sc_hd__nand2_1
X_25821_ net2512 _09183_ _09192_ _09182_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28540_ clknet_leaf_211_clock _01553_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_25752_ _09128_ VGND VGND VPWR VPWR _09153_ sky130_fd_sc_hd__clkbuf_4
X_22964_ _07391_ _07392_ _07411_ _07412_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__o2bb2a_1
X_24703_ _08535_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21915_ csr.io_mret_vector\[23\] csr.io_mem_pc\[23\] _06539_ VGND VGND VPWR VPWR
+ _06551_ sky130_fd_sc_hd__mux2_1
X_28471_ clknet_leaf_148_clock _01484_ VGND VGND VPWR VPWR decode.io_id_pc\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25683_ _08982_ _09112_ VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__nand2_1
X_22895_ _06032_ _07345_ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__nor2_2
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27422_ clknet_leaf_28_clock _00451_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[31\]
+ sky130_fd_sc_hd__dfxtp_2
X_24634_ net1323 execute.io_target_pc\[6\] _08497_ VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21846_ _06501_ _06494_ _06495_ _06502_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27353_ clknet_leaf_47_clock _00382_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[26\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_216_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24565_ _08464_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_216_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21777_ net1268 _10759_ _06450_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26304_ net680 _09475_ _09483_ _09484_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__o211a_1
X_23516_ net2471 _07890_ _07887_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__or3b_1
XFILLER_0_148_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1086 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27284_ clknet_leaf_33_clock _00313_ VGND VGND VPWR VPWR decode.regfile.registers_31\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20728_ _03728_ decode.id_ex_rs1_data_reg\[22\] VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24496_ _08055_ net1361 _08428_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29023_ clknet_leaf_180_clock _02036_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26235_ _09443_ _09372_ VGND VGND VPWR VPWR _09444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23447_ net4 _07846_ _07858_ _07851_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__o211a_1
X_20659_ csr.io_mret_vector\[31\] _05580_ _05581_ csr.mscratch\[31\] _05787_ VGND
+ VGND VPWR VPWR _05788_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14180_ net2420 _10359_ _10362_ _10357_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__o211a_1
X_26166_ _10030_ VGND VGND VPWR VPWR _09396_ sky130_fd_sc_hd__buf_4
X_23378_ csr._csr_read_data_T_8\[28\] _07416_ _07790_ _07801_ _07802_ VGND VGND VPWR
+ VPWR _07803_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25117_ _06134_ net1793 _08778_ VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22329_ _06790_ _06923_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26097_ _08943_ _09340_ VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_72_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25048_ _06331_ _08744_ _08745_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__nor3_1
X_29925_ clknet_leaf_337_clock _02938_ VGND VGND VPWR VPWR decode.regfile.registers_21\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_167_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17870_ _10614_ decode.regfile.registers_2\[27\] VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_109_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29856_ clknet_leaf_305_clock _02869_ VGND VGND VPWR VPWR decode.regfile.registers_19\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28807_ clknet_leaf_119_clock _01820_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16821_ decode.regfile.registers_4\[2\] _12618_ _12620_ decode.regfile.registers_5\[2\]
+ _12737_ VGND VGND VPWR VPWR _12784_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_181_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_181_clock
+ sky130_fd_sc_hd__clkbuf_8
X_26999_ clknet_leaf_337_clock _00028_ VGND VGND VPWR VPWR decode.regfile.registers_22\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_29787_ clknet_leaf_309_clock _02800_ VGND VGND VPWR VPWR decode.regfile.registers_17\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_21_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16752_ _12681_ VGND VGND VPWR VPWR _12716_ sky130_fd_sc_hd__clkbuf_4
X_19540_ _04095_ _04820_ _04822_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__a211o_1
X_28738_ clknet_leaf_135_clock _01751_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13964_ net2407 _10226_ _10236_ _10232_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15703_ _11689_ VGND VGND VPWR VPWR _11690_ sky130_fd_sc_hd__clkbuf_4
X_28669_ clknet_leaf_177_clock _01682_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16683_ decode.regfile.registers_9\[0\] _12603_ _12608_ _12647_ VGND VGND VPWR VPWR
+ _12648_ sky130_fd_sc_hd__o22a_1
X_19471_ _04745_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__nand2_1
X_13895_ decode.io_wb_rd\[0\] decode.io_wb_rd\[1\] VGND VGND VPWR VPWR _10196_ sky130_fd_sc_hd__nor2_8
XFILLER_0_115_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15634_ _11136_ _11621_ _11622_ _11166_ VGND VGND VPWR VPWR _11623_ sky130_fd_sc_hd__a211o_1
X_18422_ csr.io_csr_address\[0\] VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__clkinv_4
Xclkbuf_leaf_196_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_196_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_303 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_314 decode.regfile.registers_10\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_325 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_336 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_347 _03580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18353_ decode.id_ex_ex_rs1_reg\[4\] VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__inv_2
X_15565_ decode.regfile.registers_18\[6\] _10642_ _11112_ _10652_ _10633_ VGND VGND
+ VPWR VPWR _11556_ sky130_fd_sc_hd__o2111a_1
XINSDIODE1_358 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_369 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17304_ _13091_ _13176_ decode.regfile.registers_27\[12\] _13050_ VGND VGND VPWR
+ VPWR _13257_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14516_ fetch.btb.btbTable\[8\]\[0\] fetch.btb.btbTable\[9\]\[0\] fetch.btb.btbTable\[10\]\[0\]
+ fetch.btb.btbTable\[11\]\[0\] _09891_ _09888_ VGND VGND VPWR VPWR _10561_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ decode.id_ex_rs2_data_reg\[8\] _03605_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15496_ _11238_ VGND VGND VPWR VPWR _11489_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_61_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17235_ decode.regfile.registers_11\[11\] _12724_ _12587_ _12550_ VGND VGND VPWR
+ VPWR _13189_ sky130_fd_sc_hd__a22o_1
X_14447_ net434 _10506_ _10516_ _10509_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17166_ decode.regfile.registers_17\[9\] _12580_ _12826_ VGND VGND VPWR VPWR _13122_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14378_ _10462_ VGND VGND VPWR VPWR _10477_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold906 decode.regfile.registers_4\[16\] VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 fetch.bht.bhtTable_target_pc\[6\]\[27\] VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__dlygate4sd3_1
X_16117_ _11646_ _11834_ _11944_ decode.regfile.registers_29\[20\] _12093_ VGND VGND
+ VPWR VPWR _12094_ sky130_fd_sc_hd__o221a_1
Xhold928 csr.mcycle\[9\] VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold939 fetch.bht.bhtTable_target_pc\[8\]\[31\] VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_134_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_134_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17097_ net434 _12709_ _13009_ _13054_ _12705_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16048_ decode.regfile.registers_4\[19\] _11375_ _12021_ _12025_ VGND VGND VPWR VPWR
+ _12026_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_161_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2307 csr._csr_read_data_T_8\[14\] VGND VGND VPWR VPWR net2534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2318 decode.regfile.registers_2\[17\] VGND VGND VPWR VPWR net2545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2329 decode.regfile.registers_26\[20\] VGND VGND VPWR VPWR net2556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1606 decode.regfile.registers_14\[20\] VGND VGND VPWR VPWR net1833 sky130_fd_sc_hd__dlygate4sd3_1
X_19807_ _05045_ _05046_ _05049_ _03814_ _03852_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__o2111ai_1
Xclkbuf_leaf_149_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_149_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1617 decode.regfile.registers_10\[7\] VGND VGND VPWR VPWR net1844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1628 fetch.bht.bhtTable_target_pc\[15\]\[21\] VGND VGND VPWR VPWR net1855 sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ decode.regfile.registers_17\[30\] _12719_ _03378_ _03395_ _12826_ VGND VGND
+ VPWR VPWR _03396_ sky130_fd_sc_hd__o221a_1
Xhold1639 decode.regfile.registers_25\[19\] VGND VGND VPWR VPWR net1866 sky130_fd_sc_hd__dlygate4sd3_1
X_19738_ _05004_ _05005_ _05011_ _05013_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_223_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19669_ _04509_ _04550_ _04879_ _04947_ _04595_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__a32o_1
XFILLER_0_177_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21700_ csr.minstret\[17\] csr.minstret\[18\] _06400_ _06401_ VGND VGND VPWR VPWR
+ _06402_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22680_ net2423 _07222_ _07227_ _07221_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21631_ _03580_ _06348_ _06350_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__nor3_1
XFILLER_0_158_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24350_ _08351_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21562_ _06301_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23301_ _07089_ _07726_ _07727_ _07730_ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_211_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20513_ csr.minstret\[10\] _05658_ _05659_ _05662_ _05537_ VGND VGND VPWR VPWR _05663_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24281_ _08109_ net983 _06218_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21493_ _06122_ net1894 _06263_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26020_ _08941_ _09297_ VGND VGND VPWR VPWR _09308_ sky130_fd_sc_hd__nand2_1
X_23232_ _07665_ _07110_ VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__or2b_1
X_20444_ csr._minstret_T_3\[35\] _05577_ _05578_ _05600_ VGND VGND VPWR VPWR _05601_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23163_ _06025_ _07573_ _03546_ _07600_ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__a31o_1
X_20375_ _05526_ _05536_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__nand2_4
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22114_ _06685_ _06708_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__and2b_1
X_27971_ clknet_leaf_216_clock _00993_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_23094_ net69 _07343_ _07344_ _07534_ _07535_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__o311a_1
XFILLER_0_28_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22045_ _00003_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__clkbuf_8
X_29710_ clknet_leaf_283_clock _02723_ VGND VGND VPWR VPWR decode.regfile.registers_14\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_26922_ net2250 _09839_ _09841_ _09836_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29641_ clknet_leaf_277_clock _02654_ VGND VGND VPWR VPWR decode.regfile.registers_12\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_26853_ net896 _09795_ _09801_ _09799_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_162_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25804_ _08952_ _09179_ VGND VGND VPWR VPWR _09184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29572_ clknet_leaf_267_clock _02585_ VGND VGND VPWR VPWR decode.regfile.registers_10\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_26784_ net1420 _09752_ _09761_ _09758_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o211a_1
X_23996_ net1277 VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28523_ clknet_leaf_169_clock _01536_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_218_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25735_ _08958_ _09136_ VGND VGND VPWR VPWR _09144_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_218_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22947_ execute.io_target_pc\[3\] _03592_ _03590_ _07396_ VGND VGND VPWR VPWR _07397_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_206_Right_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28454_ clknet_leaf_148_clock _01467_ VGND VGND VPWR VPWR decode.io_id_pc\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13680_ _10012_ memory.io_wb_aluresult\[11\] _09978_ memory.io_wb_reg_pc\[11\] _09977_
+ VGND VGND VPWR VPWR _10034_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25666_ net2454 _09095_ _09103_ _09100_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_863 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22878_ net1784 _10773_ _07335_ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27405_ clknet_leaf_9_clock _00434_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[14\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_171_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24617_ net868 execute.io_target_pc\[30\] _09897_ VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28385_ clknet_leaf_145_clock _01398_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_4
X_21829_ _06479_ csr._mcycle_T_2\[2\] _06396_ net735 VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25597_ net1142 _09052_ _09063_ _09059_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27336_ clknet_leaf_46_clock _00365_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_15350_ _10962_ decode.regfile.registers_30\[2\] _11039_ _11032_ _11033_ VGND VGND
+ VPWR VPWR _11345_ sky130_fd_sc_hd__o2111a_1
X_24548_ _08455_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14301_ _10025_ _10431_ VGND VGND VPWR VPWR _10433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27267_ clknet_leaf_13_clock _00296_ VGND VGND VPWR VPWR decode.regfile.registers_30\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_15281_ _11035_ _11043_ _11143_ VGND VGND VPWR VPWR _11277_ sky130_fd_sc_hd__and3_1
X_24479_ _08419_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29006_ clknet_leaf_110_clock _02019_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17020_ decode.regfile.registers_10\[6\] _12600_ _12976_ _12978_ _12724_ VGND VGND
+ VPWR VPWR _12979_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_130_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ _10042_ _10387_ VGND VGND VPWR VPWR _10393_ sky130_fd_sc_hd__nand2_1
X_26218_ _10116_ VGND VGND VPWR VPWR _09432_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_51_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_51_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27198_ clknet_leaf_361_clock _00227_ VGND VGND VPWR VPWR decode.regfile.registers_28\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire177 net178 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_169_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14163_ net1305 _10346_ _10352_ _10344_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__o211a_1
X_26149_ _09383_ _09374_ VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_95_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18971_ _04269_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14094_ _10074_ _10312_ VGND VGND VPWR VPWR _10313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_66_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_66_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17922_ decode.regfile.registers_14\[28\] _12984_ _03306_ _03320_ _12874_ VGND VGND
+ VPWR VPWR _03321_ sky130_fd_sc_hd__o221a_1
X_29908_ clknet_leaf_301_clock _02921_ VGND VGND VPWR VPWR decode.regfile.registers_20\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17853_ _12712_ decode.regfile.registers_24\[26\] _12997_ _12998_ _13367_ VGND VGND
+ VPWR VPWR _03254_ sky130_fd_sc_hd__o2111a_1
X_29839_ clknet_leaf_299_clock _02852_ VGND VGND VPWR VPWR decode.regfile.registers_18\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16804_ _12766_ VGND VGND VPWR VPWR _12767_ sky130_fd_sc_hd__buf_2
X_17784_ decode.regfile.registers_20\[25\] _12525_ _12552_ _12823_ _12824_ VGND VGND
+ VPWR VPWR _03186_ sky130_fd_sc_hd__a41o_1
X_14996_ _11008_ VGND VGND VPWR VPWR _11009_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19523_ _04349_ _04273_ _04468_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__and3_1
X_13947_ net2310 _10226_ _10227_ _10219_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__o211a_1
X_16735_ decode.regfile.registers_29\[0\] _12493_ _12496_ decode.regfile.registers_28\[0\]
+ _12699_ VGND VGND VPWR VPWR _12700_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16666_ _12630_ VGND VGND VPWR VPWR _12631_ sky130_fd_sc_hd__buf_4
X_19454_ _04169_ _04637_ _04740_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_198_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13878_ _10112_ _10177_ VGND VGND VPWR VPWR _10186_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_100 _10660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_111 _10994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18405_ _03703_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__clkbuf_4
XINSDIODE1_122 _11085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15617_ _10960_ decode.regfile.registers_28\[7\] _11067_ _11038_ _11440_ VGND VGND
+ VPWR VPWR _11607_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_69_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_133 _11347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19385_ _04393_ _04534_ _04674_ _04371_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16597_ _12561_ VGND VGND VPWR VPWR _12562_ sky130_fd_sc_hd__clkbuf_4
XINSDIODE1_144 _12504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_155 _12690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_166 decode.id_ex_rs1_data_reg\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15548_ _11538_ VGND VGND VPWR VPWR _11539_ sky130_fd_sc_hd__clkbuf_4
X_18336_ decode.id_ex_aluop_reg\[3\] VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__buf_2
XINSDIODE1_177 execute.csr_read_data_out_reg\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_188 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_199 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18267_ _03597_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__clkbuf_1
X_15479_ decode.regfile.registers_10\[4\] _11184_ _11468_ _11469_ _11471_ VGND VGND
+ VPWR VPWR _11472_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_19_clock
+ sky130_fd_sc_hd__clkbuf_8
X_17218_ _12915_ decode.regfile.registers_25\[10\] _13045_ _12812_ VGND VGND VPWR
+ VPWR _13173_ sky130_fd_sc_hd__or4_1
XFILLER_0_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18198_ _10943_ _03528_ decode.control.io_funct7\[5\] VGND VGND VPWR VPWR _03536_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold703 fetch.bht.bhtTable_target_pc\[5\]\[11\] VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 fetch.bht.bhtTable_target_pc\[14\]\[19\] VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17149_ decode.regfile.registers_3\[9\] _12628_ _13102_ _13104_ VGND VGND VPWR VPWR
+ _13105_ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold725 fetch.bht.bhtTable_tag\[12\]\[10\] VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold736 fetch.bht.bhtTable_target_pc\[9\]\[5\] VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold747 fetch.bht.bhtTable_target_pc\[12\]\[8\] VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold758 fetch.bht.bhtTable_tag\[4\]\[9\] VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__dlygate4sd3_1
X_20160_ decode.id_ex_imm_reg\[23\] _10786_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__xor2_1
Xhold769 fetch.bht.bhtTable_target_pc\[8\]\[13\] VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__dlygate4sd3_1
X_20091_ decode.id_ex_imm_reg\[11\] _10689_ _05297_ _05304_ VGND VGND VPWR VPWR _05305_
+ sky130_fd_sc_hd__o211ai_2
Xhold2104 decode.regfile.registers_30\[31\] VGND VGND VPWR VPWR net2331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2115 decode.regfile.registers_11\[11\] VGND VGND VPWR VPWR net2342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2126 decode.regfile.registers_15\[7\] VGND VGND VPWR VPWR net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2137 decode.regfile.registers_8\[28\] VGND VGND VPWR VPWR net2364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1403 _10721_ VGND VGND VPWR VPWR net1630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2148 decode.regfile.registers_12\[23\] VGND VGND VPWR VPWR net2375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 fetch.bht.bhtTable_tag\[14\]\[7\] VGND VGND VPWR VPWR net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2159 _10720_ VGND VGND VPWR VPWR net2386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1425 fetch.bht.bhtTable_target_pc\[14\]\[26\] VGND VGND VPWR VPWR net1652 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1436 decode.regfile.registers_21\[12\] VGND VGND VPWR VPWR net1663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 fetch.bht.bhtTable_tag\[6\]\[18\] VGND VGND VPWR VPWR net1674 sky130_fd_sc_hd__dlygate4sd3_1
X_23850_ _08087_ net1231 _08079_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1458 fetch.bht.bhtTable_tag\[11\]\[10\] VGND VGND VPWR VPWR net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1469 decode.regfile.registers_24\[7\] VGND VGND VPWR VPWR net1696 sky130_fd_sc_hd__dlygate4sd3_1
X_22801_ _07295_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_200_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23781_ _06143_ net2022 _08041_ VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20993_ execute.io_reg_pc\[21\] _05977_ _05973_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25520_ _08970_ _08978_ VGND VGND VPWR VPWR _09019_ sky130_fd_sc_hd__nand2_1
X_22732_ _07258_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25451_ _08978_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22663_ net2306 _07208_ _07217_ _07164_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_213_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24402_ _08378_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28170_ clknet_leaf_56_clock _01192_ VGND VGND VPWR VPWR csr.io_mret_vector\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_21614_ _06337_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25382_ _10035_ VGND VGND VPWR VPWR _08931_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22594_ csr._minstret_T_3\[46\] csr._minstret_T_3\[45\] _07170_ _06422_ VGND VGND
+ VPWR VPWR _07173_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27121_ clknet_leaf_351_clock _00150_ VGND VGND VPWR VPWR decode.regfile.registers_26\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24333_ _08095_ net1992 _08334_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21545_ _06292_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27052_ clknet_leaf_343_clock _00081_ VGND VGND VPWR VPWR decode.regfile.registers_23\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_24264_ _08307_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__clkbuf_1
X_21476_ _06105_ net2089 _06252_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26003_ net2192 _09286_ _09298_ _09292_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__o211a_1
X_23215_ _07347_ _07634_ _07649_ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__or3_1
X_20427_ _05582_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24195_ _08089_ net1330 _08266_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__mux2_1
X_23146_ execute.io_target_pc\[14\] _06037_ _10970_ _03592_ VGND VGND VPWR VPWR _07585_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_164_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20358_ _05519_ csr.io_csr_address\[11\] _05520_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__or3b_1
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27954_ clknet_leaf_199_clock _00976_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_23077_ execute.io_target_pc\[10\] _07346_ _07502_ _07519_ _07348_ VGND VGND VPWR
+ VPWR _07520_ sky130_fd_sc_hd__a2111o_1
X_20289_ _10681_ decode.id_ex_pc_reg\[16\] _05462_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__and3_1
X_22028_ _06622_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__buf_4
X_26905_ net2372 _09822_ _09830_ _09825_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__o211a_1
X_27885_ clknet_leaf_22_clock _00914_ VGND VGND VPWR VPWR csr._mcycle_T_2\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_944 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14850_ net336 _10891_ _10678_ VGND VGND VPWR VPWR _10893_ sky130_fd_sc_hd__o21a_1
X_29624_ clknet_leaf_270_clock _02637_ VGND VGND VPWR VPWR decode.regfile.registers_11\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26836_ net2552 _09779_ _09790_ _09784_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_67_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _10136_ _09937_ VGND VGND VPWR VPWR _10137_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1970 decode.regfile.registers_23\[31\] VGND VGND VPWR VPWR net2197 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ _10747_ _09887_ _09890_ VGND VGND VPWR VPWR _10824_ sky130_fd_sc_hd__nor3_1
Xhold1981 decode.regfile.registers_26\[30\] VGND VGND VPWR VPWR net2208 sky130_fd_sc_hd__dlygate4sd3_1
X_29555_ clknet_leaf_274_clock _02568_ VGND VGND VPWR VPWR decode.regfile.registers_9\[25\]
+ sky130_fd_sc_hd__dfxtp_2
X_26767_ _09750_ VGND VGND VPWR VPWR _09751_ sky130_fd_sc_hd__clkbuf_4
X_23979_ _08160_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__clkbuf_1
Xhold1992 fetch.bht.bhtTable_target_pc\[13\]\[30\] VGND VGND VPWR VPWR net2219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_63_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16520_ _12133_ net775 _12451_ _12485_ _11248_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__o221a_1
X_28506_ clknet_leaf_237_clock _01519_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13732_ _10003_ _10021_ memory.io_wb_readdata\[19\] VGND VGND VPWR VPWR _10078_ sky130_fd_sc_hd__and3b_1
X_25718_ _08941_ _09122_ VGND VGND VPWR VPWR _09134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26698_ net2500 _09709_ _09712_ _09702_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__o211a_1
X_29486_ clknet_leaf_264_clock _02499_ VGND VGND VPWR VPWR decode.regfile.registers_7\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16451_ decode.regfile.registers_14\[30\] _11207_ _11273_ decode.regfile.registers_15\[30\]
+ _11361_ VGND VGND VPWR VPWR _12418_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28437_ clknet_leaf_48_clock _01450_ VGND VGND VPWR VPWR decode.control.io_funct7\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_25649_ _08948_ _09092_ VGND VGND VPWR VPWR _09094_ sky130_fd_sc_hd__nand2_1
X_13663_ _10019_ VGND VGND VPWR VPWR _10020_ sky130_fd_sc_hd__clkbuf_4
X_15402_ decode.regfile.registers_27\[2\] _11237_ _11351_ _11395_ _11396_ VGND VGND
+ VPWR VPWR _11397_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19170_ _04303_ _04305_ _04463_ _04464_ _04465_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__o32a_1
XFILLER_0_112_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28368_ clknet_leaf_203_clock _01381_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16382_ decode.regfile.registers_3\[28\] _11110_ _11141_ _11145_ VGND VGND VPWR VPWR
+ _12351_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13594_ memory.io_wb_memtoreg\[1\] memory.io_wb_aluresult\[1\] memory.io_wb_memtoreg\[0\]
+ VGND VGND VPWR VPWR _09958_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18121_ _03488_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15333_ decode.regfile.registers_21\[1\] _11267_ _11099_ _11228_ _11328_ VGND VGND
+ VPWR VPWR _11329_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_97_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27319_ clknet_leaf_38_clock _00348_ VGND VGND VPWR VPWR decode.id_ex_ex_rs1_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_186_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28299_ clknet_leaf_164_clock _00013_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18052_ _10965_ _10998_ _10969_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15264_ _11235_ VGND VGND VPWR VPWR _11260_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_10_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17003_ _12496_ _12960_ _12961_ _12962_ VGND VGND VPWR VPWR _12963_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14215_ _09993_ _10377_ VGND VGND VPWR VPWR _10383_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_93_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15195_ _11178_ VGND VGND VPWR VPWR _11192_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14146_ _10015_ _10342_ VGND VGND VPWR VPWR _10343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14077_ _10290_ VGND VGND VPWR VPWR _10304_ sky130_fd_sc_hd__buf_2
X_18954_ _04233_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17905_ decode.regfile.registers_20\[28\] _11024_ _12553_ _12554_ _12537_ VGND VGND
+ VPWR VPWR _03304_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_52_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18885_ _04180_ net256 _04183_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__a21o_1
XFILLER_0_177_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17836_ _12497_ _12539_ _12503_ decode.regfile.registers_7\[26\] _12645_ VGND VGND
+ VPWR VPWR _03237_ sky130_fd_sc_hd__o32a_1
XFILLER_0_222_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer17 net242 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17767_ decode.regfile.registers_18\[24\] _10925_ _12569_ _11023_ _11009_ VGND VGND
+ VPWR VPWR _03170_ sky130_fd_sc_hd__o2111a_1
Xrebuffer28 net254 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_1
X_14979_ _10948_ _10954_ _10997_ net677 _10999_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__o311a_1
XFILLER_0_117_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer39 net263 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19506_ _04733_ _04790_ _04324_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__mux2_1
X_16718_ decode.regfile.registers_20\[0\] _12545_ _12563_ _12680_ _12682_ VGND VGND
+ VPWR VPWR _12683_ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17698_ _13407_ decode.regfile.registers_25\[22\] _13482_ _13294_ VGND VGND VPWR
+ VPWR _03103_ sky130_fd_sc_hd__or4_1
XFILLER_0_88_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19437_ _04495_ _04717_ _04718_ _04724_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__a31o_1
X_16649_ _12613_ VGND VGND VPWR VPWR _12614_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19368_ _04415_ _04644_ _04651_ _04658_ _03595_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__o311a_1
XFILLER_0_45_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18319_ decode.id_ex_rs2_data_reg\[25\] _03616_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__and2_1
X_19299_ _04591_ _04547_ _04247_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__mux2_1
Xrebuffer107 _04077_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_2
Xrebuffer118 _11150_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21330_ _06175_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21261_ _06133_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__clkbuf_1
Xhold500 decode.regfile.registers_13\[10\] VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 decode.regfile.registers_16\[17\] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 decode.regfile.registers_18\[15\] VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__dlygate4sd3_1
X_23000_ net94 net93 _07393_ net227 VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__a31o_1
Xhold533 fetch.bht.bhtTable_tag\[11\]\[3\] VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__dlygate4sd3_1
X_20212_ _05404_ _05405_ _05407_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21192_ _06091_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__clkbuf_1
Xhold544 decode.regfile.registers_8\[9\] VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 decode.regfile.registers_18\[6\] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold566 decode.regfile.registers_17\[19\] VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold577 decode.regfile.registers_5\[9\] VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold588 fetch.bht.bhtTable_tag\[4\]\[13\] VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlygate4sd3_1
X_20143_ _00568_ _05226_ _05349_ _05239_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold599 fetch.bht.bhtTable_target_pc\[3\]\[12\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20074_ _05288_ _05289_ _05282_ _05286_ _05283_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__o221ai_1
X_24951_ csr._mcycle_T_3\[52\] csr._mcycle_T_3\[51\] csr._mcycle_T_3\[50\] _08676_
+ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_202_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 fetch.bht.bhtTable_target_pc\[2\]\[26\] VGND VGND VPWR VPWR net1427 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_202_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1211 fetch.bht.bhtTable_target_pc\[6\]\[28\] VGND VGND VPWR VPWR net1438 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23902_ net827 _08060_ _08119_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__mux2_1
Xhold1222 decode.regfile.registers_18\[9\] VGND VGND VPWR VPWR net1449 sky130_fd_sc_hd__dlygate4sd3_1
X_27670_ clknet_leaf_27_clock _00699_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_24882_ csr.mcycle\[8\] csr.mcycle\[20\] _08629_ _08631_ VGND VGND VPWR VPWR _08632_
+ sky130_fd_sc_hd__and4_1
Xhold1233 fetch.bht.bhtTable_tag\[5\]\[5\] VGND VGND VPWR VPWR net1460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1244 decode.regfile.registers_25\[14\] VGND VGND VPWR VPWR net1471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1255 decode.regfile.registers_23\[30\] VGND VGND VPWR VPWR net1482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1266 fetch.bht.bhtTable_tag\[2\]\[24\] VGND VGND VPWR VPWR net1493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26621_ _09450_ _09666_ VGND VGND VPWR VPWR _09668_ sky130_fd_sc_hd__nand2_1
X_23833_ execute.io_target_pc\[13\] VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__buf_2
XFILLER_0_213_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1277 fetch.bht.bhtTable_tag\[0\]\[25\] VGND VGND VPWR VPWR net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1288 fetch.bht.bhtTable_tag\[6\]\[24\] VGND VGND VPWR VPWR net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 fetch.bht.bhtTable_tag\[14\]\[22\] VGND VGND VPWR VPWR net1526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29340_ clknet_leaf_246_clock _02353_ VGND VGND VPWR VPWR decode.regfile.registers_3\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26552_ _09381_ _09623_ VGND VGND VPWR VPWR _09628_ sky130_fd_sc_hd__nand2_1
X_23764_ _06126_ net1333 _08030_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20976_ _05970_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25503_ _08954_ _09005_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22715_ _06578_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__buf_4
X_29271_ clknet_leaf_224_clock _02284_ VGND VGND VPWR VPWR decode.regfile.registers_0\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_157_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26483_ _09387_ _09579_ VGND VGND VPWR VPWR _09588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23695_ net1235 _10812_ _07992_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28222_ clknet_leaf_87_clock net2143 VGND VGND VPWR VPWR csr.mscratch\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25434_ _08966_ _08946_ VGND VGND VPWR VPWR _08967_ sky130_fd_sc_hd__nand2_1
X_22646_ _06457_ net217 _06458_ _06466_ VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__and4_1
XFILLER_0_165_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28153_ clknet_leaf_188_clock _01175_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25365_ _08918_ _08907_ VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22577_ csr._minstret_T_3\[33\] csr._minstret_T_3\[32\] csr.minstret\[31\] _07152_
+ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27104_ clknet_leaf_357_clock _00133_ VGND VGND VPWR VPWR decode.regfile.registers_25\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24316_ _06186_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21528_ _06282_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__buf_6
X_28084_ clknet_leaf_213_clock _01106_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25296_ _08878_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27035_ clknet_leaf_345_clock _00064_ VGND VGND VPWR VPWR decode.regfile.registers_23\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_24247_ _08298_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__clkbuf_1
X_21459_ _06245_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14000_ _10031_ _10255_ VGND VGND VPWR VPWR _10259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_14__f_clock clknet_2_1_0_clock VGND VGND VPWR VPWR clknet_5_14__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_112_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24178_ _08072_ net930 _08255_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_187_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23129_ _07391_ _07392_ _07567_ _07568_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_183_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28986_ clknet_leaf_178_clock _01999_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput75 net75 VGND VGND VPWR VPWR io_fetch_address[17] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput86 net86 VGND VGND VPWR VPWR io_fetch_address[27] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 net97 VGND VGND VPWR VPWR io_fetch_address[8] sky130_fd_sc_hd__clkbuf_4
X_27937_ clknet_leaf_216_clock _00959_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_125_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15951_ decode.regfile.registers_18\[16\] _11455_ _11456_ _11931_ VGND VGND VPWR
+ VPWR _11932_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14902_ _10936_ VGND VGND VPWR VPWR _10937_ sky130_fd_sc_hd__clkbuf_4
X_15882_ _11079_ _11244_ _11261_ _11835_ _11864_ VGND VGND VPWR VPWR _11865_ sky130_fd_sc_hd__a41o_1
X_18670_ _03967_ _03654_ _03968_ _03649_ net353 VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__a41o_2
X_27868_ clknet_leaf_325_clock _00897_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2490 decode.regfile.registers_26\[28\] VGND VGND VPWR VPWR net2717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17621_ _02990_ _13176_ decode.regfile.registers_27\[20\] _13487_ VGND VGND VPWR
+ VPWR _03028_ sky130_fd_sc_hd__or4_1
X_29607_ clknet_leaf_275_clock _02620_ VGND VGND VPWR VPWR decode.regfile.registers_11\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14833_ _10871_ _10763_ _10872_ VGND VGND VPWR VPWR _10876_ sky130_fd_sc_hd__a21oi_1
X_26819_ net2329 _09779_ _09781_ _09771_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_4_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27799_ clknet_leaf_323_clock _00828_ VGND VGND VPWR VPWR memory.io_wb_readdata\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_142_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14764_ csr.io_mem_pc\[15\] VGND VGND VPWR VPWR _10807_ sky130_fd_sc_hd__buf_4
X_17552_ decode.regfile.registers_1\[19\] _12932_ _12830_ _12882_ _02959_ VGND VGND
+ VPWR VPWR _02960_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29538_ clknet_leaf_252_clock _02551_ VGND VGND VPWR VPWR decode.regfile.registers_9\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13715_ _10063_ VGND VGND VPWR VPWR _10064_ sky130_fd_sc_hd__buf_4
X_16503_ _11364_ decode.regfile.registers_11\[31\] _11690_ _12468_ VGND VGND VPWR
+ VPWR _12469_ sky130_fd_sc_hd__o211a_1
X_17483_ decode.regfile.registers_10\[17\] _10603_ _12503_ _12597_ VGND VGND VPWR
+ VPWR _13431_ sky130_fd_sc_hd__or4b_1
XFILLER_0_86_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14695_ _10674_ decode.id_ex_pc_reg\[1\] _10710_ _10709_ _10737_ VGND VGND VPWR VPWR
+ _10738_ sky130_fd_sc_hd__o221a_1
X_29469_ clknet_leaf_253_clock _02482_ VGND VGND VPWR VPWR decode.regfile.registers_7\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19222_ _04321_ _04021_ _04228_ _04449_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_15_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16434_ _11199_ _12400_ _12401_ _11203_ VGND VGND VPWR VPWR _12402_ sky130_fd_sc_hd__a211o_1
X_13646_ _09981_ VGND VGND VPWR VPWR _10004_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_15_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19153_ _04022_ _04448_ _04228_ _04449_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__and4b_1
X_16365_ decode.regfile.registers_19\[27\] _11406_ _11325_ _12334_ VGND VGND VPWR
+ VPWR _12335_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13577_ _09941_ VGND VGND VPWR VPWR _09942_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18104_ _03478_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__clkbuf_1
X_15316_ decode.regfile.registers_10\[1\] _10638_ _11132_ _11282_ _11311_ VGND VGND
+ VPWR VPWR _11312_ sky130_fd_sc_hd__o32a_1
XFILLER_0_147_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16296_ _10958_ decode.regfile.registers_26\[25\] _11676_ _11338_ _11564_ VGND VGND
+ VPWR VPWR _12268_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_48_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19084_ _04379_ _04381_ _04352_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15247_ _11065_ VGND VGND VPWR VPWR _11244_ sky130_fd_sc_hd__clkbuf_4
X_18035_ decode.regfile.registers_17\[31\] _12719_ _12826_ VGND VGND VPWR VPWR _03431_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15178_ _11174_ VGND VGND VPWR VPWR _11175_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14129_ _09950_ _10333_ VGND VGND VPWR VPWR _10334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19986_ _03588_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18937_ _04226_ _04227_ _04232_ _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__and4_1
XFILLER_0_158_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18868_ _03708_ decode.id_ex_imm_reg\[10\] _04161_ _04163_ _04166_ VGND VGND VPWR
+ VPWR _04167_ sky130_fd_sc_hd__a221o_2
XFILLER_0_207_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17819_ _02990_ _03068_ decode.regfile.registers_27\[25\] _13487_ VGND VGND VPWR
+ VPWR _03221_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18799_ execute.csr_read_data_out_reg\[13\] _03658_ _04097_ VGND VGND VPWR VPWR _04098_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_178_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20830_ _05866_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20761_ _05849_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22500_ _06041_ _07094_ _06481_ _07065_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23480_ _04459_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__buf_2
XFILLER_0_147_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20692_ _05801_ _05808_ decode.id_ex_rs1_data_reg\[7\] _05812_ _00694_ VGND VGND
+ VPWR VPWR _00726_ sky130_fd_sc_hd__a32o_1
XFILLER_0_169_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22431_ _06700_ fetch.bht.bhtTable_tag\[14\]\[12\] _06675_ _07025_ VGND VGND VPWR
+ VPWR _07026_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25150_ _10573_ net2584 _08802_ VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__mux2_1
X_22362_ fetch.bht.bhtTable_tag\[0\]\[2\] fetch.bht.bhtTable_tag\[1\]\[2\] fetch.bht.bhtTable_tag\[2\]\[2\]
+ fetch.bht.bhtTable_tag\[3\]\[2\] _06679_ _06620_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__mux4_2
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24101_ _08223_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__clkbuf_1
X_21313_ _06166_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25081_ _08704_ _03567_ _06566_ _08768_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22293_ net226 _06877_ _06886_ _06887_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24032_ net1712 execute.io_target_pc\[4\] _08187_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__mux2_1
X_21244_ _10868_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__buf_2
Xhold330 decode.regfile.registers_30\[27\] VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 decode.regfile.registers_23\[29\] VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _01117_ VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold363 csr._mcycle_T_2\[3\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__clkbuf_2
X_28840_ clknet_leaf_101_clock _01853_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold374 decode.regfile.registers_28\[1\] VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_68_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21175_ _09955_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__buf_2
Xhold385 decode.regfile.registers_13\[11\] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold396 decode.regfile.registers_15\[9\] VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20126_ decode.id_ex_imm_reg\[15\] _10681_ _05321_ _05324_ VGND VGND VPWR VPWR _05335_
+ sky130_fd_sc_hd__o211ai_1
X_28771_ clknet_leaf_132_clock _01784_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25983_ _09285_ VGND VGND VPWR VPWR _09287_ sky130_fd_sc_hd__buf_2
X_20057_ decode.id_ex_imm_reg\[8\] decode.id_ex_pc_reg\[8\] VGND VGND VPWR VPWR _05276_
+ sky130_fd_sc_hd__xnor2_1
X_24934_ net2616 _08668_ _08669_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__o21a_1
X_27722_ clknet_leaf_23_clock _00751_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1030 fetch.bht.bhtTable_target_pc\[11\]\[23\] VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 fetch.bht.bhtTable_tag\[4\]\[21\] VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 fetch.bht.bhtTable_tag\[9\]\[7\] VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 fetch.bht.bhtTable_target_pc\[5\]\[24\] VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__dlygate4sd3_1
X_24865_ _08620_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_159_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27653_ clknet_leaf_48_clock _00682_ VGND VGND VPWR VPWR execute.io_reg_pc\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1074 decode.regfile.registers_23\[3\] VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 fetch.bht.bhtTable_target_pc\[5\]\[26\] VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1096 fetch.bht.bhtTable_target_pc\[12\]\[6\] VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__dlygate4sd3_1
X_23816_ _08064_ net1906 _08058_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26604_ _09434_ _09645_ VGND VGND VPWR VPWR _09657_ sky130_fd_sc_hd__nand2_1
X_27584_ clknet_leaf_136_clock _00613_ VGND VGND VPWR VPWR csr.io_mem_pc\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24796_ _08584_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29323_ clknet_leaf_226_clock _02336_ VGND VGND VPWR VPWR decode.regfile.registers_2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_26535_ _09441_ _09577_ VGND VGND VPWR VPWR _09617_ sky130_fd_sc_hd__nand2_1
X_23747_ _06109_ net1680 _09907_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20959_ _03582_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_81_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13500_ csr.io_mem_pc\[5\] VGND VGND VPWR VPWR _09882_ sky130_fd_sc_hd__clkbuf_4
X_29254_ clknet_leaf_233_clock _02267_ VGND VGND VPWR VPWR decode.regfile.registers_0\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14480_ _10092_ _10530_ VGND VGND VPWR VPWR _10536_ sky130_fd_sc_hd__nand2_1
X_26466_ _09577_ VGND VGND VPWR VPWR _09578_ sky130_fd_sc_hd__clkbuf_4
X_23678_ net1493 _10777_ _07983_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28205_ clknet_leaf_63_clock net2020 VGND VGND VPWR VPWR csr.mscratch\[7\] sky130_fd_sc_hd__dfxtp_1
X_25417_ net818 _08951_ _08955_ _08950_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__o211a_1
X_22629_ _06377_ _07194_ _07196_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__nor3_1
X_29185_ clknet_leaf_162_clock _02198_ VGND VGND VPWR VPWR fetch.btb.btbTable\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26397_ net555 _09534_ _09538_ _09525_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28136_ clknet_leaf_206_clock _01158_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16150_ decode.regfile.registers_23\[21\] _11088_ _12100_ _12125_ VGND VGND VPWR
+ VPWR _12126_ sky130_fd_sc_hd__o22a_1
XFILLER_0_183_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25348_ _09950_ _08907_ VGND VGND VPWR VPWR _08908_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_114_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer8 _03744_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
X_15101_ _11097_ VGND VGND VPWR VPWR _11098_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_224_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28067_ clknet_leaf_169_clock _01089_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_16081_ decode.regfile.registers_3\[20\] _11110_ _11142_ _11146_ VGND VGND VPWR VPWR
+ _12058_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25279_ _08869_ net2470 VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_185_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15032_ net451 _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__a31o_1
X_27018_ clknet_leaf_342_clock _00047_ VGND VGND VPWR VPWR decode.regfile.registers_22\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19840_ _05089_ _05110_ _05111_ _05041_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19771_ _03852_ _03839_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__nand2_2
XFILLER_0_208_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28969_ clknet_leaf_96_clock _01982_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16983_ _12611_ _12941_ _12942_ VGND VGND VPWR VPWR _12943_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_88_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18722_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_144_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15934_ decode.regfile.registers_1\[16\] _11116_ _11137_ _11157_ VGND VGND VPWR VPWR
+ _11915_ sky130_fd_sc_hd__and4_1
XFILLER_0_218_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18653_ _03715_ _03725_ _03951_ _03727_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__o31a_1
X_15865_ _11845_ _11846_ _11847_ VGND VGND VPWR VPWR _11848_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_189_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17604_ decode.regfile.registers_10\[20\] _12652_ _12791_ VGND VGND VPWR VPWR _03011_
+ sky130_fd_sc_hd__o21a_1
X_14816_ _10779_ _10826_ _10697_ VGND VGND VPWR VPWR _10859_ sky130_fd_sc_hd__a21o_1
X_18584_ memory.csr_read_data_out_reg\[22\] _09987_ _10095_ VGND VGND VPWR VPWR _03883_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15796_ decode.regfile.registers_15\[12\] _11037_ _11205_ _11208_ decode.regfile.registers_14\[12\]
+ VGND VGND VPWR VPWR _11781_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_47_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17535_ _12505_ VGND VGND VPWR VPWR _13482_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_47_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14747_ decode.id_ex_pc_reg\[25\] VGND VGND VPWR VPWR _10790_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_103_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14678_ decode.id_ex_pc_reg\[10\] VGND VGND VPWR VPWR _10721_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17466_ net399 _12709_ _13377_ _13414_ _13219_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19205_ _04499_ _04454_ _04500_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16417_ decode.regfile.registers_9\[29\] _11365_ decode.regfile.registers_8\[29\]
+ _11285_ _11382_ VGND VGND VPWR VPWR _12385_ sky130_fd_sc_hd__o221ai_1
X_13629_ _09988_ VGND VGND VPWR VPWR _09989_ sky130_fd_sc_hd__buf_6
X_17397_ _13343_ _13345_ _13346_ VGND VGND VPWR VPWR _13347_ sky130_fd_sc_hd__o21a_2
XFILLER_0_171_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19136_ _04431_ _04432_ net242 VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__mux2_1
X_16348_ decode.regfile.registers_2\[27\] _11190_ _11148_ _11151_ _12317_ VGND VGND
+ VPWR VPWR _12318_ sky130_fd_sc_hd__o311a_1
XFILLER_0_27_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19067_ _04363_ _04364_ _04277_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__mux2_1
X_16279_ decode.regfile.registers_8\[25\] _11165_ _11547_ decode.regfile.registers_9\[25\]
+ _11182_ VGND VGND VPWR VPWR _12251_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18018_ decode.regfile.registers_1\[31\] _12778_ _12634_ _03413_ VGND VGND VPWR VPWR
+ _03414_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_23_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19969_ _05215_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22980_ net93 net92 net89 net94 VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_220_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21931_ csr._mcycle_T_2\[28\] _06545_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24650_ _07284_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21862_ csr.io_mret_vector\[8\] _10881_ _06040_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__mux2_1
X_23601_ _07946_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20813_ net125 _05879_ _05875_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__and3_1
X_24581_ _08472_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__clkbuf_1
X_21793_ _06462_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26320_ net583 _09491_ _09494_ _09484_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23532_ net2184 _07904_ _07901_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20744_ _05818_ decode.id_ex_rs1_data_reg\[29\] _05780_ VGND VGND VPWR VPWR _05843_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26251_ net657 _09447_ _09454_ _09440_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_189_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23463_ net10 _07861_ _07868_ _07865_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_189_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20675_ _05792_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_169_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25202_ _09880_ _09883_ _10569_ VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22414_ fetch.bht.bhtTable_tag\[4\]\[1\] fetch.bht.bhtTable_tag\[5\]\[1\] fetch.bht.bhtTable_tag\[6\]\[1\]
+ fetch.bht.bhtTable_tag\[7\]\[1\] _06680_ _06684_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__mux4_1
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26182_ _09406_ _09390_ VGND VGND VPWR VPWR _09407_ sky130_fd_sc_hd__nand2_1
X_23394_ _07619_ _07345_ _07620_ _07817_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__a31o_1
XFILLER_0_162_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25133_ _06151_ net1872 _08562_ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__mux2_1
X_22345_ fetch.bht.bhtTable_tag\[14\]\[10\] fetch.bht.bhtTable_tag\[15\]\[10\] _06809_
+ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_76_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_227_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25064_ _03555_ csr.mcycle\[21\] _08745_ VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__and3_1
X_29941_ clknet_leaf_340_clock _02954_ VGND VGND VPWR VPWR decode.regfile.registers_21\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_22276_ fetch.bht.bhtTable_tag\[0\]\[6\] fetch.bht.bhtTable_tag\[1\]\[6\] fetch.bht.bhtTable_tag\[2\]\[6\]
+ fetch.bht.bhtTable_tag\[3\]\[6\] _06645_ _06651_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_148_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24015_ net925 execute.io_target_pc\[28\] _07960_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21227_ _06110_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__clkbuf_1
Xhold160 io_fetch_data[2] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold171 fetch.bht.bhtTable_valid\[1\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29872_ clknet_leaf_300_clock _02885_ VGND VGND VPWR VPWR decode.regfile.registers_19\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_180_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold182 decode.regfile.registers_31\[13\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_218_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold193 fetch.btb.btbTable\[14\]\[0\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28823_ clknet_leaf_133_clock _01836_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21158_ _06062_ _06070_ execute.csr_write_data_out_reg\[23\] VGND VGND VPWR VPWR
+ _06073_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_70_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20109_ decode.id_ex_imm_reg\[16\] decode.id_ex_pc_reg\[16\] VGND VGND VPWR VPWR
+ _05320_ sky130_fd_sc_hd__nand2_1
X_28754_ clknet_leaf_106_clock _01767_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_13980_ net2401 _10243_ _10247_ _10232_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__o211a_1
X_21089_ _10971_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__buf_4
X_25966_ _09263_ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27705_ clknet_leaf_20_clock _00734_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_24917_ csr._mcycle_T_3\[40\] csr._mcycle_T_3\[39\] csr._mcycle_T_3\[38\] _08654_
+ VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_107_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28685_ clknet_leaf_108_clock _01698_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_107_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25897_ net2740 _09226_ _09236_ _09235_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27636_ clknet_leaf_155_clock _00665_ VGND VGND VPWR VPWR execute.io_reg_pc\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_15650_ decode.regfile.registers_23\[8\] _11088_ _11612_ _11638_ VGND VGND VPWR VPWR
+ _11639_ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24848_ _06126_ net1875 _08607_ VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_178_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_50 _09983_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_61 _10121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_72 _10198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_83 _10588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14601_ _10626_ _10634_ _10641_ _10643_ VGND VGND VPWR VPWR _10644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_94 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15581_ _10961_ VGND VGND VPWR VPWR _11571_ sky130_fd_sc_hd__clkbuf_4
X_24779_ _08072_ net1468 _08574_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27567_ clknet_leaf_157_clock _00596_ VGND VGND VPWR VPWR csr.io_mem_pc\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14532_ net66 VGND VGND VPWR VPWR _10575_ sky130_fd_sc_hd__buf_4
X_29306_ clknet_leaf_243_clock _02319_ VGND VGND VPWR VPWR decode.regfile.registers_2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_17320_ decode.regfile.registers_4\[13\] _12549_ _12532_ decode.regfile.registers_5\[13\]
+ _12626_ VGND VGND VPWR VPWR _13272_ sky130_fd_sc_hd__a221o_1
X_26518_ net2274 _09605_ _09607_ _09608_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27498_ clknet_leaf_29_clock _00527_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29237_ clknet_leaf_180_clock _02250_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17251_ decode.regfile.registers_19\[11\] _12678_ _13185_ _13204_ _12906_ VGND VGND
+ VPWR VPWR _13205_ sky130_fd_sc_hd__o221a_1
X_14463_ _10053_ _10517_ VGND VGND VPWR VPWR _10526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26449_ net2758 _09561_ _09568_ _09567_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16202_ decode.regfile.registers_1\[23\] _11117_ _11057_ _11109_ VGND VGND VPWR VPWR
+ _12176_ sky130_fd_sc_hd__and4_1
XFILLER_0_126_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17182_ net441 _12709_ _13098_ _13137_ _12705_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__o221a_1
XFILLER_0_226_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29168_ clknet_leaf_168_clock _02181_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14394_ _10069_ _10474_ VGND VGND VPWR VPWR _10486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16133_ decode.regfile.registers_5\[21\] _11291_ _12107_ _12108_ VGND VGND VPWR VPWR
+ _12109_ sky130_fd_sc_hd__a22oi_2
X_28119_ clknet_leaf_90_clock _01141_ VGND VGND VPWR VPWR csr.minstret\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29099_ clknet_leaf_71_clock _02112_ VGND VGND VPWR VPWR csr._mcycle_T_3\[47\] sky130_fd_sc_hd__dfxtp_1
X_16064_ decode.regfile.registers_19\[19\] _11048_ _11215_ _11216_ _11325_ VGND VGND
+ VPWR VPWR _12042_ sky130_fd_sc_hd__o41a_1
XFILLER_0_80_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15015_ _11024_ VGND VGND VPWR VPWR _11025_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19823_ _04921_ _04371_ _04392_ _05094_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_36_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19754_ _05019_ _05020_ _05028_ _04667_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__o211a_1
X_16966_ decode.regfile.registers_15\[5\] _12555_ _10923_ _12876_ _12672_ VGND VGND
+ VPWR VPWR _12926_ sky130_fd_sc_hd__a41o_1
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18705_ _03816_ _04000_ _04001_ _03998_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15917_ _11225_ _11125_ _11216_ decode.regfile.registers_17\[15\] _11128_ VGND VGND
+ VPWR VPWR _11899_ sky130_fd_sc_hd__o32a_1
X_19685_ _04589_ _04954_ _04961_ _04962_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__a22o_1
XFILLER_0_216_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16897_ decode.regfile.registers_21\[3\] _12822_ _12825_ _12858_ _12806_ VGND VGND
+ VPWR VPWR _12859_ sky130_fd_sc_hd__o221a_1
XFILLER_0_194_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18636_ _03890_ decode.id_ex_imm_reg\[17\] _03906_ _03907_ VGND VGND VPWR VPWR _03935_
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_189_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15848_ _11646_ _11253_ _11064_ decode.regfile.registers_29\[13\] _11831_ VGND VGND
+ VPWR VPWR _11832_ sky130_fd_sc_hd__o221a_1
XFILLER_0_91_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18567_ _03853_ _03854_ _03865_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15779_ _11435_ decode.regfile.registers_22\[12\] _11450_ _10979_ _10991_ VGND VGND
+ VPWR VPWR _11764_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_364_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_364_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17518_ _12790_ _13464_ VGND VGND VPWR VPWR _13465_ sky130_fd_sc_hd__nand2_1
X_18498_ net308 VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17449_ decode.regfile.registers_15\[16\] _12666_ _12773_ _12575_ _13397_ VGND VGND
+ VPWR VPWR _13398_ sky130_fd_sc_hd__o311a_1
XFILLER_0_89_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20460_ _05595_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19119_ net190 _04254_ _04265_ _04352_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__o211a_1
X_20391_ net294 _05534_ _05525_ _05536_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22130_ fetch.bht.bhtTable_tag\[14\]\[4\] fetch.bht.bhtTable_tag\[15\]\[4\] _06680_
+ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_302_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_302_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22061_ _06630_ _06638_ _06655_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_227_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21012_ _05990_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_222_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25820_ _08968_ _09155_ VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_317_clock clknet_5_18__leaf_clock VGND VGND VPWR VPWR clknet_leaf_317_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_215_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25751_ _08975_ _09110_ VGND VGND VPWR VPWR _09152_ sky130_fd_sc_hd__nand2_1
X_22963_ net92 net89 net93 VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24702_ _08064_ net1865 _08531_ VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__mux2_1
X_21914_ _06549_ _06543_ _06544_ _06550_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__o211a_1
X_28470_ clknet_leaf_138_clock _01483_ VGND VGND VPWR VPWR decode.io_id_pc\[28\] sky130_fd_sc_hd__dfxtp_1
X_25682_ net1134 _09111_ _09113_ _09100_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__o211a_1
X_22894_ _03592_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24633_ _08499_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__clkbuf_1
X_27421_ clknet_leaf_29_clock _00450_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[30\]
+ sky130_fd_sc_hd__dfxtp_2
X_21845_ net2581 _06497_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_216_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24564_ net1226 execute.io_target_pc\[4\] _08462_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27352_ clknet_leaf_46_clock _00381_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[25\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_216_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21776_ _06451_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_173_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23515_ net2255 _07889_ _07898_ _07893_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26303_ _09417_ VGND VGND VPWR VPWR _09484_ sky130_fd_sc_hd__buf_4
XFILLER_0_93_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27283_ clknet_leaf_32_clock _00312_ VGND VGND VPWR VPWR decode.regfile.registers_31\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20727_ _05831_ _05808_ decode.id_ex_rs1_data_reg\[21\] _05833_ _00708_ VGND VGND
+ VPWR VPWR _00740_ sky130_fd_sc_hd__a32o_1
X_24495_ _09901_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_1098 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29022_ clknet_leaf_135_clock _02035_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26234_ _10146_ VGND VGND VPWR VPWR _09443_ sky130_fd_sc_hd__clkbuf_4
X_23446_ _10941_ _07847_ _05206_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__or3b_1
X_20658_ _05585_ _05552_ csr.mcycle\[31\] VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26165_ _09372_ VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__clkbuf_4
X_23377_ _06038_ csr.io_mret_vector\[28\] _06041_ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__or3b_1
XFILLER_0_34_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20589_ net2006 _05593_ _05625_ _05727_ _05728_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__o32a_1
XFILLER_0_162_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25116_ _08786_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22328_ fetch.bht.bhtTable_tag\[4\]\[8\] fetch.bht.bhtTable_tag\[5\]\[8\] fetch.bht.bhtTable_tag\[6\]\[8\]
+ fetch.bht.bhtTable_tag\[7\]\[8\] _06878_ _06677_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__mux4_1
X_26096_ net2357 _09343_ _09351_ _09346_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25047_ net342 _03562_ _03554_ csr.mcycle\[20\] VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__and4_1
X_29924_ clknet_leaf_337_clock _02937_ VGND VGND VPWR VPWR decode.regfile.registers_21\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_22259_ _06853_ _06650_ _06686_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_167_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29855_ clknet_leaf_306_clock _02868_ VGND VGND VPWR VPWR decode.regfile.registers_19\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28806_ clknet_leaf_94_clock _01819_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16820_ _12780_ _12781_ _12782_ VGND VGND VPWR VPWR _12783_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_219_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29786_ clknet_leaf_309_clock _02799_ VGND VGND VPWR VPWR decode.regfile.registers_17\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_26998_ clknet_leaf_334_clock _00027_ VGND VGND VPWR VPWR decode.regfile.registers_22\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28737_ clknet_leaf_174_clock _01750_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16751_ _10926_ decode.regfile.registers_22\[1\] _12554_ _11009_ _12546_ VGND VGND
+ VPWR VPWR _12715_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_219_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13963_ _10128_ _10198_ VGND VGND VPWR VPWR _10236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25949_ _09241_ VGND VGND VPWR VPWR _09267_ sky130_fd_sc_hd__buf_2
XFILLER_0_216_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15702_ _11191_ _10630_ _11051_ VGND VGND VPWR VPWR _11689_ sky130_fd_sc_hd__or3_2
X_19470_ net316 VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__inv_2
X_28668_ clknet_leaf_176_clock _01681_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_13894_ _10194_ VGND VGND VPWR VPWR _10195_ sky130_fd_sc_hd__clkbuf_4
X_16682_ _12612_ _12643_ _12646_ VGND VGND VPWR VPWR _12647_ sky130_fd_sc_hd__o21a_1
XFILLER_0_186_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18421_ _03642_ _03718_ execute.io_mem_rd\[3\] _03719_ VGND VGND VPWR VPWR _03720_
+ sky130_fd_sc_hd__a22oi_2
X_27619_ clknet_leaf_153_clock _00648_ VGND VGND VPWR VPWR execute.io_target_pc\[28\]
+ sky130_fd_sc_hd__dfxtp_4
X_15633_ decode.regfile.registers_7\[8\] _11092_ _11167_ _11170_ decode.regfile.registers_6\[8\]
+ VGND VGND VPWR VPWR _11622_ sky130_fd_sc_hd__a32o_1
XFILLER_0_186_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_304 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28599_ clknet_leaf_124_clock _01612_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_315 decode.regfile.registers_11\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_326 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_337 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18352_ _09920_ decode.id_ex_ex_rs1_reg\[4\] VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_348 _03580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15564_ _11554_ decode.regfile.registers_17\[6\] _11356_ VGND VGND VPWR VPWR _11555_
+ sky130_fd_sc_hd__mux2_1
XINSDIODE1_359 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17303_ _13183_ _13252_ _13253_ _13255_ VGND VGND VPWR VPWR _13256_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_29_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ fetch.btb.btbTable\[12\]\[0\] fetch.btb.btbTable\[13\]\[0\] fetch.btb.btbTable\[14\]\[0\]
+ fetch.btb.btbTable\[15\]\[0\] _10556_ _10557_ VGND VGND VPWR VPWR _10560_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15495_ _11251_ _11259_ decode.regfile.registers_27\[4\] _11449_ _11487_ VGND VGND
+ VPWR VPWR _11488_ sky130_fd_sc_hd__o32a_1
X_18283_ _03606_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17234_ decode.regfile.registers_13\[11\] _12927_ _12583_ VGND VGND VPWR VPWR _13188_
+ sky130_fd_sc_hd__and3_1
X_14446_ _10008_ _10507_ VGND VGND VPWR VPWR _10516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17165_ _11023_ _12569_ _12535_ _13120_ VGND VGND VPWR VPWR _13121_ sky130_fd_sc_hd__a31o_1
X_14377_ net458 _10463_ _10476_ _10468_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold907 decode.regfile.registers_5\[0\] VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 fetch.bht.bhtTable_tag\[9\]\[25\] VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16116_ _11396_ _12090_ _12091_ _12092_ VGND VGND VPWR VPWR _12093_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold929 fetch.bht.bhtTable_target_pc\[1\]\[11\] VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__dlygate4sd3_1
X_17096_ _12765_ _12768_ _12493_ decode.regfile.registers_29\[7\] _13053_ VGND VGND
+ VPWR VPWR _13054_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_38_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16047_ decode.regfile.registers_2\[19\] _10646_ _11298_ _11151_ _12024_ VGND VGND
+ VPWR VPWR _12025_ sky130_fd_sc_hd__o311a_1
XFILLER_0_228_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2308 csr.minstret\[21\] VGND VGND VPWR VPWR net2535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2319 decode.regfile.registers_26\[22\] VGND VGND VPWR VPWR net2546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19806_ _03852_ _05048_ _05049_ _03814_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__a31o_1
Xhold1607 csr.mscratch\[15\] VGND VGND VPWR VPWR net1834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1618 fetch.bht.bhtTable_tag\[13\]\[15\] VGND VGND VPWR VPWR net1845 sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ decode.regfile.registers_15\[30\] _12874_ _03379_ _03394_ _12576_ VGND VGND
+ VPWR VPWR _03395_ sky130_fd_sc_hd__o221a_1
Xhold1629 decode.regfile.registers_1\[2\] VGND VGND VPWR VPWR net1856 sky130_fd_sc_hd__dlygate4sd3_1
X_19737_ _04805_ _04806_ _05012_ _04628_ _04729_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__o221ai_4
X_16949_ decode.regfile.registers_21\[4\] _12682_ _12909_ VGND VGND VPWR VPWR _12910_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_205_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19668_ _04281_ _04283_ _04945_ _04946_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__o31a_1
XFILLER_0_56_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18619_ decode.id_ex_rs1_data_reg\[18\] _03908_ _03913_ _03914_ _03917_ VGND VGND
+ VPWR VPWR _03918_ sky130_fd_sc_hd__o221a_4
XFILLER_0_172_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19599_ _04674_ _04546_ _04428_ _04880_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21630_ _05613_ csr.minstret\[5\] _06338_ _06349_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21561_ _06132_ net1845 _06295_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23300_ _07728_ _07729_ _07063_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__and3b_1
X_20512_ csr.mscratch\[10\] _05591_ _05611_ _05660_ _05661_ VGND VGND VPWR VPWR _05662_
+ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_211_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24280_ _08315_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21492_ _06251_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__buf_4
XFILLER_0_105_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23231_ fetch.bht.bhtTable_target_pc\[2\]\[19\] fetch.bht.bhtTable_target_pc\[3\]\[19\]
+ _07067_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__mux2_1
X_20443_ csr.minstret\[3\] _05594_ _05599_ csr.ie _05552_ VGND VGND VPWR VPWR _05600_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_241_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_241_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23162_ _05246_ _07591_ _07597_ _07599_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__o31a_1
X_20374_ net296 _05534_ _05525_ _05536_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_113_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22113_ fetch.bht.bhtTable_tag\[4\]\[3\] fetch.bht.bhtTable_tag\[5\]\[3\] _06707_
+ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27970_ clknet_leaf_212_clock _00992_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_23093_ _09956_ VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22044_ fetch.bht.bhtTable_tag\[0\]\[22\] fetch.bht.bhtTable_tag\[1\]\[22\] fetch.bht.bhtTable_tag\[2\]\[22\]
+ fetch.bht.bhtTable_tag\[3\]\[22\] _06619_ _06624_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__mux4_1
X_26921_ _10245_ _09840_ VGND VGND VPWR VPWR _09841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_256_clock clknet_5_19__leaf_clock VGND VGND VPWR VPWR clknet_leaf_256_clock
+ sky130_fd_sc_hd__clkbuf_8
X_29640_ clknet_leaf_278_clock _02653_ VGND VGND VPWR VPWR decode.regfile.registers_12\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_26852_ _09379_ _09796_ VGND VGND VPWR VPWR _09801_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_162_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25803_ _09155_ VGND VGND VPWR VPWR _09183_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29571_ clknet_leaf_252_clock _02584_ VGND VGND VPWR VPWR decode.regfile.registers_10\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_104_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23995_ net1276 execute.io_target_pc\[18\] _08164_ VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26783_ _09385_ _09753_ VGND VGND VPWR VPWR _09761_ sky130_fd_sc_hd__nand2_1
X_28522_ clknet_leaf_188_clock _01535_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22946_ _07390_ _07367_ _07090_ _07395_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__a211o_1
X_25734_ net2432 _09139_ _09143_ _09142_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_218_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28453_ clknet_leaf_147_clock _01466_ VGND VGND VPWR VPWR decode.io_id_pc\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22877_ _09896_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25665_ _08964_ _09092_ VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27404_ clknet_leaf_28_clock _00433_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_24616_ _08490_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21828_ _06480_ csr._csr_read_data_T_9\[2\] _06488_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28384_ clknet_leaf_145_clock _01397_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_4
X_25596_ _08970_ _09023_ VGND VGND VPWR VPWR _09063_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24547_ _08107_ net1799 _09902_ VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__mux2_1
X_27335_ clknet_leaf_46_clock _00364_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21759_ _06442_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14300_ net2228 _10419_ _10432_ _10427_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__o211a_1
X_15280_ _11275_ VGND VGND VPWR VPWR _11276_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24478_ _08105_ net1293 _08411_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27266_ clknet_leaf_0_clock _00295_ VGND VGND VPWR VPWR decode.regfile.registers_30\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29005_ clknet_leaf_103_clock _02018_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_14231_ net694 _10390_ _10392_ _10385_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23429_ _06422_ _10910_ _03500_ net26 VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_24_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26217_ decode.regfile.registers_11\[25\] _09419_ _09431_ _09418_ VGND VGND VPWR
+ VPWR _02632_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27197_ clknet_leaf_3_clock _00226_ VGND VGND VPWR VPWR decode.regfile.registers_28\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_209_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_209_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_130_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire178 _00664_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14162_ _10058_ _10342_ VGND VGND VPWR VPWR _10352_ sky130_fd_sc_hd__nand2_1
X_26148_ _09992_ VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_95_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18970_ _04268_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__clkbuf_4
X_14093_ _10286_ VGND VGND VPWR VPWR _10312_ sky130_fd_sc_hd__clkbuf_4
X_26079_ _08925_ _09340_ VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _12512_ _12772_ _12794_ _03318_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__o221a_1
X_29907_ clknet_leaf_340_clock _02920_ VGND VGND VPWR VPWR decode.regfile.registers_20\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17852_ _11014_ _10936_ decode.regfile.registers_23\[26\] _12995_ VGND VGND VPWR
+ VPWR _03253_ sky130_fd_sc_hd__or4_1
X_29838_ clknet_leaf_300_clock _02851_ VGND VGND VPWR VPWR decode.regfile.registers_18\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16803_ _10939_ _10606_ _10937_ _10933_ VGND VGND VPWR VPWR _12766_ sky130_fd_sc_hd__or4_1
XFILLER_0_227_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29769_ clknet_leaf_293_clock _02782_ VGND VGND VPWR VPWR decode.regfile.registers_16\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17783_ _13451_ net610 _13492_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__o21a_1
X_14995_ _10612_ VGND VGND VPWR VPWR _11008_ sky130_fd_sc_hd__buf_2
X_19522_ _04359_ _04306_ _03704_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_50_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16734_ _12693_ _12696_ _12698_ VGND VGND VPWR VPWR _12699_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_50_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13946_ _10087_ _10223_ VGND VGND VPWR VPWR _10227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19453_ _04155_ _04168_ _04738_ _04739_ _04154_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__a32o_1
XFILLER_0_158_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16665_ _12556_ _10601_ _10591_ _10614_ VGND VGND VPWR VPWR _12630_ sky130_fd_sc_hd__nand4_4
X_13877_ net2607 _10180_ _10185_ _10175_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_101 _10668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_112 _10994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18404_ _03656_ _03668_ _03670_ _03702_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__o211a_4
X_15616_ _11250_ decode.regfile.registers_27\[7\] _11258_ VGND VGND VPWR VPWR _11606_
+ sky130_fd_sc_hd__or3_1
XINSDIODE1_123 _11097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19384_ _04673_ _04554_ _04269_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__mux2_1
XINSDIODE1_134 _11347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16596_ _12560_ VGND VGND VPWR VPWR _12561_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_145 _12512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_156 _12690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18335_ decode.id_ex_aluop_reg\[2\] VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__clkbuf_4
XINSDIODE1_167 decode.id_ex_rs1_data_reg\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15547_ _11115_ _11055_ _11107_ VGND VGND VPWR VPWR _11538_ sky130_fd_sc_hd__and3_1
XINSDIODE1_178 execute.csr_read_data_out_reg\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_189 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18266_ decode.id_ex_rs2_data_reg\[0\] _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15478_ decode.regfile.registers_11\[4\] _11070_ _11470_ _11186_ VGND VGND VPWR VPWR
+ _11471_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17217_ _12516_ _13167_ _13169_ _13171_ VGND VGND VPWR VPWR _13172_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14429_ _10505_ VGND VGND VPWR VPWR _10506_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18197_ decode.control.io_funct7\[6\] decode.control.io_funct7\[4\] decode.control.io_funct7\[3\]
+ _03529_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__nor4_1
X_17148_ decode.regfile.registers_1\[9\] _12932_ _12933_ _10615_ _13103_ VGND VGND
+ VPWR VPWR _13104_ sky130_fd_sc_hd__o221a_1
Xhold704 decode.regfile.registers_28\[5\] VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold715 fetch.bht.bhtTable_target_pc\[8\]\[24\] VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold726 decode.id_ex_regwrite_reg VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold737 fetch.bht.bhtTable_tag\[11\]\[5\] VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold748 fetch.bht.bhtTable_tag\[1\]\[23\] VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 fetch.bht.bhtTable_target_pc\[2\]\[4\] VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17079_ decode.regfile.registers_20\[7\] _12545_ _13010_ _13036_ VGND VGND VPWR VPWR
+ _13037_ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20090_ _05283_ _05292_ _05298_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2105 decode.regfile.registers_5\[7\] VGND VGND VPWR VPWR net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2116 decode.regfile.registers_15\[26\] VGND VGND VPWR VPWR net2343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2127 csr._mcycle_T_3\[55\] VGND VGND VPWR VPWR net2354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2138 csr._mcycle_T_3\[59\] VGND VGND VPWR VPWR net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1404 fetch.bht.bhtTable_target_pc\[9\]\[23\] VGND VGND VPWR VPWR net1631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2149 decode.regfile.registers_12\[21\] VGND VGND VPWR VPWR net2376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1415 decode.regfile.registers_18\[30\] VGND VGND VPWR VPWR net1642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_204_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1426 fetch.bht.bhtTable_target_pc\[6\]\[14\] VGND VGND VPWR VPWR net1653 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1437 fetch.bht.bhtTable_tag\[15\]\[3\] VGND VGND VPWR VPWR net1664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1448 fetch.bht.bhtTable_tag\[5\]\[8\] VGND VGND VPWR VPWR net1675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 fetch.bht.bhtTable_target_pc\[10\]\[1\] VGND VGND VPWR VPWR net1686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22800_ net1071 _10872_ _07286_ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23780_ _08042_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_200_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20992_ _05979_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_200_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22731_ _06105_ net1962 _09903_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25450_ _08977_ VGND VGND VPWR VPWR _08978_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_220_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22662_ net1733 _07210_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_213_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24401_ net1442 execute.io_target_pc\[23\] _09911_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21613_ _06317_ _06333_ csr.io_inst_retired VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__and3_1
X_25381_ net2567 _08928_ _08930_ _08927_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__o211a_1
X_22593_ csr._minstret_T_3\[45\] csr._minstret_T_3\[44\] csr._minstret_T_3\[43\] _07166_
+ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__and4_1
XFILLER_0_34_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24332_ _08342_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27120_ clknet_leaf_351_clock _00149_ VGND VGND VPWR VPWR decode.regfile.registers_26\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21544_ _06115_ net2001 _06284_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_180_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_180_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27051_ clknet_leaf_338_clock _00080_ VGND VGND VPWR VPWR decode.regfile.registers_23\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24263_ _08091_ net1564 _08300_ VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21475_ _06254_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26002_ _08922_ _09297_ VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__nand2_1
X_23214_ execute.io_target_pc\[18\] _03592_ _03590_ _07648_ VGND VGND VPWR VPWR _07649_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20426_ _05576_ _05579_ _05584_ _05414_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__o31a_1
X_24194_ _08271_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23145_ _07391_ _07392_ _07582_ _07583_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_113_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20357_ csr.io_csr_address\[10\] csr.io_csr_address\[9\] csr.io_csr_address\[8\]
+ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__and3b_2
XFILLER_0_101_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_195_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_195_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_164_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27953_ clknet_leaf_202_clock _00975_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_23076_ _05246_ _07505_ _07518_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__nor3_1
XFILLER_0_140_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20288_ _10681_ _05462_ decode.id_ex_pc_reg\[16\] VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22027_ _06621_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__buf_4
X_26904_ _09432_ _09819_ VGND VGND VPWR VPWR _09830_ sky130_fd_sc_hd__nand2_1
X_27884_ clknet_leaf_23_clock _00913_ VGND VGND VPWR VPWR csr._mcycle_T_2\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29623_ clknet_leaf_277_clock _02636_ VGND VGND VPWR VPWR decode.regfile.registers_11\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_26835_ _09438_ _09751_ VGND VGND VPWR VPWR _09790_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1960 decode.regfile.registers_29\[1\] VGND VGND VPWR VPWR net2187 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _10135_ VGND VGND VPWR VPWR _10136_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_123_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29554_ clknet_leaf_274_clock _02567_ VGND VGND VPWR VPWR decode.regfile.registers_9\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1971 fetch.bht.bhtTable_tag\[10\]\[24\] VGND VGND VPWR VPWR net2198 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ net269 _10818_ decode.id_ex_pc_reg\[9\] VGND VGND VPWR VPWR _10823_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_123_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26766_ _10149_ _10150_ _03672_ VGND VGND VPWR VPWR _09750_ sky130_fd_sc_hd__and3_1
XFILLER_0_202_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23978_ net1775 execute.io_target_pc\[10\] _08153_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__mux2_1
Xhold1982 decode.regfile.registers_6\[12\] VGND VGND VPWR VPWR net2209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1993 decode.regfile.registers_19\[2\] VGND VGND VPWR VPWR net2220 sky130_fd_sc_hd__dlygate4sd3_1
X_28505_ clknet_leaf_239_clock _01518_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13731_ net2101 _10027_ _10076_ _10077_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__o211a_1
X_25717_ net616 _09125_ _09133_ _09129_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__o211a_1
X_22929_ _07130_ net89 VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__and2_1
X_29485_ clknet_leaf_264_clock _02498_ VGND VGND VPWR VPWR decode.regfile.registers_7\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26697_ _09450_ _09710_ VGND VGND VPWR VPWR _09712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_133_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_133_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28436_ clknet_leaf_48_clock _01449_ VGND VGND VPWR VPWR decode.control.io_funct7\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16450_ _11263_ decode.regfile.registers_22\[30\] _11404_ _11264_ _11265_ VGND VGND
+ VPWR VPWR _12417_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_39_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13662_ _10018_ VGND VGND VPWR VPWR _10019_ sky130_fd_sc_hd__buf_6
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25648_ net2550 _09082_ _09093_ _09087_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15401_ _11238_ VGND VGND VPWR VPWR _11396_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_26_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28367_ clknet_leaf_202_clock _01380_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13593_ net1891 _09938_ _09952_ _09957_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__o211a_1
X_16381_ decode.regfile.registers_5\[28\] _10636_ _11138_ _11169_ VGND VGND VPWR VPWR
+ _12350_ sky130_fd_sc_hd__a31o_1
X_25579_ _08954_ _09049_ VGND VGND VPWR VPWR _09054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18120_ _03482_ _03480_ _03487_ decode.io_id_pc\[16\] VGND VGND VPWR VPWR _03488_
+ sky130_fd_sc_hd__and4bb_1
X_15332_ decode.regfile.registers_20\[1\] _11102_ _11324_ _11326_ _11327_ VGND VGND
+ VPWR VPWR _11328_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27318_ clknet_leaf_38_clock _00347_ VGND VGND VPWR VPWR decode.id_ex_ex_rd_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_152_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28298_ clknet_leaf_164_clock _00014_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_148_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_148_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18051_ net775 _12872_ _03409_ _03446_ _03073_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__o221a_1
XFILLER_0_81_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15263_ _11258_ VGND VGND VPWR VPWR _11259_ sky130_fd_sc_hd__clkbuf_4
X_27249_ clknet_leaf_32_clock _00278_ VGND VGND VPWR VPWR decode.regfile.registers_30\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17002_ _12701_ decode.regfile.registers_28\[5\] _12698_ VGND VGND VPWR VPWR _12962_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_93_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14214_ net982 _10376_ _10382_ _10369_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__o211a_1
X_15194_ _11190_ VGND VGND VPWR VPWR _11191_ sky130_fd_sc_hd__buf_4
XANTENNA_6 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_227_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14145_ _10331_ VGND VGND VPWR VPWR _10342_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14076_ _10031_ _10299_ VGND VGND VPWR VPWR _10303_ sky130_fd_sc_hd__nand2_1
X_18953_ _03998_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17904_ _10926_ decode.regfile.registers_22\[28\] _12554_ _11009_ _12546_ VGND VGND
+ VPWR VPWR _03303_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_52_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18884_ _04181_ _04182_ _04180_ net255 VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__o22a_1
XFILLER_0_218_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17835_ decode.regfile.registers_6\[26\] _10603_ _12615_ _03231_ _03235_ VGND VGND
+ VPWR VPWR _03236_ sky130_fd_sc_hd__o32a_1
XFILLER_0_206_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer18 net242 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_1
X_17766_ decode.regfile.registers_17\[24\] _12580_ _03150_ _03168_ VGND VGND VPWR
+ VPWR _03169_ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14978_ _10948_ _10954_ _10997_ net451 _10999_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__o311a_1
Xrebuffer29 net255 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19505_ _04181_ net285 _04253_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__mux2_1
X_16717_ _12681_ VGND VGND VPWR VPWR _12682_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_187_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13929_ _10048_ _10210_ VGND VGND VPWR VPWR _10217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17697_ _13339_ _03099_ _03100_ _03101_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19436_ _04715_ _04722_ net351 _04723_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16648_ decode.immGen._imm_T_24\[19\] _10597_ _10934_ VGND VGND VPWR VPWR _12613_
+ sky130_fd_sc_hd__or3_4
XFILLER_0_202_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19367_ _04652_ _04654_ _04656_ _04657_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16579_ _12543_ VGND VGND VPWR VPWR _12544_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18318_ _03624_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19298_ _04045_ _04070_ _04274_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer108 net334 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_1
Xrebuffer119 net345 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18249_ _03582_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__buf_2
XFILLER_0_199_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21260_ net1128 _06132_ _06120_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold501 decode.regfile.registers_18\[12\] VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold512 decode.regfile.registers_3\[1\] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20211_ decode.id_ex_imm_reg\[30\] decode.id_ex_pc_reg\[30\] VGND VGND VPWR VPWR
+ _05407_ sky130_fd_sc_hd__nand2_1
Xhold523 decode.regfile.registers_29\[19\] VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 decode.regfile.registers_7\[11\] VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__dlygate4sd3_1
X_21191_ _06086_ _06082_ net1847 VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__and3_1
Xhold545 decode.regfile.registers_4\[4\] VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold556 decode.regfile.registers_23\[21\] VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold567 fetch.bht.bhtTable_tag\[2\]\[15\] VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20142_ _05345_ _05348_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__xnor2_1
Xhold578 decode.regfile.registers_28\[3\] VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold589 decode.regfile.registers_19\[5\] VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20073_ decode.id_ex_imm_reg\[11\] _10689_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__nor2_1
X_24950_ net1109 _08678_ net502 VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_202_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 fetch.bht.bhtTable_target_pc\[15\]\[26\] VGND VGND VPWR VPWR net1428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 fetch.bht.bhtTable_target_pc\[10\]\[6\] VGND VGND VPWR VPWR net1439 sky130_fd_sc_hd__dlygate4sd3_1
X_23901_ _08120_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_198_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_198_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 fetch.bht.bhtTable_tag\[1\]\[2\] VGND VGND VPWR VPWR net1450 sky130_fd_sc_hd__dlygate4sd3_1
X_24881_ csr.mcycle\[28\] csr.mcycle\[27\] csr.mcycle\[29\] _08630_ VGND VGND VPWR
+ VPWR _08631_ sky130_fd_sc_hd__and4_1
Xhold1234 fetch.bht.bhtTable_tag\[3\]\[4\] VGND VGND VPWR VPWR net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1245 fetch.bht.bhtTable_tag\[2\]\[5\] VGND VGND VPWR VPWR net1472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26620_ net2117 _09665_ _09667_ _09660_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__o211a_1
Xhold1256 decode.regfile.registers_4\[7\] VGND VGND VPWR VPWR net1483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23832_ _08075_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__clkbuf_1
Xhold1267 fetch.bht.bhtTable_target_pc\[13\]\[3\] VGND VGND VPWR VPWR net1494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1278 fetch.bht.bhtTable_tag\[14\]\[25\] VGND VGND VPWR VPWR net1505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1289 fetch.bht.bhtTable_target_pc\[11\]\[16\] VGND VGND VPWR VPWR net1516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23763_ _08033_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26551_ net716 _09622_ _09627_ _09619_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__o211a_1
X_20975_ execute.io_reg_pc\[13\] _05965_ _05961_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25502_ net2450 _09008_ _09009_ _09004_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22714_ net2803 _07236_ VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__or2_1
X_29270_ clknet_leaf_232_clock _02283_ VGND VGND VPWR VPWR decode.regfile.registers_0\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23694_ _07997_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__clkbuf_1
X_26482_ net1854 _09578_ _09587_ _09582_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28221_ clknet_leaf_86_clock net724 VGND VGND VPWR VPWR csr.mscratch\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22645_ net2762 _07205_ _07206_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__o21ba_1
X_25433_ _10121_ VGND VGND VPWR VPWR _08966_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_65_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_65_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28152_ clknet_leaf_169_clock _01174_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25364_ _09998_ VGND VGND VPWR VPWR _08918_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22576_ csr._minstret_T_3\[40\] csr._minstret_T_3\[32\] _07157_ _07159_ VGND VGND
+ VPWR VPWR _07160_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27103_ clknet_leaf_348_clock _00132_ VGND VGND VPWR VPWR decode.regfile.registers_25\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_24315_ _08333_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__clkbuf_1
X_21527_ _10557_ _09900_ _06281_ _10556_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__or4b_4
X_28083_ clknet_leaf_205_clock _01105_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_25295_ _08869_ net2578 VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24246_ _08074_ net1475 _08289_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__mux2_1
X_27034_ clknet_5_4__leaf_clock _00063_ VGND VGND VPWR VPWR decode.regfile.registers_23\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_21458_ _06149_ net1851 _06241_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20409_ csr.mcycle\[0\] _05552_ _05553_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24177_ _08262_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_187_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21389_ _06207_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_187_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23128_ net226 _07530_ net225 VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__a21oi_1
X_28985_ clknet_leaf_127_clock _01998_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_183_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput76 net76 VGND VGND VPWR VPWR io_fetch_address[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_183_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput87 net87 VGND VGND VPWR VPWR io_fetch_address[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_183_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27936_ clknet_leaf_214_clock _00958_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_23059_ csr._csr_read_data_T_8\[10\] _06039_ csr.io_mret_vector\[10\] _06463_ VGND
+ VGND VPWR VPWR _07502_ sky130_fd_sc_hd__a22o_1
X_15950_ _11059_ _11149_ _11128_ decode.regfile.registers_17\[16\] _11930_ VGND VGND
+ VPWR VPWR _11931_ sky130_fd_sc_hd__o221a_1
Xoutput98 net98 VGND VGND VPWR VPWR io_fetch_address[9] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_125_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14901_ _10935_ VGND VGND VPWR VPWR _10936_ sky130_fd_sc_hd__buf_2
X_15881_ decode.regfile.registers_23\[14\] _11262_ _11836_ _11863_ _11335_ VGND VGND
+ VPWR VPWR _11864_ sky130_fd_sc_hd__o221a_1
X_27867_ clknet_leaf_327_clock _00896_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17620_ _13183_ _03024_ _03025_ _03026_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__a31o_1
X_29606_ clknet_leaf_276_clock _02619_ VGND VGND VPWR VPWR decode.regfile.registers_11\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2480 decode.id_ex_rs1_data_reg\[9\] VGND VGND VPWR VPWR net2707 sky130_fd_sc_hd__dlygate4sd3_1
X_14832_ _10804_ _10873_ VGND VGND VPWR VPWR _10875_ sky130_fd_sc_hd__nand2_1
X_26818_ _09422_ _09776_ VGND VGND VPWR VPWR _09781_ sky130_fd_sc_hd__nand2_1
Xhold2491 decode.regfile.registers_13\[22\] VGND VGND VPWR VPWR net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_18_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_4_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27798_ clknet_leaf_335_clock _00827_ VGND VGND VPWR VPWR memory.io_wb_readdata\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1790 fetch.bht.bhtTable_tag\[15\]\[2\] VGND VGND VPWR VPWR net2017 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _12934_ _10592_ _12558_ decode.regfile.registers_0\[19\] VGND VGND VPWR VPWR
+ _02959_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29537_ clknet_leaf_251_clock _02550_ VGND VGND VPWR VPWR decode.regfile.registers_9\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_14763_ decode.id_ex_pc_reg\[17\] VGND VGND VPWR VPWR _10806_ sky130_fd_sc_hd__clkbuf_4
X_26749_ _09428_ _09733_ VGND VGND VPWR VPWR _09741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16502_ _11070_ _11470_ _11509_ decode.regfile.registers_10\[31\] _12467_ VGND VGND
+ VPWR VPWR _12468_ sky130_fd_sc_hd__a221o_1
XFILLER_0_224_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13714_ memory.csr_read_data_out_reg\[16\] _09987_ _10061_ _10062_ VGND VGND VPWR
+ VPWR _10063_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17482_ decode.regfile.registers_9\[17\] _12606_ _13428_ _13429_ VGND VGND VPWR VPWR
+ _13430_ sky130_fd_sc_hd__a22o_1
X_29468_ clknet_leaf_250_clock _02481_ VGND VGND VPWR VPWR decode.regfile.registers_7\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14694_ execute.io_target_pc\[17\] _10736_ _10688_ _10689_ VGND VGND VPWR VPWR _10737_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19221_ _04038_ _04054_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__and2_2
XFILLER_0_116_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28419_ clknet_leaf_39_clock _01432_ VGND VGND VPWR VPWR decode.immGen._imm_T_10\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16433_ decode.regfile.registers_15\[29\] _11036_ _11205_ _11208_ decode.regfile.registers_14\[29\]
+ VGND VGND VPWR VPWR _12401_ sky130_fd_sc_hd__a32o_1
XFILLER_0_195_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13645_ _09943_ VGND VGND VPWR VPWR _10003_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_183_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29399_ clknet_leaf_258_clock _02412_ VGND VGND VPWR VPWR decode.regfile.registers_4\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19152_ _04006_ _03983_ _03988_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_45_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16364_ decode.regfile.registers_18\[27\] _11269_ _11271_ _12333_ VGND VGND VPWR
+ VPWR _12334_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13576_ _09939_ _09940_ VGND VGND VPWR VPWR _09941_ sky130_fd_sc_hd__nand2_2
XFILLER_0_137_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18103_ _03469_ _03467_ _03474_ decode.io_id_pc\[9\] VGND VGND VPWR VPWR _03478_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_109_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15315_ decode.regfile.registers_8\[1\] _11285_ _11287_ _11310_ VGND VGND VPWR VPWR
+ _11311_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19083_ _04233_ _04180_ _04380_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16295_ _11050_ decode.regfile.registers_25\[25\] _11089_ VGND VGND VPWR VPWR _12267_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_87_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18034_ decode.regfile.registers_16\[31\] _12674_ _12901_ _03429_ VGND VGND VPWR
+ VPWR _03430_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15246_ _11242_ VGND VGND VPWR VPWR _11243_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_83_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15177_ _11173_ VGND VGND VPWR VPWR _11174_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14128_ _10331_ VGND VGND VPWR VPWR _10333_ sky130_fd_sc_hd__clkbuf_4
X_19985_ net426 _05217_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14059_ net927 _10287_ _10293_ _10291_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__o211a_1
X_18936_ _03977_ _03979_ _03982_ _04234_ _03775_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__a311o_1
XFILLER_0_20_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_105_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18867_ decode.id_ex_rs1_data_reg\[10\] _03687_ _04156_ _03914_ _04159_ VGND VGND
+ VPWR VPWR _04166_ sky130_fd_sc_hd__o221a_4
XFILLER_0_94_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17818_ _12968_ _03217_ _03218_ _03219_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__a31o_1
X_18798_ execute.io_reg_pc\[13\] _03776_ net104 _03664_ VGND VGND VPWR VPWR _04097_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_171_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17749_ decode.regfile.registers_7\[24\] _12611_ _12623_ decode.regfile.registers_6\[24\]
+ _12888_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_178_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20760_ _03452_ _05425_ _05577_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__and3b_1
XFILLER_0_175_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19419_ _04268_ _04705_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20691_ _05809_ decode.id_ex_rs1_data_reg\[7\] _05798_ VGND VGND VPWR VPWR _05812_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_114_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22430_ fetch.bht.bhtTable_tag\[15\]\[12\] _06707_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22361_ net79 _06955_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24100_ net1454 execute.io_target_pc\[5\] _08221_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21312_ net1135 _10872_ _06157_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__mux2_1
X_25080_ csr._mcycle_T_2\[30\] _08704_ _08766_ csr.mcycle\[30\] VGND VGND VPWR VPWR
+ _08768_ sky130_fd_sc_hd__a211o_1
X_22292_ net75 VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24031_ _07990_ VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21243_ _06121_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold320 decode.regfile.registers_29\[15\] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold331 decode.regfile.registers_19\[12\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold342 csr.mcycle\[0\] VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 decode.regfile.registers_31\[0\] VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 decode.regfile.registers_24\[8\] VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21174_ _06081_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__clkbuf_1
Xhold375 decode.regfile.registers_29\[30\] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 decode.regfile.registers_16\[8\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold397 decode.regfile.registers_15\[8\] VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_225_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20125_ _05332_ _05333_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_225_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28770_ clknet_leaf_134_clock _01783_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25982_ _09285_ VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27721_ clknet_leaf_20_clock _00750_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_20056_ decode.id_ex_imm_reg\[7\] _10730_ _05272_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__a21oi_1
X_24933_ csr._mcycle_T_3\[46\] _08668_ _06318_ VGND VGND VPWR VPWR _08669_ sky130_fd_sc_hd__a21oi_1
Xhold1020 fetch.bht.bhtTable_target_pc\[2\]\[22\] VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 csr._minstret_T_3\[51\] VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 execute.csr_write_address_out_reg\[3\] VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27652_ clknet_leaf_48_clock net168 VGND VGND VPWR VPWR execute.io_reg_pc\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold1053 decode.regfile.registers_6\[20\] VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24864_ _06143_ net2094 _08388_ VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1064 fetch.bht.bhtTable_tag\[12\]\[18\] VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1075 fetch.bht.bhtTable_tag\[8\]\[21\] VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1086 fetch.bht.bhtTable_tag\[5\]\[24\] VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26603_ net2681 _09649_ _09656_ _09648_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__o211a_1
X_23815_ execute.io_target_pc\[7\] VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__buf_2
Xhold1097 decode.regfile.registers_30\[17\] VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__dlygate4sd3_1
X_27583_ clknet_leaf_171_clock _00612_ VGND VGND VPWR VPWR csr.io_mem_pc\[24\] sky130_fd_sc_hd__dfxtp_1
X_24795_ _08089_ net941 _08574_ VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29322_ clknet_leaf_225_clock _02335_ VGND VGND VPWR VPWR decode.regfile.registers_2\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_155_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26534_ net2502 _09605_ _09616_ _09608_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__o211a_1
X_23746_ _08024_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__clkbuf_1
X_20958_ _05960_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_81_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Left_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29253_ clknet_leaf_218_clock _02266_ VGND VGND VPWR VPWR decode.regfile.registers_0\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26465_ _09576_ VGND VGND VPWR VPWR _09577_ sky130_fd_sc_hd__clkbuf_4
X_23677_ _07987_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__clkbuf_1
X_20889_ _05923_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__clkbuf_1
X_28204_ clknet_leaf_68_clock net778 VGND VGND VPWR VPWR csr.mscratch\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25416_ _08954_ _08946_ VGND VGND VPWR VPWR _08955_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22628_ _07195_ VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__clkbuf_2
X_29184_ clknet_leaf_157_clock _02197_ VGND VGND VPWR VPWR fetch.btb.btbTable\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26396_ _09377_ _09535_ VGND VGND VPWR VPWR _09538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28135_ clknet_leaf_221_clock _01157_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22559_ net713 csr._minstret_T_3\[36\] _07144_ _07146_ _06336_ VGND VGND VPWR VPWR
+ _01259_ sky130_fd_sc_hd__a311oi_1
X_25347_ _08905_ VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_114_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15100_ _10628_ _11042_ _11082_ VGND VGND VPWR VPWR _11097_ sky130_fd_sc_hd__or3_4
XFILLER_0_134_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer9 net235 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_6
X_28066_ clknet_leaf_175_clock _01088_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_16080_ decode.regfile.registers_10\[20\] _11184_ _11181_ VGND VGND VPWR VPWR _12057_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25278_ _10018_ VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_79_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_185_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_185_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15031_ net449 _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27017_ clknet_leaf_342_clock _00046_ VGND VGND VPWR VPWR decode.regfile.registers_22\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24229_ _06217_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_141_Left_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19770_ _04442_ _03852_ _03839_ _04667_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__a31o_1
X_28968_ clknet_leaf_103_clock _01981_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16982_ _11017_ _12539_ _12502_ decode.regfile.registers_7\[5\] _12644_ VGND VGND
+ VPWR VPWR _12942_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_88_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18721_ _04015_ _04016_ _04017_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27919_ clknet_leaf_69_clock _00948_ VGND VGND VPWR VPWR csr.io_csr_write_address\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_15933_ _10660_ _10655_ _11297_ decode.regfile.registers_3\[16\] VGND VGND VPWR VPWR
+ _11914_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_144_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28899_ clknet_leaf_130_clock _01912_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18652_ execute.io_reg_pc\[20\] _03776_ _03664_ net112 _03950_ VGND VGND VPWR VPWR
+ _03951_ sky130_fd_sc_hd__o221a_1
X_15864_ _11042_ decode.regfile.registers_4\[14\] _10646_ _10628_ _11082_ VGND VGND
+ VPWR VPWR _11847_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_118_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17603_ _03009_ _12653_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__nand2_1
X_14815_ _10760_ _10792_ VGND VGND VPWR VPWR _10858_ sky130_fd_sc_hd__nor2_1
X_18583_ _03872_ _03881_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__and2_1
X_15795_ decode.regfile.registers_13\[12\] _10642_ _11187_ _11778_ _11779_ VGND VGND
+ VPWR VPWR _11780_ sky130_fd_sc_hd__a32o_1
XFILLER_0_188_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_150_Left_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17534_ _12691_ _13453_ _13479_ _13480_ VGND VGND VPWR VPWR _13481_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _10768_ _10788_ VGND VGND VPWR VPWR _10789_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17465_ _13099_ _13262_ _13182_ decode.regfile.registers_29\[16\] _13413_ VGND VGND
+ VPWR VPWR _13414_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14677_ decode.id_ex_pc_reg\[26\] VGND VGND VPWR VPWR _10720_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19204_ _04008_ _03976_ _04497_ _04498_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__o22ai_4
X_16416_ _11493_ decode.regfile.registers_22\[29\] _11450_ _10978_ _10991_ VGND VGND
+ VPWR VPWR _12384_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13628_ _09987_ VGND VGND VPWR VPWR _09988_ sky130_fd_sc_hd__buf_8
XFILLER_0_73_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17396_ decode.regfile.registers_3\[15\] _12628_ _10609_ _12625_ VGND VGND VPWR VPWR
+ _13346_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19135_ _04335_ _04340_ _04247_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16347_ _12315_ _11371_ _10646_ _11298_ _12316_ VGND VGND VPWR VPWR _12317_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13559_ net132 net327 _09922_ _09925_ VGND VGND VPWR VPWR _09926_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_27_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19066_ _03835_ _03812_ _03989_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16278_ decode.regfile.registers_7\[25\] _11462_ _11297_ decode.regfile.registers_6\[25\]
+ _11534_ VGND VGND VPWR VPWR _12250_ sky130_fd_sc_hd__o32a_1
XFILLER_0_125_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18017_ _12934_ _10592_ _12558_ decode.regfile.registers_0\[31\] VGND VGND VPWR VPWR
+ _03413_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15229_ _11059_ _11065_ _11225_ _11085_ VGND VGND VPWR VPWR _11226_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19968_ _10694_ _05214_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__and2_1
XFILLER_0_226_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18919_ net349 _03809_ _04217_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__o21a_1
X_19899_ _05166_ _05167_ _04620_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_220_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21930_ csr.io_mret_vector\[28\] _10771_ _06539_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__mux2_1
X_21861_ _06511_ _06494_ _06495_ _06512_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23600_ _06130_ net1205 _07941_ VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20812_ _05881_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24580_ net1790 execute.io_target_pc\[12\] _08462_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__mux2_1
X_21792_ _06461_ _10970_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__and2_2
XFILLER_0_136_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23531_ net2793 _07903_ _07908_ _07907_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20743_ _05831_ _05813_ decode.id_ex_rs1_data_reg\[28\] _05842_ _00715_ VGND VGND
+ VPWR VPWR _00747_ sky130_fd_sc_hd__a32o_1
XFILLER_0_175_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23462_ _11015_ _07862_ _07859_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26250_ _09381_ _09448_ VGND VGND VPWR VPWR _09454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20674_ _05798_ _05799_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_189_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_189_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25201_ _08829_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__clkbuf_1
X_22413_ fetch.bht.bhtTable_tag\[0\]\[1\] fetch.bht.bhtTable_tag\[1\]\[1\] fetch.bht.bhtTable_tag\[2\]\[1\]
+ fetch.bht.bhtTable_tag\[3\]\[1\] _06680_ _06684_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23393_ csr._csr_read_data_T_8\[29\] _07416_ csr.io_mret_vector\[29\] _07417_ _07816_
+ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__o221a_1
X_26181_ _10057_ VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25132_ _08794_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__clkbuf_1
X_22344_ _06730_ _06938_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__and2b_1
XFILLER_0_190_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25063_ net1911 _08754_ _08755_ _06327_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__a211oi_1
X_29940_ clknet_leaf_341_clock _02953_ VGND VGND VPWR VPWR decode.regfile.registers_21\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_227_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22275_ _06866_ _06868_ _06869_ _06632_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_227_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24014_ _08178_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21226_ net841 _06109_ _09912_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__mux2_1
Xhold150 io_fetch_data[27] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29871_ clknet_leaf_300_clock _02884_ VGND VGND VPWR VPWR decode.regfile.registers_19\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold161 fetch.bht.bhtTable_valid\[6\] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold172 decode.regfile.registers_31\[16\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_180_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold183 fetch.btb.btbTable\[9\]\[0\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
X_28822_ clknet_leaf_126_clock _01835_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_180_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold194 fetch.btb.btbTable\[12\]\[0\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21157_ _06072_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20108_ decode.id_ex_imm_reg\[16\] decode.id_ex_pc_reg\[16\] VGND VGND VPWR VPWR
+ _05319_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_70_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28753_ clknet_leaf_104_clock _01766_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21088_ net328 net132 _09922_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__a21oi_1
X_25965_ _08962_ _09267_ VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__nand2_1
X_27704_ clknet_leaf_20_clock _00733_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_20039_ decode.id_ex_imm_reg\[6\] _10678_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24916_ net524 _08656_ csr._mcycle_T_3\[40\] VGND VGND VPWR VPWR _08658_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_107_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28684_ clknet_leaf_87_clock _01697_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_107_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25896_ _08968_ _09198_ VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27635_ clknet_leaf_45_clock net176 VGND VGND VPWR VPWR execute.io_reg_pc\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24847_ _08611_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_40 _08956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_51 _10041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_62 _10121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_178_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _10642_ decode.id_ex_ex_rd_reg\[0\] VGND VGND VPWR VPWR _10643_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_73 _10240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27566_ clknet_leaf_158_clock _00595_ VGND VGND VPWR VPWR csr.io_mem_pc\[7\] sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_84 _10594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15580_ _11344_ net508 _11528_ _11570_ _11249_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__o221a_1
X_24778_ _08575_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__clkbuf_1
XINSDIODE1_95 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29305_ clknet_leaf_242_clock _02318_ VGND VGND VPWR VPWR decode.regfile.registers_1\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14531_ _10574_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__clkbuf_1
X_26517_ _09566_ VGND VGND VPWR VPWR _09608_ sky130_fd_sc_hd__clkbuf_4
X_23729_ net1131 _10759_ _08014_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27497_ clknet_leaf_33_clock _00526_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29236_ clknet_leaf_181_clock _02249_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_17250_ decode.regfile.registers_17\[11\] _12719_ _13186_ _13203_ _12826_ VGND VGND
+ VPWR VPWR _13204_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_42_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26448_ _09428_ _09558_ VGND VGND VPWR VPWR _09568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14462_ net409 _10520_ _10525_ _10522_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ decode.regfile.registers_3\[23\] _11111_ _11142_ _11146_ VGND VGND VPWR VPWR
+ _12175_ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29167_ clknet_leaf_198_clock _02180_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_137_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17181_ _13099_ _12768_ _12493_ decode.regfile.registers_29\[9\] _13136_ VGND VGND
+ VPWR VPWR _13137_ sky130_fd_sc_hd__o221a_1
XFILLER_0_92_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26379_ net2099 _09518_ _09527_ _09525_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__o211a_1
X_14393_ net402 _10477_ _10485_ _10481_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28118_ clknet_leaf_89_clock net844 VGND VGND VPWR VPWR csr.minstret\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_180_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16132_ _11313_ decode.regfile.registers_4\[21\] _11191_ _10630_ _11462_ VGND VGND
+ VPWR VPWR _12108_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_3_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29098_ clknet_leaf_71_clock _02111_ VGND VGND VPWR VPWR csr._mcycle_T_3\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28049_ clknet_leaf_236_clock _01071_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16063_ _11106_ _12039_ _12040_ VGND VGND VPWR VPWR _12041_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_219_Left_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15014_ _11023_ VGND VGND VPWR VPWR _11024_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_184_Right_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19822_ _04330_ _05007_ _04304_ _05093_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_36_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16965_ decode.regfile.registers_18\[5\] _10925_ _12569_ _11023_ _11008_ VGND VGND
+ VPWR VPWR _12925_ sky130_fd_sc_hd__o2111a_1
X_19753_ _03851_ _05026_ _05027_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__a21o_1
X_15916_ _11094_ _11113_ _11119_ _11897_ VGND VGND VPWR VPWR _11898_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18704_ _03997_ _03998_ _03999_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__o2bb2a_1
X_19684_ _03947_ _03639_ _04667_ _04191_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__a211o_1
X_16896_ _12562_ _12856_ _12857_ _12545_ VGND VGND VPWR VPWR _12858_ sky130_fd_sc_hd__o211a_1
X_18635_ _03909_ _03914_ _03908_ decode.id_ex_rs1_data_reg\[17\] _03910_ VGND VGND
+ VPWR VPWR _03934_ sky130_fd_sc_hd__o221a_4
XFILLER_0_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15847_ _11403_ _11828_ _11829_ _11830_ VGND VGND VPWR VPWR _11831_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_228_Left_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18566_ _03862_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__nor2_1
X_15778_ _11446_ decode.regfile.registers_26\[12\] _11447_ _11348_ _10993_ VGND VGND
+ VPWR VPWR _11763_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17517_ decode.regfile.registers_9\[18\] _12602_ _13454_ _13463_ VGND VGND VPWR VPWR
+ _13464_ sky130_fd_sc_hd__o22ai_2
X_14729_ csr.io_mem_pc\[24\] VGND VGND VPWR VPWR _10772_ sky130_fd_sc_hd__buf_4
XFILLER_0_115_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18497_ net206 net207 VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__nor2_4
XFILLER_0_129_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17448_ _12555_ _10923_ _12876_ _13395_ _13396_ VGND VGND VPWR VPWR _13397_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17379_ _12716_ decode.regfile.registers_21\[14\] _12909_ _13329_ VGND VGND VPWR
+ VPWR _13330_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19118_ _04242_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20390_ _05550_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__clkbuf_1
X_19049_ _04242_ _04293_ _04295_ _04315_ _04347_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__a311o_1
XFILLER_0_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22060_ _06639_ _06629_ _06642_ _06654_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__a211o_1
XFILLER_0_207_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21011_ execute.io_reg_pc\[29\] _05989_ _05985_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_222_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_222_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25750_ net2091 _09112_ _09151_ _09142_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__o211a_1
X_22962_ net93 net92 net89 VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__and3_1
XFILLER_0_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24701_ _08534_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21913_ net1093 _06545_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__or2_1
X_25681_ _09025_ _09112_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22893_ _03500_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27420_ clknet_leaf_9_clock _00449_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[29\]
+ sky130_fd_sc_hd__dfxtp_2
X_24632_ net1040 execute.io_target_pc\[5\] _08497_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21844_ csr.io_mret_vector\[2\] _10556_ _06040_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27351_ clknet_leaf_46_clock _00380_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[24\]
+ sky130_fd_sc_hd__dfxtp_2
X_21775_ net1016 _10760_ _06450_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__mux2_1
X_24563_ _08463_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_216_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26302_ _09434_ _09472_ VGND VGND VPWR VPWR _09483_ sky130_fd_sc_hd__nand2_1
X_23514_ net2769 _07890_ _07887_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__or3b_1
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20726_ _05809_ decode.id_ex_rs1_data_reg\[21\] _03585_ VGND VGND VPWR VPWR _05833_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27282_ clknet_leaf_33_clock _00311_ VGND VGND VPWR VPWR decode.regfile.registers_31\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24494_ _08427_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29021_ clknet_leaf_179_clock _02034_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26233_ net1587 _09374_ _09442_ _09440_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20657_ _05785_ _05786_ _03595_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__o21a_2
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23445_ net3 _07846_ _07857_ _07851_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23376_ execute.io_target_pc\[28\] _07090_ _07089_ _07800_ _06032_ VGND VGND VPWR
+ VPWR _07801_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26164_ net2761 _09373_ _09393_ _09394_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__o211a_1
X_20588_ _05627_ csr.io_mret_vector\[20\] _05603_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25115_ _06132_ net1905 _08778_ VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22327_ _06672_ _06921_ _06635_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26095_ _08941_ _09340_ VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22258_ fetch.bht.bhtTable_tag\[6\]\[17\] fetch.bht.bhtTable_tag\[7\]\[17\] _06616_
+ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__mux2_1
X_25046_ csr._mcycle_T_2\[20\] _08712_ _08742_ _03554_ net2733 VGND VGND VPWR VPWR
+ _08744_ sky130_fd_sc_hd__a221oi_1
X_29923_ clknet_leaf_335_clock _02936_ VGND VGND VPWR VPWR decode.regfile.registers_21\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21209_ _06099_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__clkbuf_1
X_29854_ clknet_leaf_305_clock _02867_ VGND VGND VPWR VPWR decode.regfile.registers_19\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_22189_ _06740_ _06773_ _06777_ _06783_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_109_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28805_ clknet_leaf_135_clock _01818_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_29785_ clknet_leaf_313_clock _02798_ VGND VGND VPWR VPWR decode.regfile.registers_16\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_26997_ clknet_leaf_333_clock _00026_ VGND VGND VPWR VPWR decode.regfile.registers_22\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_28736_ clknet_leaf_170_clock _01749_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16750_ _11013_ _10935_ _12667_ _10595_ VGND VGND VPWR VPWR _12714_ sky130_fd_sc_hd__or4_4
X_13962_ net2485 _10226_ _10235_ _10232_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_31_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25948_ net2240 _09256_ _09266_ _09264_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15701_ decode.regfile.registers_18\[10\] _10955_ _11114_ _11094_ _10977_ VGND VGND
+ VPWR VPWR _11688_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_220_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28667_ clknet_leaf_135_clock _01680_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_16681_ _12497_ _12539_ _12503_ decode.regfile.registers_7\[0\] _12645_ VGND VGND
+ VPWR VPWR _12646_ sky130_fd_sc_hd__o32a_1
XFILLER_0_216_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25879_ _08952_ _09223_ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__nand2_1
X_13893_ decode.io_wb_rd\[3\] VGND VGND VPWR VPWR _10194_ sky130_fd_sc_hd__buf_12
X_18420_ csr.io_csr_address\[3\] VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__inv_2
X_27618_ clknet_leaf_149_clock _00647_ VGND VGND VPWR VPWR execute.io_target_pc\[27\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15632_ decode.regfile.registers_5\[8\] _10637_ _11139_ _11619_ _11620_ VGND VGND
+ VPWR VPWR _11621_ sky130_fd_sc_hd__a32o_1
X_28598_ clknet_leaf_125_clock _01611_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_305 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_316 decode.regfile.registers_12\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_327 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18351_ execute.io_mem_regwrite decode.id_ex_ex_use_rs1_reg VGND VGND VPWR VPWR _03650_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_139_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ decode.regfile.registers_16\[6\] _11123_ _11531_ _11553_ VGND VGND VPWR VPWR
+ _11554_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_338 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27549_ clknet_leaf_43_clock _00578_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_349 _03580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17302_ _13087_ decode.regfile.registers_26\[12\] _13254_ _13047_ _13088_ VGND VGND
+ VPWR VPWR _13255_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_51_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14514_ _10555_ _09917_ _09916_ _10558_ VGND VGND VPWR VPWR _10559_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ decode.id_ex_rs2_data_reg\[7\] _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15494_ _11075_ _11482_ _11485_ _11486_ VGND VGND VPWR VPWR _11487_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29219_ clknet_leaf_93_clock _02232_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17233_ decode.regfile.registers_14\[11\] _10619_ _12589_ _10612_ VGND VGND VPWR
+ VPWR _13187_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14445_ net508 _10506_ _10515_ _10509_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17164_ decode.regfile.registers_16\[9\] _12576_ _13101_ _13119_ VGND VGND VPWR VPWR
+ _13120_ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14376_ _10025_ _10474_ VGND VGND VPWR VPWR _10476_ sky130_fd_sc_hd__nand2_1
X_16115_ _11756_ decode.regfile.registers_28\[20\] _11871_ _11681_ _11448_ VGND VGND
+ VPWR VPWR _12092_ sky130_fd_sc_hd__o2111a_1
Xhold908 fetch.bht.bhtTable_tag\[1\]\[8\] VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold919 fetch.bht.bhtTable_target_pc\[14\]\[16\] VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17095_ _12496_ _13049_ _13051_ _13052_ VGND VGND VPWR VPWR _13053_ sky130_fd_sc_hd__a31o_1
XFILLER_0_161_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16046_ _11298_ _10646_ _12022_ _12023_ VGND VGND VPWR VPWR _12024_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_126_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2309 _01139_ VGND VGND VPWR VPWR net2536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19805_ _05076_ _05052_ _03814_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__o21ai_1
Xhold1608 _01235_ VGND VGND VPWR VPWR net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_17997_ _10604_ _10619_ _12773_ _03380_ _03393_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__o32a_1
XFILLER_0_193_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1619 fetch.bht.bhtTable_tag\[10\]\[6\] VGND VGND VPWR VPWR net1846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19736_ _04618_ _04245_ _04386_ _04515_ _03705_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__o32a_1
X_16948_ _12755_ VGND VGND VPWR VPWR _12909_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19667_ _04790_ _04249_ _04272_ _04848_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__a211o_1
X_16879_ _12832_ _12839_ _12840_ VGND VGND VPWR VPWR _12841_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18618_ _03817_ _03916_ _03774_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_204_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19598_ _04317_ _04393_ _04879_ _04539_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18549_ _03844_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21560_ _06300_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20511_ _05540_ csr.io_mret_vector\[10\] _05602_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_220_Right_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21491_ _06262_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_211_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23230_ _07371_ _07661_ _07663_ _06637_ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20442_ _05527_ _05540_ _05524_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_891 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23161_ csr._csr_read_data_T_8\[15\] _06461_ csr.io_mret_vector\[15\] _07417_ _07598_
+ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20373_ csr.io_csr_address\[9\] _05535_ csr.io_csr_address\[11\] csr.io_csr_address\[10\]
+ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_144_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22112_ _06706_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__buf_4
X_23092_ execute.io_target_pc\[11\] _07346_ _07521_ _07533_ _07348_ VGND VGND VPWR
+ VPWR _07534_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_2_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22043_ _06633_ _06634_ _06637_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__a21o_1
X_26920_ _09838_ VGND VGND VPWR VPWR _09840_ sky130_fd_sc_hd__buf_2
XFILLER_0_101_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26851_ net993 _09795_ _09800_ _09799_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25802_ net2553 _09170_ _09181_ _09182_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29570_ clknet_leaf_270_clock _02583_ VGND VGND VPWR VPWR decode.regfile.registers_10\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_26782_ net816 _09752_ _09760_ _09758_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23994_ net1023 VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28521_ clknet_leaf_167_clock _01534_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25733_ _08956_ _09136_ VGND VGND VPWR VPWR _09143_ sky130_fd_sc_hd__nand2_1
X_22945_ _07391_ _07392_ _07393_ _07394_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_134_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28452_ clknet_leaf_146_clock _01465_ VGND VGND VPWR VPWR decode.io_id_pc\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25664_ net2594 _09095_ _09102_ _09100_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__o211a_1
X_22876_ _07334_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27403_ clknet_leaf_29_clock _00432_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_24615_ net871 execute.io_target_pc\[29\] _09897_ VGND VGND VPWR VPWR _08490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28383_ clknet_leaf_55_clock _01396_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_4
X_21827_ _06481_ net734 _06316_ _06470_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25595_ net2605 _09052_ _09062_ _09059_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27334_ clknet_leaf_46_clock _00363_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24546_ _08454_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21758_ net1388 csr.io_mem_pc\[18\] _06439_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20709_ _05822_ _05823_ _05414_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__o21a_1
X_27265_ clknet_leaf_0_clock _00294_ VGND VGND VPWR VPWR decode.regfile.registers_30\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_24477_ _08418_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__clkbuf_1
X_21689_ net526 _06321_ _06392_ csr.minstret\[25\] VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_34_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29004_ clknet_leaf_109_clock _02017_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ _10036_ _10387_ VGND VGND VPWR VPWR _10392_ sky130_fd_sc_hd__nand2_1
X_26216_ _09430_ _09413_ VGND VGND VPWR VPWR _09431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23428_ net23 _07846_ _07848_ _05454_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_24_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27196_ clknet_leaf_360_clock _00225_ VGND VGND VPWR VPWR decode.regfile.registers_28\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire168 _00681_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire179 net180 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14161_ net2557 _10346_ _10351_ _10344_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26147_ net1812 _09373_ _09382_ _09370_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__o211a_1
X_23359_ _07783_ _07784_ _07063_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_95_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14092_ net2069 _10302_ _10311_ _10304_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__o211a_1
X_26078_ net1137 _09329_ _09341_ _09333_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_91_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25029_ csr.mcycle\[14\] csr.mcycle\[13\] _08730_ VGND VGND VPWR VPWR _08733_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_363_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_363_clock
+ sky130_fd_sc_hd__clkbuf_8
X_17920_ decode.regfile.registers_12\[28\] _12489_ _11019_ _12540_ VGND VGND VPWR
+ VPWR _03319_ sky130_fd_sc_hd__or4_1
X_29906_ clknet_leaf_340_clock _02919_ VGND VGND VPWR VPWR decode.regfile.registers_20\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17851_ _03250_ _03251_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_128_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29837_ clknet_leaf_298_clock _02850_ VGND VGND VPWR VPWR decode.regfile.registers_18\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16802_ _10930_ VGND VGND VPWR VPWR _12765_ sky130_fd_sc_hd__buf_4
X_17782_ net478 _12872_ _03147_ _03184_ _03073_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__o221a_1
X_14994_ _10931_ _11004_ _11006_ _11007_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__a31o_1
X_29768_ clknet_leaf_293_clock _02781_ VGND VGND VPWR VPWR decode.regfile.registers_16\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_19521_ _04346_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__clkbuf_4
X_16733_ _12697_ VGND VGND VPWR VPWR _12698_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28719_ clknet_leaf_111_clock _01732_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13945_ _10198_ VGND VGND VPWR VPWR _10226_ sky130_fd_sc_hd__clkbuf_4
X_29699_ clknet_leaf_291_clock _02712_ VGND VGND VPWR VPWR decode.regfile.registers_14\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19452_ _04149_ _04152_ _04166_ _04164_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16664_ _12628_ VGND VGND VPWR VPWR _12629_ sky130_fd_sc_hd__buf_4
X_13876_ _10107_ _10177_ VGND VGND VPWR VPWR _10185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_102 _10668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_5__f_clock clknet_2_0_0_clock VGND VGND VPWR VPWR clknet_5_5__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_15615_ _11236_ _11602_ _11603_ _11604_ VGND VGND VPWR VPWR _11605_ sky130_fd_sc_hd__a31o_1
X_18403_ decode.id_ex_rs1_data_reg\[31\] _03689_ _03690_ _03701_ VGND VGND VPWR VPWR
+ _03702_ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_301_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_301_clock
+ sky130_fd_sc_hd__clkbuf_8
XINSDIODE1_113 _11036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19383_ _04251_ _04252_ _04671_ _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__a31o_1
XINSDIODE1_124 _11149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16595_ _11020_ _12555_ _10923_ _12559_ VGND VGND VPWR VPWR _12560_ sky130_fd_sc_hd__and4_1
XINSDIODE1_135 _11549_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_146 _12512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18334_ decode.id_ex_aluop_reg\[1\] VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__clkbuf_4
XINSDIODE1_157 _12690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15546_ decode.regfile.registers_2\[6\] _11155_ _11150_ _11120_ VGND VGND VPWR VPWR
+ _11537_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_29_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_168 decode.id_ex_rs1_data_reg\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_179 execute.io_reg_pc\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18265_ _03595_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15477_ _11167_ VGND VGND VPWR VPWR _11470_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17216_ _10927_ decode.regfile.registers_24\[10\] _13170_ _13083_ _12862_ VGND VGND
+ VPWR VPWR _13171_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_4_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_316_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_316_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14428_ _10504_ VGND VGND VPWR VPWR _10505_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18196_ _10965_ _10964_ _10951_ _10946_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__o31a_1
XFILLER_0_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17147_ _12934_ _12616_ _12557_ decode.regfile.registers_0\[9\] VGND VGND VPWR VPWR
+ _13103_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold705 fetch.bht.bhtTable_tag\[3\]\[14\] VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14359_ net665 _10463_ _10466_ _10453_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__o211a_1
Xhold716 fetch.bht.bhtTable_tag\[8\]\[8\] VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 fetch.bht.bhtTable_target_pc\[2\]\[21\] VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold738 fetch.bht.bhtTable_target_pc\[3\]\[2\] VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold749 fetch.bht.bhtTable_target_pc\[1\]\[0\] VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17078_ decode.regfile.registers_18\[7\] _12566_ _12678_ _13035_ VGND VGND VPWR VPWR
+ _13036_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16029_ decode.regfile.registers_21\[18\] _11062_ _11100_ _11229_ _12007_ VGND VGND
+ VPWR VPWR _12008_ sky130_fd_sc_hd__o311a_1
XFILLER_0_23_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2106 decode.regfile.registers_25\[5\] VGND VGND VPWR VPWR net2333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2117 decode.regfile.registers_6\[22\] VGND VGND VPWR VPWR net2344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2128 decode.regfile.registers_20\[28\] VGND VGND VPWR VPWR net2355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2139 _03574_ VGND VGND VPWR VPWR net2366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1405 fetch.bht.bhtTable_target_pc\[9\]\[12\] VGND VGND VPWR VPWR net1632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 fetch.bht.bhtTable_target_pc\[9\]\[24\] VGND VGND VPWR VPWR net1643 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1427 fetch.bht.bhtTable_target_pc\[0\]\[28\] VGND VGND VPWR VPWR net1654 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1438 fetch.bht.bhtTable_tag\[7\]\[8\] VGND VGND VPWR VPWR net1665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1449 fetch.bht.bhtTable_target_pc\[5\]\[12\] VGND VGND VPWR VPWR net1676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19719_ _04194_ _03882_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__or2_2
X_20991_ execute.io_reg_pc\[20\] _05977_ _05973_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__and3_1
XFILLER_0_205_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22730_ _07257_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22661_ net2235 _07208_ _07216_ _07164_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_213_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24400_ _08377_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_213_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21612_ _05613_ _06323_ _06333_ _06335_ _06336_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__a311oi_1
X_25380_ _08929_ _08923_ VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1003 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22592_ csr._minstret_T_3\[45\] _07170_ _07171_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_36_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24331_ _08093_ net1363 _08334_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21543_ _06291_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27050_ clknet_leaf_342_clock _00079_ VGND VGND VPWR VPWR decode.regfile.registers_23\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_24262_ _08306_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__clkbuf_1
X_21474_ _06103_ net1649 _06252_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26001_ _09285_ VGND VGND VPWR VPWR _09297_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23213_ _07130_ _07637_ _07647_ _07090_ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__a211o_1
X_20425_ csr.io_mret_vector\[1\] _05580_ _05581_ csr.mscratch\[1\] _05583_ VGND VGND
+ VPWR VPWR _05584_ sky130_fd_sc_hd__a221o_1
X_24193_ _08087_ net1943 _08266_ VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23144_ net72 _07567_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__nor2_1
X_20356_ csr.io_csr_address\[4\] csr.io_csr_address\[5\] csr.io_csr_address\[7\] csr.io_csr_address\[6\]
+ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_164_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27952_ clknet_leaf_199_clock _00974_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_23075_ _07085_ _07508_ _07517_ _07130_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_164_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20287_ _05412_ _05318_ _05466_ _03517_ _03551_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_105_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22026_ _06620_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__buf_4
X_26903_ decode.regfile.registers_20\[25\] _09822_ _09829_ _09825_ VGND VGND VPWR
+ VPWR _02920_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27883_ clknet_leaf_65_clock _00912_ VGND VGND VPWR VPWR csr._mcycle_T_2\[4\] sky130_fd_sc_hd__dfxtp_2
X_29622_ clknet_leaf_280_clock _02635_ VGND VGND VPWR VPWR decode.regfile.registers_11\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_26834_ net2405 _09779_ _09789_ _09784_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1950 fetch.bht.bhtTable_tag\[10\]\[5\] VGND VGND VPWR VPWR net2177 sky130_fd_sc_hd__dlygate4sd3_1
X_29553_ clknet_leaf_274_clock _02566_ VGND VGND VPWR VPWR decode.regfile.registers_9\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_123_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1961 decode.regfile.registers_15\[13\] VGND VGND VPWR VPWR net2188 sky130_fd_sc_hd__dlygate4sd3_1
X_26765_ net2070 _09710_ _09749_ _09743_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__o211a_1
X_23977_ _08159_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_123_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1972 decode.regfile.registers_7\[0\] VGND VGND VPWR VPWR net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1983 decode.io_id_pc\[20\] VGND VGND VPWR VPWR net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28504_ clknet_leaf_219_clock _01517_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13730_ _10019_ VGND VGND VPWR VPWR _10077_ sky130_fd_sc_hd__buf_2
Xhold1994 decode.regfile.registers_13\[31\] VGND VGND VPWR VPWR net2221 sky130_fd_sc_hd__dlygate4sd3_1
X_25716_ _08939_ _09122_ VGND VGND VPWR VPWR _09133_ sky130_fd_sc_hd__nand2_1
X_22928_ _07372_ _07085_ _07378_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__a21oi_2
X_29484_ clknet_leaf_263_clock _02497_ VGND VGND VPWR VPWR decode.regfile.registers_7\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26696_ net2258 _09709_ _09711_ _09702_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28435_ clknet_leaf_49_clock _01448_ VGND VGND VPWR VPWR decode.control.io_funct7\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13661_ _09954_ VGND VGND VPWR VPWR _10018_ sky130_fd_sc_hd__buf_4
X_25647_ _08945_ _09092_ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22859_ net1685 _10868_ _07324_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15400_ _11076_ decode.regfile.registers_25\[2\] _11090_ _11235_ _11394_ VGND VGND
+ VPWR VPWR _11395_ sky130_fd_sc_hd__o311a_1
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28366_ clknet_leaf_212_clock _01379_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16380_ _11071_ _11204_ _11184_ decode.regfile.registers_10\[28\] VGND VGND VPWR
+ VPWR _12349_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25578_ net2394 _09052_ _09053_ _09046_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13592_ _09956_ VGND VGND VPWR VPWR _09957_ sky130_fd_sc_hd__buf_4
XFILLER_0_183_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15331_ _11221_ VGND VGND VPWR VPWR _11327_ sky130_fd_sc_hd__clkbuf_4
X_27317_ clknet_leaf_327_clock _00346_ VGND VGND VPWR VPWR decode.id_ex_ex_rd_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24529_ _08089_ net1369 _08439_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__mux2_1
X_28297_ clknet_leaf_164_clock _00015_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18050_ _10930_ _12767_ _12965_ decode.regfile.registers_29\[31\] _03445_ VGND VGND
+ VPWR VPWR _03446_ sky130_fd_sc_hd__o221a_1
X_15262_ _11257_ VGND VGND VPWR VPWR _11258_ sky130_fd_sc_hd__buf_2
X_27248_ clknet_leaf_7_clock _00277_ VGND VGND VPWR VPWR decode.regfile.registers_30\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17001_ _10940_ _12706_ decode.regfile.registers_27\[5\] _12507_ VGND VGND VPWR VPWR
+ _12961_ sky130_fd_sc_hd__or4_1
XFILLER_0_227_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14213_ _09984_ _10377_ VGND VGND VPWR VPWR _10382_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_93_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15193_ _11129_ VGND VGND VPWR VPWR _11190_ sky130_fd_sc_hd__buf_4
X_27179_ clknet_leaf_361_clock _00208_ VGND VGND VPWR VPWR decode.regfile.registers_27\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14144_ net453 _10332_ _10341_ _10328_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14075_ _10286_ VGND VGND VPWR VPWR _10302_ sky130_fd_sc_hd__buf_2
X_18952_ _03997_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17903_ _10927_ decode.regfile.registers_24\[28\] _10933_ _12759_ _12862_ VGND VGND
+ VPWR VPWR _03302_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_197_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18883_ _04083_ _04084_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17834_ _10610_ _12626_ _12629_ decode.regfile.registers_3\[26\] _03234_ VGND VGND
+ VPWR VPWR _03235_ sky130_fd_sc_hd__o221a_2
XFILLER_0_20_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14977_ _10948_ _10954_ _10997_ net449 _10999_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__o311a_1
X_17765_ _12585_ _03166_ _03167_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__o21a_1
XFILLER_0_221_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer19 _03686_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__buf_1
XFILLER_0_18_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19504_ _04454_ _04783_ _04784_ _04788_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13928_ net627 _10213_ _10216_ _10206_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__o211a_1
X_16716_ _10595_ _10599_ _10935_ _12512_ VGND VGND VPWR VPWR _12681_ sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_240_clock clknet_5_25__leaf_clock VGND VGND VPWR VPWR clknet_leaf_240_clock
+ sky130_fd_sc_hd__clkbuf_8
X_17696_ _13250_ decode.regfile.registers_24\[22\] _13170_ _12998_ _13367_ VGND VGND
+ VPWR VPWR _03101_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_92_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16647_ _12611_ VGND VGND VPWR VPWR _12612_ sky130_fd_sc_hd__clkbuf_4
X_19435_ _04160_ _04164_ _04155_ _04721_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__a211o_1
X_13859_ net742 _10167_ _10174_ _10175_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19366_ _04271_ _04546_ _04295_ _04362_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__a211o_1
X_16578_ _10594_ _10598_ _10935_ _12542_ VGND VGND VPWR VPWR _12543_ sky130_fd_sc_hd__or4_4
XFILLER_0_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15529_ decode.regfile.registers_23\[5\] _11086_ _11495_ _11520_ _11335_ VGND VGND
+ VPWR VPWR _11521_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18317_ decode.id_ex_rs2_data_reg\[24\] _03616_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_255_clock clknet_5_19__leaf_clock VGND VGND VPWR VPWR clknet_leaf_255_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19297_ _04073_ _04070_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer109 _10761_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_178_Left_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18248_ _09954_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18179_ _10944_ _03516_ _03517_ _03518_ _10972_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold502 decode.regfile.registers_8\[11\] VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap210 _09974_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_4
X_20210_ _05178_ _05247_ _05406_ _05267_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_124_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold513 decode.regfile.registers_29\[23\] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold524 decode.regfile.registers_6\[11\] VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__dlygate4sd3_1
X_21190_ _06090_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold535 csr.minstret\[28\] VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 fetch.bht.bhtTable_target_pc\[1\]\[28\] VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold557 decode.regfile.registers_24\[0\] VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 csr.mscratch\[1\] VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__dlygate4sd3_1
X_20141_ decode.id_ex_imm_reg\[19\] _05340_ _05347_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_206_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold579 csr._mcycle_T_2\[14\] VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_1206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20072_ decode.id_ex_imm_reg\[11\] _10689_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__and2_1
Xhold1202 fetch.bht.bhtTable_target_pc\[0\]\[29\] VGND VGND VPWR VPWR net1429 sky130_fd_sc_hd__dlygate4sd3_1
X_23900_ net1253 _08057_ _08119_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_187_Left_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_198_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 fetch.bht.bhtTable_target_pc\[11\]\[24\] VGND VGND VPWR VPWR net1440 sky130_fd_sc_hd__dlygate4sd3_1
X_24880_ csr.mcycle\[23\] csr.mcycle\[26\] csr.mcycle\[25\] csr.mcycle\[30\] VGND
+ VGND VPWR VPWR _08630_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_198_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 fetch.bht.bhtTable_target_pc\[3\]\[3\] VGND VGND VPWR VPWR net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 fetch.bht.bhtTable_target_pc\[15\]\[13\] VGND VGND VPWR VPWR net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 fetch.bht.bhtTable_tag\[2\]\[10\] VGND VGND VPWR VPWR net1473 sky130_fd_sc_hd__dlygate4sd3_1
X_23831_ _08074_ net1670 _08058_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__mux2_1
Xhold1257 fetch.bht.bhtTable_target_pc\[7\]\[19\] VGND VGND VPWR VPWR net1484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1268 fetch.bht.bhtTable_target_pc\[7\]\[13\] VGND VGND VPWR VPWR net1495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1279 fetch.bht.bhtTable_target_pc\[7\]\[29\] VGND VGND VPWR VPWR net1506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_208_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_208_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26550_ _09379_ _09623_ VGND VGND VPWR VPWR _09627_ sky130_fd_sc_hd__nand2_1
X_23762_ _06124_ net1782 _08030_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20974_ _05969_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25501_ _08952_ _09005_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22713_ net2632 _07235_ _07245_ _07234_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26481_ _09385_ _09579_ VGND VGND VPWR VPWR _09587_ sky130_fd_sc_hd__nand2_1
X_23693_ net1461 _10878_ _07992_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28220_ clknet_leaf_86_clock net1094 VGND VGND VPWR VPWR csr.mscratch\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_157_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25432_ net577 _08951_ _08965_ _08950_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__o211a_1
X_22644_ csr._minstret_T_3\[63\] csr._minstret_T_3\[62\] csr._minstret_T_3\[61\] _07202_
+ _07148_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__a41o_1
XFILLER_0_211_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28151_ clknet_leaf_175_clock _01173_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_196_Left_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25363_ net2636 _08906_ _08917_ _07247_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22575_ csr._minstret_T_3\[38\] csr._minstret_T_3\[37\] csr._minstret_T_3\[36\] _07158_
+ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27102_ clknet_leaf_348_clock _00131_ VGND VGND VPWR VPWR decode.regfile.registers_25\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_24314_ _08076_ net1495 _08323_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28082_ clknet_leaf_204_clock _01104_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_21526_ _09879_ _09882_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__nand2_2
X_25294_ _08877_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27033_ clknet_leaf_350_clock _00062_ VGND VGND VPWR VPWR decode.regfile.registers_23\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24245_ _08297_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_116_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21457_ _06244_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20408_ csr._minstret_T_3\[32\] _05526_ _05536_ _05558_ _05567_ VGND VGND VPWR VPWR
+ _05568_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21388_ _06136_ net2039 _06199_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__mux2_1
X_24176_ _08070_ net1245 _08255_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23127_ net225 net226 _07530_ VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__and3_1
X_20339_ decode.id_ex_pc_reg\[28\] _05502_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28984_ clknet_leaf_122_clock _01997_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput77 net77 VGND VGND VPWR VPWR io_fetch_address[19] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput88 net88 VGND VGND VPWR VPWR io_fetch_address[29] sky130_fd_sc_hd__clkbuf_4
X_27935_ clknet_leaf_165_clock _00019_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_23058_ _06718_ _07343_ _07344_ _07501_ _06566_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__o311a_1
XFILLER_0_101_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput99 net99 VGND VGND VPWR VPWR io_load_store_unsigned sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_125_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14900_ _10934_ VGND VGND VPWR VPWR _10935_ sky130_fd_sc_hd__buf_4
X_22009_ csr._mcycle_T_2\[26\] _06600_ _06609_ _06605_ VGND VGND VPWR VPWR _01246_
+ sky130_fd_sc_hd__o211a_1
X_15880_ decode.regfile.registers_21\[14\] _11060_ _11098_ _11227_ _11862_ VGND VGND
+ VPWR VPWR _11863_ sky130_fd_sc_hd__o311a_1
X_27866_ clknet_leaf_324_clock _00895_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2470 decode.regfile.registers_14\[14\] VGND VGND VPWR VPWR net2697 sky130_fd_sc_hd__dlygate4sd3_1
X_14831_ _10804_ _10873_ _10675_ VGND VGND VPWR VPWR _10874_ sky130_fd_sc_hd__a21o_1
Xhold2481 csr._mcycle_T_2\[10\] VGND VGND VPWR VPWR net2708 sky130_fd_sc_hd__dlygate4sd3_1
X_29605_ clknet_leaf_276_clock _02618_ VGND VGND VPWR VPWR decode.regfile.registers_11\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_26817_ net2527 _09779_ _09780_ _09771_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__o211a_1
X_27797_ clknet_leaf_323_clock _00826_ VGND VGND VPWR VPWR memory.io_wb_readdata\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2492 decode.regfile.registers_9\[1\] VGND VGND VPWR VPWR net2719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1780 _01240_ VGND VGND VPWR VPWR net2007 sky130_fd_sc_hd__dlygate4sd3_1
X_17550_ decode.regfile.registers_2\[19\] _10609_ _12636_ _12639_ VGND VGND VPWR VPWR
+ _13496_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_86_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1791 fetch.bht.bhtTable_target_pc\[4\]\[30\] VGND VGND VPWR VPWR net2018 sky130_fd_sc_hd__dlygate4sd3_1
X_14762_ _10803_ _10804_ VGND VGND VPWR VPWR _10805_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_142_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26748_ net2299 _09736_ _09740_ _09730_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__o211a_1
X_29536_ clknet_leaf_312_clock _02549_ VGND VGND VPWR VPWR decode.regfile.registers_9\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_23__f_clock clknet_2_2_0_clock VGND VGND VPWR VPWR clknet_5_23__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_16501_ _11381_ _12465_ _12466_ VGND VGND VPWR VPWR _12467_ sky130_fd_sc_hd__and3_1
X_13713_ _10003_ memory.io_wb_aluresult\[16\] _10001_ memory.io_wb_reg_pc\[16\] _10005_
+ VGND VGND VPWR VPWR _10062_ sky130_fd_sc_hd__a221o_1
X_17481_ _11017_ _12502_ _12509_ decode.regfile.registers_8\[17\] _12725_ VGND VGND
+ VPWR VPWR _13429_ sky130_fd_sc_hd__o32a_1
X_29467_ clknet_leaf_253_clock _02480_ VGND VGND VPWR VPWR decode.regfile.registers_7\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14693_ decode.id_ex_pc_reg\[17\] VGND VGND VPWR VPWR _10736_ sky130_fd_sc_hd__inv_2
X_26679_ _09434_ _09689_ VGND VGND VPWR VPWR _09700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19220_ _04467_ _04507_ _04513_ _04515_ _04459_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__o221a_2
X_16432_ decode.regfile.registers_13\[29\] _10640_ _11187_ _12398_ _12399_ VGND VGND
+ VPWR VPWR _12400_ sky130_fd_sc_hd__a32o_1
X_28418_ clknet_leaf_38_clock _01431_ VGND VGND VPWR VPWR decode.immGen._imm_T_10\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13644_ memory.io_wb_reg_pc\[7\] _10001_ VGND VGND VPWR VPWR _10002_ sky130_fd_sc_hd__and2_1
XFILLER_0_224_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29398_ clknet_leaf_259_clock _02411_ VGND VGND VPWR VPWR decode.regfile.registers_4\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19151_ _04321_ _04021_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28349_ clknet_leaf_186_clock _01362_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_16363_ _12313_ _12332_ _11059_ _11149_ VGND VGND VPWR VPWR _12333_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_45_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13575_ memory.io_wb_memtoreg\[0\] VGND VGND VPWR VPWR _09940_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18102_ _03477_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ _11289_ _11306_ _11309_ VGND VGND VPWR VPWR _11310_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19082_ _04233_ _04209_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__nand2_1
X_16294_ _11079_ _11244_ _11080_ _12238_ _12265_ VGND VGND VPWR VPWR _12266_ sky130_fd_sc_hd__a41o_1
XFILLER_0_227_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18033_ decode.regfile.registers_15\[31\] _12667_ _12773_ _13011_ _03428_ VGND VGND
+ VPWR VPWR _03429_ sky130_fd_sc_hd__o311a_1
XFILLER_0_124_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15245_ _11062_ _11066_ _11076_ _11054_ VGND VGND VPWR VPWR _11242_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15176_ _10645_ _10654_ _10627_ _10659_ VGND VGND VPWR VPWR _11173_ sky130_fd_sc_hd__or4b_1
X_14127_ _10331_ VGND VGND VPWR VPWR _10332_ sky130_fd_sc_hd__clkbuf_4
X_19984_ net2735 _05217_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14058_ _09970_ _10288_ VGND VGND VPWR VPWR _10293_ sky130_fd_sc_hd__nand2_1
X_18935_ _04233_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__buf_4
XFILLER_0_207_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18866_ _04160_ _04164_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__or2_2
XFILLER_0_98_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17817_ _02986_ decode.regfile.registers_26\[25\] _13002_ _13484_ _02987_ VGND VGND
+ VPWR VPWR _03219_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18797_ _10045_ _10044_ _09942_ _10046_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_118_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_193_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17748_ decode.regfile.registers_13\[24\] _12534_ _12876_ _12664_ VGND VGND VPWR
+ VPWR _03151_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17679_ _03081_ _03082_ _03083_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19418_ _04623_ _04486_ _04247_ _04624_ _04268_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_194_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_194_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20690_ _05801_ _05808_ net1999 _05811_ _00693_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19349_ _04612_ _04621_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22360_ _06946_ _06951_ _06640_ _06954_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_116_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_198_Right_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21311_ _06165_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22291_ _06636_ _06881_ _06883_ _06885_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24030_ _08186_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__clkbuf_1
X_21242_ net835 _06119_ _06120_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold310 decode.regfile.registers_18\[10\] VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold321 execute.csr_write_data_out_reg\[28\] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold332 csr._mcycle_T_2\[0\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__buf_2
XFILLER_0_29_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold343 decode.regfile.registers_1\[27\] VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold354 csr._mcycle_T_3\[34\] VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__dlygate4sd3_1
X_21173_ _06074_ _06070_ net709 VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_132_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_132_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold365 decode.regfile.registers_30\[12\] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 decode.regfile.registers_13\[0\] VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 decode.regfile.registers_28\[7\] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__dlygate4sd3_1
X_20124_ decode.id_ex_imm_reg\[18\] decode.id_ex_pc_reg\[18\] VGND VGND VPWR VPWR
+ _05333_ sky130_fd_sc_hd__nand2_1
Xhold398 decode.regfile.registers_4\[8\] VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25981_ _09284_ VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_225_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27720_ clknet_leaf_16_clock _00749_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20055_ _00555_ _05228_ _05274_ _05231_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__o22a_1
X_24932_ _07199_ _08667_ _08668_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__nor3_1
XFILLER_0_102_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_1312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1010 fetch.bht.bhtTable_tag\[12\]\[7\] VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 fetch.bht.bhtTable_tag\[9\]\[3\] VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1032 fetch.bht.bhtTable_tag\[12\]\[21\] VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_147_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_147_clock
+ sky130_fd_sc_hd__clkbuf_8
X_27651_ clknet_leaf_48_clock net169 VGND VGND VPWR VPWR execute.io_reg_pc\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold1043 fetch.bht.bhtTable_target_pc\[4\]\[29\] VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__dlygate4sd3_1
X_24863_ _08619_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__clkbuf_1
Xhold1054 fetch.bht.bhtTable_target_pc\[5\]\[27\] VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1065 fetch.bht.bhtTable_tag\[8\]\[1\] VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 fetch.bht.bhtTable_target_pc\[5\]\[29\] VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26602_ _09432_ _09645_ VGND VGND VPWR VPWR _09656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23814_ _08063_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27582_ clknet_leaf_136_clock _00611_ VGND VGND VPWR VPWR csr.io_mem_pc\[23\] sky130_fd_sc_hd__dfxtp_4
Xhold1087 fetch.bht.bhtTable_tag\[6\]\[6\] VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1098 fetch.bht.bhtTable_target_pc\[7\]\[15\] VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__dlygate4sd3_1
X_24794_ _08583_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__clkbuf_1
X_29321_ clknet_leaf_226_clock _02334_ VGND VGND VPWR VPWR decode.regfile.registers_2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26533_ _09438_ _09577_ VGND VGND VPWR VPWR _09616_ sky130_fd_sc_hd__nand2_1
X_23745_ _06107_ net1248 _09907_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__mux2_1
X_20957_ net2505 _05915_ _05911_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29252_ clknet_leaf_232_clock _02265_ VGND VGND VPWR VPWR decode.regfile.registers_0\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_26464_ net333 _10195_ _10150_ _08903_ VGND VGND VPWR VPWR _09576_ sky130_fd_sc_hd__and4_1
XFILLER_0_83_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23676_ net812 csr.io_mem_pc\[29\] _07983_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20888_ _05858_ _05921_ net61 VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__and3_1
X_28203_ clknet_leaf_63_clock _01225_ VGND VGND VPWR VPWR csr.mscratch\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25415_ _10091_ VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__buf_4
XFILLER_0_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22627_ csr._minstret_T_3\[57\] csr._minstret_T_3\[56\] csr._minstret_T_3\[55\] _07190_
+ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__and4_1
X_29183_ clknet_leaf_162_clock _02196_ VGND VGND VPWR VPWR fetch.btb.btbTable\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26395_ net2388 _09534_ _09537_ _09525_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28134_ clknet_leaf_237_clock _01156_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25346_ _08905_ VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__clkbuf_4
X_22558_ csr._minstret_T_3\[36\] _07144_ net713 VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21509_ _06138_ net2246 _06263_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__mux2_1
X_28065_ clknet_leaf_188_clock _01087_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_40_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25277_ _08868_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_79_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22489_ _06637_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15030_ net437 _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__a31o_1
X_27016_ clknet_leaf_341_clock _00045_ VGND VGND VPWR VPWR decode.regfile.registers_22\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_24228_ _08288_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_185_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24159_ _08053_ net1797 _06274_ VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28967_ clknet_leaf_114_clock _01980_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_1311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16981_ decode.regfile.registers_6\[5\] _10602_ _12614_ _12939_ _12940_ VGND VGND
+ VPWR VPWR _12941_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_88_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18720_ _03726_ _04018_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_88_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27918_ clknet_leaf_66_clock _00947_ VGND VGND VPWR VPWR csr.io_csr_write_address\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_15932_ decode.regfile.registers_15\[16\] _11036_ _11204_ _11361_ VGND VGND VPWR
+ VPWR _11913_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_144_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28898_ clknet_leaf_135_clock _01911_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15863_ decode.regfile.registers_3\[14\] _11614_ _11367_ _11178_ VGND VGND VPWR VPWR
+ _11846_ sky130_fd_sc_hd__o2bb2a_1
X_18651_ execute.csr_read_data_out_reg\[20\] _03661_ _03660_ VGND VGND VPWR VPWR _03950_
+ sky130_fd_sc_hd__or3_1
X_27849_ clknet_leaf_325_clock _00878_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14814_ _10852_ _10855_ _10856_ VGND VGND VPWR VPWR _10857_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17602_ decode.regfile.registers_9\[20\] _12606_ _03007_ _03008_ VGND VGND VPWR VPWR
+ _03009_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_99_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15794_ _11047_ decode.regfile.registers_12\[12\] _10651_ _11053_ _10633_ VGND VGND
+ VPWR VPWR _11779_ sky130_fd_sc_hd__a2111o_1
X_18582_ _03708_ decode.id_ex_imm_reg\[23\] _03873_ _03880_ VGND VGND VPWR VPWR _03881_
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_188_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14745_ _10787_ _10767_ csr.io_mem_pc\[23\] VGND VGND VPWR VPWR _10788_ sky130_fd_sc_hd__a21oi_1
X_17533_ _10938_ _12542_ _12505_ decode.regfile.registers_23\[18\] _12714_ VGND VGND
+ VPWR VPWR _13480_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_47_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29519_ clknet_leaf_266_clock _02532_ VGND VGND VPWR VPWR decode.regfile.registers_8\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17464_ _13221_ _13410_ _13411_ _13412_ VGND VGND VPWR VPWR _13413_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_103_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14676_ _10703_ decode.id_ex_pc_reg\[0\] _10716_ execute.io_target_pc\[20\] _10718_
+ VGND VGND VPWR VPWR _10719_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19203_ _04008_ _03976_ _04497_ _04498_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__or4_1
X_16415_ _11446_ decode.regfile.registers_26\[29\] _11447_ _11348_ _10993_ VGND VGND
+ VPWR VPWR _12383_ sky130_fd_sc_hd__o2111a_1
X_13627_ _09986_ VGND VGND VPWR VPWR _09987_ sky130_fd_sc_hd__clkbuf_8
X_17395_ decode.regfile.registers_1\[15\] _12932_ _12933_ _10615_ _13344_ VGND VGND
+ VPWR VPWR _13345_ sky130_fd_sc_hd__o221a_1
XFILLER_0_229_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16346_ _11371_ decode.regfile.registers_0\[27\] VGND VGND VPWR VPWR _12316_ sky130_fd_sc_hd__nand2_1
X_19134_ _04250_ _04339_ _04277_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__mux2_1
X_13558_ csr.mtie csr.ie csr.mtip execute.exception_out_reg _09924_ VGND VGND VPWR
+ VPWR _09925_ sky130_fd_sc_hd__a311o_1
XFILLER_0_229_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19065_ net188 net189 _03988_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_915 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16277_ _12241_ _12248_ _11135_ VGND VGND VPWR VPWR _12249_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15228_ _10642_ VGND VGND VPWR VPWR _11225_ sky130_fd_sc_hd__buf_4
X_18016_ decode.regfile.registers_4\[31\] _12618_ _12620_ decode.regfile.registers_5\[31\]
+ _12737_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15159_ _11155_ VGND VGND VPWR VPWR _11156_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19967_ _03594_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_64_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_64_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18918_ _03835_ _03838_ _03821_ _03825_ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__o221a_1
XFILLER_0_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19898_ _03861_ _04618_ _04445_ _03865_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_220_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18849_ _03816_ _04147_ net353 VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21860_ net2483 _06497_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_79_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_79_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20811_ net122 _05879_ _05875_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21791_ _06037_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23530_ net2129 _07904_ _07901_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__or3b_1
XFILLER_0_33_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20742_ _05818_ decode.id_ex_rs1_data_reg\[28\] _03585_ VGND VGND VPWR VPWR _05842_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23461_ net9 _07861_ _07867_ _07865_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_150_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20673_ decode.id_ex_rs1_data_reg\[2\] decode.id_ex_ex_rs1_reg\[2\] _05056_ VGND
+ VGND VPWR VPWR _05799_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_189_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25200_ _10572_ net2442 _08828_ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__mux2_1
X_22412_ _06991_ _07006_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__or2b_1
XFILLER_0_163_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26180_ net2610 _09395_ _09405_ _09394_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23392_ _07089_ _07811_ _07812_ _07815_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_171_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25131_ _06149_ net1634 _08562_ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22343_ fetch.bht.bhtTable_tag\[12\]\[10\] fetch.bht.bhtTable_tag\[13\]\[10\] _06643_
+ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_17_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25062_ csr._mcycle_T_2\[25\] _08710_ _08754_ csr.mcycle\[25\] VGND VGND VPWR VPWR
+ _08755_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_227_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22274_ fetch.bht.bhtTable_tag\[8\]\[6\] fetch.bht.bhtTable_tag\[9\]\[6\] fetch.bht.bhtTable_tag\[10\]\[6\]
+ fetch.bht.bhtTable_tag\[11\]\[6\] _06645_ _06651_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_227_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24013_ net1433 execute.io_target_pc\[27\] _07960_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21225_ _10878_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold151 io_fetch_data[26] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
X_29870_ clknet_leaf_300_clock _02883_ VGND VGND VPWR VPWR decode.regfile.registers_19\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold162 fetch.bht.bhtTable_valid\[4\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_180_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold173 fetch.bht.bhtTable_valid\[5\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28821_ clknet_leaf_116_clock _01834_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_180_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold184 decode.regfile.registers_31\[17\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_180_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold195 fetch.btb.btbTable\[2\]\[0\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
X_21156_ _06062_ _06070_ net2748 VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20107_ _00563_ _05227_ _05318_ _05267_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__a2bb2oi_1
XTAP_TAPCELL_ROW_6_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28752_ clknet_leaf_121_clock _01765_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_21087_ _06030_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25964_ net2686 _09270_ _09275_ _09264_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20038_ _00553_ _05228_ _05259_ _05231_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__o22a_1
X_24915_ net524 _08656_ _08657_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__o21ba_1
X_27703_ clknet_leaf_19_clock _00732_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28683_ clknet_leaf_89_clock _01696_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_107_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25895_ net2105 _09226_ _09234_ _09235_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_30 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24846_ _06124_ net2077 _08607_ VGND VGND VPWR VPWR _08611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27634_ clknet_leaf_45_clock _00663_ VGND VGND VPWR VPWR execute.io_reg_pc\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_41 _08968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_52 _10041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_63 _10127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27565_ clknet_leaf_157_clock _00594_ VGND VGND VPWR VPWR csr.io_mem_pc\[6\] sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_74 _10240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24777_ _08070_ net1931 _08574_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__mux2_1
XINSDIODE1_85 _10594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21989_ net1950 _06588_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__or2_1
XFILLER_0_200_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_96 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_205_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14530_ _10573_ net2675 _10570_ VGND VGND VPWR VPWR _10574_ sky130_fd_sc_hd__mux2_1
X_29304_ clknet_leaf_242_clock _02317_ VGND VGND VPWR VPWR decode.regfile.registers_1\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_26516_ _09422_ _09602_ VGND VGND VPWR VPWR _09607_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23728_ _08015_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27496_ clknet_leaf_33_clock _00525_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29235_ clknet_leaf_172_clock _02248_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26447_ decode.regfile.registers_14\[23\] _09561_ _09565_ _09567_ VGND VGND VPWR
+ VPWR _02726_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_42_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _10048_ _10517_ VGND VGND VPWR VPWR _10525_ sky130_fd_sc_hd__nand2_1
X_23659_ net794 csr.io_mem_pc\[21\] _07972_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16200_ decode.regfile.registers_5\[23\] _10637_ _11139_ _11170_ VGND VGND VPWR VPWR
+ _12174_ sky130_fd_sc_hd__a31o_1
X_29166_ clknet_leaf_186_clock _02179_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_137_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17180_ _12496_ _13133_ _13134_ _13135_ VGND VGND VPWR VPWR _13136_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_137_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26378_ _09434_ _09515_ VGND VGND VPWR VPWR _09527_ sky130_fd_sc_hd__nand2_1
X_14392_ _10064_ _10474_ VGND VGND VPWR VPWR _10485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28117_ clknet_leaf_89_clock net2536 VGND VGND VPWR VPWR csr.minstret\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_141_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16131_ _12103_ _12105_ _12106_ VGND VGND VPWR VPWR _12107_ sky130_fd_sc_hd__o21ai_2
X_25329_ _08895_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29097_ clknet_leaf_70_clock _02110_ VGND VGND VPWR VPWR csr._mcycle_T_3\[45\] sky130_fd_sc_hd__dfxtp_1
X_28048_ clknet_leaf_235_clock _01070_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16062_ decode.regfile.registers_18\[19\] _10955_ _11113_ _11094_ _10976_ VGND VGND
+ VPWR VPWR _12040_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_224_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15013_ _11022_ VGND VGND VPWR VPWR _11023_ sky130_fd_sc_hd__clkbuf_4
X_19821_ _04338_ _05061_ _05092_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_209_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19752_ _03851_ _05026_ net212 VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__o21ai_1
X_16964_ decode.regfile.registers_20\[5\] _11024_ _12553_ _12823_ _12824_ VGND VGND
+ VPWR VPWR _12924_ sky130_fd_sc_hd__a41o_1
XFILLER_0_159_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18703_ net202 _04000_ _04001_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_155_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15915_ decode.regfile.registers_16\[15\] _11124_ _11878_ _11896_ VGND VGND VPWR
+ VPWR _11897_ sky130_fd_sc_hd__o22a_1
X_19683_ _04496_ _04955_ _04956_ _04960_ _04445_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__a311o_1
XFILLER_0_95_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16895_ decode.regfile.registers_19\[3\] _10599_ _10589_ _12518_ VGND VGND VPWR VPWR
+ _12857_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18634_ _03708_ decode.id_ex_imm_reg\[16\] _03932_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__a21oi_4
X_15846_ _11756_ decode.regfile.registers_28\[13\] _11067_ _11681_ _11440_ VGND VGND
+ VPWR VPWR _11830_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_95_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_201_Right_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18565_ _03863_ _03861_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15777_ _11571_ decode.regfile.registers_30\[12\] _11722_ _11723_ _11724_ VGND VGND
+ VPWR VPWR _11762_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_148_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17516_ _12645_ _13461_ _13462_ VGND VGND VPWR VPWR _13463_ sky130_fd_sc_hd__a21oi_1
X_14728_ csr.io_mem_pc\[28\] VGND VGND VPWR VPWR _10771_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18496_ net191 _03772_ _03775_ _03794_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_59_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14659_ decode.id_ex_pc_reg\[14\] VGND VGND VPWR VPWR _10702_ sky130_fd_sc_hd__inv_2
X_17447_ decode.regfile.registers_14\[16\] _10603_ _10618_ _12722_ VGND VGND VPWR
+ VPWR _13396_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17378_ decode.regfile.registers_20\[14\] _12770_ _13328_ _12537_ VGND VGND VPWR
+ VPWR _13329_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19117_ _04409_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16329_ decode.regfile.registers_22\[26\] _11096_ _12299_ VGND VGND VPWR VPWR _12300_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19048_ _04331_ _04344_ _04242_ _04346_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21010_ _05864_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_222_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_222_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22961_ _07097_ _07403_ _07405_ _07409_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_173_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24700_ _08062_ net2312 _08531_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21912_ csr.io_mret_vector\[22\] _10787_ _06539_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__mux2_1
X_25680_ _09110_ VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__buf_2
X_22892_ _06248_ VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24631_ _08498_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__clkbuf_1
X_21843_ _06499_ _06494_ _06495_ _06500_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27350_ clknet_leaf_46_clock _00379_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[23\]
+ sky130_fd_sc_hd__dfxtp_2
X_24562_ net1806 execute.io_target_pc\[3\] _08462_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__mux2_1
X_21774_ _06426_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_173_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26301_ net2448 _09475_ _09482_ _09471_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23513_ net96 _07889_ _07897_ _07893_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27281_ clknet_leaf_33_clock _00310_ VGND VGND VPWR VPWR decode.regfile.registers_31\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20725_ _05831_ _05808_ decode.id_ex_rs1_data_reg\[20\] _05832_ _00707_ VGND VGND
+ VPWR VPWR _00739_ sky130_fd_sc_hd__a32o_1
X_24493_ _08053_ net1585 _07276_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29020_ clknet_leaf_181_clock _02033_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26232_ _09441_ _09372_ VGND VGND VPWR VPWR _09442_ sky130_fd_sc_hd__nand2_1
X_23444_ decode.immGen._imm_T_10\[4\] _07847_ _05206_ VGND VGND VPWR VPWR _07857_
+ sky130_fd_sc_hd__or3b_1
X_20656_ csr.mcycle\[30\] _05588_ _05575_ csr.minstret\[30\] VGND VGND VPWR VPWR _05786_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26163_ _09263_ VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__buf_2
X_23375_ _07792_ _07796_ _07084_ _07799_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20587_ csr.minstret\[20\] _05574_ _05586_ csr.mcycle\[20\] VGND VGND VPWR VPWR _05727_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25114_ _08785_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22326_ fetch.bht.bhtTable_tag\[12\]\[8\] fetch.bht.bhtTable_tag\[13\]\[8\] fetch.bht.bhtTable_tag\[14\]\[8\]
+ fetch.bht.bhtTable_tag\[15\]\[8\] _06809_ _06649_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__mux4_2
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26094_ net1925 _09343_ _09350_ _09346_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25045_ _03554_ _08644_ _08743_ _06419_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__a211oi_1
X_29922_ clknet_5_5__leaf_clock _02935_ VGND VGND VPWR VPWR decode.regfile.registers_21\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22257_ _06650_ _06851_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21208_ decode.id_ex_ex_rd_reg\[2\] _05214_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__and2_1
X_29853_ clknet_leaf_306_clock _02866_ VGND VGND VPWR VPWR decode.regfile.registers_19\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22188_ _06633_ _06778_ _06780_ _06782_ _06642_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__o221ai_1
XTAP_TAPCELL_ROW_109_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28804_ clknet_leaf_131_clock _01817_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21139_ _06062_ _06058_ net2229 VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__and3_1
X_29784_ clknet_leaf_313_clock _02797_ VGND VGND VPWR VPWR decode.regfile.registers_16\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_26996_ clknet_leaf_334_clock _00025_ VGND VGND VPWR VPWR decode.regfile.registers_22\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_28735_ clknet_leaf_180_clock _01748_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13961_ _10122_ _10223_ VGND VGND VPWR VPWR _10235_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25947_ _08943_ _09253_ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15700_ _11435_ decode.regfile.registers_24\[10\] VGND VGND VPWR VPWR _11687_ sky130_fd_sc_hd__or2_1
X_16680_ _12644_ VGND VGND VPWR VPWR _12645_ sky130_fd_sc_hd__clkbuf_4
X_28666_ clknet_leaf_130_clock _01679_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_13892_ net2197 _10154_ _10193_ _10188_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__o211a_1
X_25878_ _09198_ VGND VGND VPWR VPWR _09226_ sky130_fd_sc_hd__buf_2
XFILLER_0_214_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24829_ _06107_ net1010 _08422_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27617_ clknet_leaf_151_clock _00646_ VGND VGND VPWR VPWR execute.io_target_pc\[26\]
+ sky130_fd_sc_hd__dfxtp_4
X_15631_ _11313_ decode.regfile.registers_4\[8\] _11191_ _10630_ _11462_ VGND VGND
+ VPWR VPWR _11620_ sky130_fd_sc_hd__a2111o_1
X_28597_ clknet_leaf_118_clock _01610_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_306 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_317 decode.regfile.registers_5\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15562_ _10650_ _10625_ _11053_ _11532_ _11552_ VGND VGND VPWR VPWR _11553_ sky130_fd_sc_hd__o32a_1
X_18350_ _03642_ decode.id_ex_ex_rs1_reg\[0\] _03646_ _03647_ _03648_ VGND VGND VPWR
+ VPWR _03649_ sky130_fd_sc_hd__o2111a_2
XTAP_TAPCELL_ROW_100_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_328 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27548_ clknet_leaf_41_clock _00577_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_139_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_339 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14513_ fetch.btb.btbTable\[4\]\[0\] fetch.btb.btbTable\[5\]\[0\] fetch.btb.btbTable\[6\]\[0\]
+ fetch.btb.btbTable\[7\]\[0\] _10556_ _10557_ VGND VGND VPWR VPWR _10558_ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17301_ _12759_ VGND VGND VPWR VPWR _13254_ sky130_fd_sc_hd__buf_2
XFILLER_0_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27479_ clknet_leaf_25_clock _00508_ VGND VGND VPWR VPWR decode.csr_read_reg sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15493_ _11235_ VGND VGND VPWR VPWR _11486_ sky130_fd_sc_hd__clkbuf_4
X_18281_ _03595_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__buf_2
XFILLER_0_194_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29218_ clknet_leaf_97_clock _02231_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17232_ _11022_ _12567_ _12586_ _12673_ decode.regfile.registers_16\[11\] VGND VGND
+ VPWR VPWR _13186_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_61_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _09999_ _10507_ VGND VGND VPWR VPWR _10515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17163_ _12667_ _12773_ _12670_ decode.regfile.registers_14\[9\] _13118_ VGND VGND
+ VPWR VPWR _13119_ sky130_fd_sc_hd__o221a_1
X_29149_ clknet_leaf_218_clock _02162_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14375_ net446 _10463_ _10475_ _10468_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16114_ _11679_ decode.regfile.registers_27\[20\] _11869_ VGND VGND VPWR VPWR _12091_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_52_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold909 fetch.bht.bhtTable_target_pc\[13\]\[27\] VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__dlygate4sd3_1
X_17094_ _12701_ decode.regfile.registers_28\[7\] _12698_ VGND VGND VPWR VPWR _13052_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16045_ _11300_ decode.regfile.registers_0\[19\] VGND VGND VPWR VPWR _12023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19804_ _03814_ _05076_ _05052_ net213 VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__o31a_1
XFILLER_0_209_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17996_ _12794_ _03391_ _03392_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__o21a_1
Xhold1609 decode.regfile.registers_10\[18\] VGND VGND VPWR VPWR net1836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19735_ _04546_ _04626_ _04924_ _04515_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__o311a_1
X_16947_ decode.regfile.registers_20\[4\] _12771_ _12905_ _12907_ _12538_ VGND VGND
+ VPWR VPWR _12908_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19666_ _04944_ _04896_ _04248_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16878_ decode.regfile.registers_4\[3\] _12548_ _12531_ decode.regfile.registers_5\[3\]
+ _12625_ VGND VGND VPWR VPWR _12840_ sky130_fd_sc_hd__a221o_1
XFILLER_0_172_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18617_ net109 _03665_ _03915_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15829_ _11547_ _11811_ _11812_ VGND VGND VPWR VPWR _11813_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19597_ _04878_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__buf_2
XFILLER_0_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18548_ _03709_ decode.id_ex_imm_reg\[24\] _03846_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_75_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18479_ execute.csr_read_data_out_reg\[29\] _03661_ _03660_ VGND VGND VPWR VPWR _03778_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_30_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20510_ csr.minstret\[10\] _05572_ _05582_ csr.mcycle\[10\] VGND VGND VPWR VPWR _05660_
+ sky130_fd_sc_hd__a22o_1
X_21490_ _06119_ net1289 _06252_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20441_ _05589_ _05590_ _05598_ _04459_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__o31a_1
XFILLER_0_132_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23160_ execute.io_target_pc\[15\] _06037_ _10970_ _03592_ VGND VGND VPWR VPWR _07598_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_28_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20372_ csr.io_csr_address\[4\] csr.io_csr_address\[5\] csr.io_csr_address\[6\] csr.io_csr_address\[8\]
+ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22111_ net275 VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23091_ _07368_ _07529_ _05246_ _07532_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_105_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22042_ _06636_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__buf_6
XFILLER_0_220_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26850_ _09377_ _09796_ VGND VGND VPWR VPWR _09800_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25801_ _09128_ VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__buf_2
X_26781_ _09383_ _09753_ VGND VGND VPWR VPWR _09760_ sky130_fd_sc_hd__nand2_1
X_23993_ net1022 execute.io_target_pc\[17\] _08164_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28520_ clknet_leaf_167_clock _01533_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25732_ net1948 _09139_ _09141_ _09142_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__o211a_1
X_22944_ net92 net89 VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_214_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28451_ clknet_leaf_147_clock _01464_ VGND VGND VPWR VPWR decode.io_id_pc\[9\] sky130_fd_sc_hd__dfxtp_1
X_25663_ _08962_ _09092_ VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__nand2_1
X_22875_ net1018 _10772_ _07324_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24614_ _08489_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27402_ clknet_leaf_28_clock _00431_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_28382_ clknet_leaf_184_clock _01395_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_21826_ _06479_ net512 _06396_ _06487_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25594_ _08968_ _09023_ VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__nand2_1
X_27333_ clknet_leaf_46_clock _00362_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24545_ _08105_ net1479 _09902_ VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21757_ _06441_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20708_ _05681_ _05684_ _05821_ _05804_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__o211a_1
X_27264_ clknet_leaf_0_clock _00293_ VGND VGND VPWR VPWR decode.regfile.registers_30\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_24476_ _08103_ net1464 _08411_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21688_ _06377_ _06390_ _06392_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_134_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29003_ clknet_leaf_94_clock _02016_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26215_ net192 VGND VGND VPWR VPWR _09430_ sky130_fd_sc_hd__buf_4
X_23427_ decode.control.io_opcode\[2\] _07847_ _05206_ VGND VGND VPWR VPWR _07848_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20639_ csr._minstret_T_3\[60\] _05616_ _05618_ csr._csr_read_data_T_8\[28\] _05770_
+ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27195_ clknet_leaf_360_clock _00224_ VGND VGND VPWR VPWR decode.regfile.registers_28\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire169 _00680_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14160_ _10053_ _10342_ VGND VGND VPWR VPWR _10351_ sky130_fd_sc_hd__nand2_1
X_26146_ _09381_ _09374_ VGND VGND VPWR VPWR _09382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23358_ net85 net220 _07740_ net86 VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22309_ fetch.bht.bhtTable_tag\[0\]\[0\] fetch.bht.bhtTable_tag\[1\]\[0\] _06706_
+ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14091_ _10069_ _10299_ VGND VGND VPWR VPWR _10311_ sky130_fd_sc_hd__nand2_1
X_26077_ _08922_ _09340_ VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__nand2_1
X_23289_ csr._csr_read_data_T_8\[22\] _07416_ csr.io_mret_vector\[22\] _07621_ _07719_
+ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25028_ net2789 _08712_ _08730_ csr.mcycle\[13\] csr.mcycle\[14\] VGND VGND VPWR
+ VPWR _08732_ sky130_fd_sc_hd__a221oi_1
X_29905_ clknet_leaf_340_clock _02918_ VGND VGND VPWR VPWR decode.regfile.registers_20\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_17850_ decode.regfile.registers_22\[26\] _12527_ _12687_ VGND VGND VPWR VPWR _03251_
+ sky130_fd_sc_hd__a21oi_1
X_29836_ clknet_leaf_298_clock _02849_ VGND VGND VPWR VPWR decode.regfile.registers_18\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16801_ _10931_ net604 _12487_ VGND VGND VPWR VPWR _12764_ sky130_fd_sc_hd__o21a_1
X_29767_ clknet_leaf_293_clock _02780_ VGND VGND VPWR VPWR decode.regfile.registers_16\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_17781_ _02997_ _12767_ _12965_ decode.regfile.registers_29\[24\] _03183_ VGND VGND
+ VPWR VPWR _03184_ sky130_fd_sc_hd__o221a_1
X_14993_ _10946_ _11004_ _11006_ _11007_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26979_ _10116_ _09862_ VGND VGND VPWR VPWR _09873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19520_ _04804_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__buf_1
XFILLER_0_195_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28718_ clknet_leaf_110_clock _01731_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_16732_ _10933_ _11012_ _11015_ _11026_ VGND VGND VPWR VPWR _12697_ sky130_fd_sc_hd__and4_2
XFILLER_0_117_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13944_ net2523 _10213_ _10225_ _10219_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_50_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29698_ clknet_leaf_291_clock _02711_ VGND VGND VPWR VPWR decode.regfile.registers_14\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19451_ _04664_ _04142_ _04177_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__o21ai_1
X_28649_ clknet_leaf_89_clock _01662_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16663_ _12627_ VGND VGND VPWR VPWR _12628_ sky130_fd_sc_hd__buf_4
X_13875_ net2106 _10180_ _10184_ _10175_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18402_ _03700_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__clkbuf_8
XINSDIODE1_103 _10771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15614_ _11436_ decode.regfile.registers_26\[7\] _11349_ _10980_ _11564_ VGND VGND
+ VPWR VPWR _11604_ sky130_fd_sc_hd__o2111a_1
XINSDIODE1_114 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19382_ _04254_ _04062_ _04487_ _04352_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16594_ _12558_ VGND VGND VPWR VPWR _12559_ sky130_fd_sc_hd__buf_4
XINSDIODE1_125 _11149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_136 _11896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_147 _12512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18333_ _03632_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__clkbuf_1
XINSDIODE1_158 _13085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15545_ decode.regfile.registers_5\[6\] _11313_ _11410_ VGND VGND VPWR VPWR _11536_
+ sky130_fd_sc_hd__or3_1
XINSDIODE1_169 decode.id_ex_rs1_data_reg\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18264_ _03594_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15476_ decode.regfile.registers_8\[4\] _11285_ _11365_ decode.regfile.registers_9\[4\]
+ _11132_ VGND VGND VPWR VPWR _11469_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17215_ _10604_ VGND VGND VPWR VPWR _13170_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14427_ _10373_ _10195_ _09933_ _10150_ VGND VGND VPWR VPWR _10504_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18195_ _10946_ _03532_ _03526_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__and3b_1
XFILLER_0_154_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17146_ decode.regfile.registers_2\[9\] _10608_ _12636_ _12639_ VGND VGND VPWR VPWR
+ _13102_ sky130_fd_sc_hd__a31o_1
X_14358_ _09964_ _10464_ VGND VGND VPWR VPWR _10466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold706 csr.minstret\[31\] VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold717 fetch.bht.bhtTable_tag\[11\]\[15\] VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold728 fetch.bht.bhtTable_target_pc\[8\]\[11\] VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17077_ decode.regfile.registers_17\[7\] _12901_ _12571_ _13034_ VGND VGND VPWR VPWR
+ _13035_ sky130_fd_sc_hd__a211o_1
Xhold739 fetch.bht.bhtTable_target_pc\[4\]\[25\] VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ _10130_ VGND VGND VPWR VPWR _10426_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16028_ decode.regfile.registers_20\[18\] _11452_ _11223_ _12006_ VGND VGND VPWR
+ VPWR _12007_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2107 execute.io_reg_pc\[26\] VGND VGND VPWR VPWR net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2118 decode.regfile.registers_8\[30\] VGND VGND VPWR VPWR net2345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2129 decode.regfile.registers_5\[20\] VGND VGND VPWR VPWR net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1406 fetch.bht.bhtTable_target_pc\[14\]\[25\] VGND VGND VPWR VPWR net1633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1417 fetch.bht.bhtTable_target_pc\[0\]\[20\] VGND VGND VPWR VPWR net1644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1428 fetch.bht.bhtTable_tag\[1\]\[10\] VGND VGND VPWR VPWR net1655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17979_ decode.regfile.registers_20\[30\] _12525_ _12552_ _12823_ _12824_ VGND VGND
+ VPWR VPWR _03376_ sky130_fd_sc_hd__a41o_1
XFILLER_0_137_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1439 decode.regfile.registers_11\[12\] VGND VGND VPWR VPWR net1666 sky130_fd_sc_hd__dlygate4sd3_1
X_19718_ _04973_ _04982_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20990_ _05978_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_196_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19649_ _04201_ _03938_ _04911_ _04860_ _04861_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__o2111ai_2
XTAP_TAPCELL_ROW_217_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22660_ net2775 _07210_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_213_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21611_ _10576_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__buf_4
XFILLER_0_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22591_ csr._minstret_T_3\[45\] csr._minstret_T_3\[44\] csr._minstret_T_3\[43\] _07166_
+ _07148_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__a41o_1
XFILLER_0_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24330_ _08341_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_1203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21542_ _06113_ net1722 _06284_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24261_ _08089_ net2175 _08300_ VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__mux2_1
X_21473_ _06253_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26000_ net2446 _09286_ _09296_ _09292_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__o211a_1
X_23212_ _07127_ _07640_ _07646_ _07367_ VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20424_ _05582_ _05551_ csr.mcycle\[1\] VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24192_ _08270_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23143_ net72 net225 net226 _07530_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__and4_2
X_20355_ _03741_ _03755_ _05517_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23074_ _07406_ _07510_ _07512_ _07097_ _07516_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__o311a_1
X_27951_ clknet_leaf_213_clock _00973_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_164_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20286_ _05464_ _05465_ _05411_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22025_ _00001_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__buf_4
X_26902_ _09430_ _09819_ VGND VGND VPWR VPWR _09829_ sky130_fd_sc_hd__nand2_1
X_27882_ clknet_leaf_25_clock _00911_ VGND VGND VPWR VPWR csr._mcycle_T_2\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29621_ clknet_leaf_280_clock _02634_ VGND VGND VPWR VPWR decode.regfile.registers_11\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_26833_ _09436_ _09751_ VGND VGND VPWR VPWR _09789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1940 decode.regfile.registers_9\[9\] VGND VGND VPWR VPWR net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1951 decode.io_id_pc\[11\] VGND VGND VPWR VPWR net2178 sky130_fd_sc_hd__dlygate4sd3_1
X_29552_ clknet_leaf_274_clock _02565_ VGND VGND VPWR VPWR decode.regfile.registers_9\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23976_ net1923 execute.io_target_pc\[9\] _08153_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__mux2_1
X_26764_ _09443_ _09708_ VGND VGND VPWR VPWR _09749_ sky130_fd_sc_hd__nand2_1
Xhold1962 fetch.bht.bhtTable_target_pc\[6\]\[4\] VGND VGND VPWR VPWR net2189 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1973 decode.io_id_pc\[12\] VGND VGND VPWR VPWR net2200 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1984 decode.io_id_pc\[19\] VGND VGND VPWR VPWR net2211 sky130_fd_sc_hd__dlygate4sd3_1
X_28503_ clknet_leaf_234_clock _01516_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_22927_ _07374_ _07376_ _07377_ _07122_ _06740_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__o221a_1
Xhold1995 decode.regfile.registers_19\[31\] VGND VGND VPWR VPWR net2222 sky130_fd_sc_hd__dlygate4sd3_1
X_25715_ net1149 _09125_ _09132_ _09129_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26695_ _10245_ _09710_ VGND VGND VPWR VPWR _09711_ sky130_fd_sc_hd__nand2_1
X_29483_ clknet_leaf_263_clock _02496_ VGND VGND VPWR VPWR decode.regfile.registers_7\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28434_ clknet_leaf_244_clock _01447_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_13660_ _10015_ _10016_ VGND VGND VPWR VPWR _10017_ sky130_fd_sc_hd__nand2_1
X_22858_ _07325_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__clkbuf_1
X_25646_ _09067_ VGND VGND VPWR VPWR _09092_ sky130_fd_sc_hd__buf_2
XFILLER_0_156_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21809_ csr._mcycle_T_2\[11\] _06467_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_26_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28365_ clknet_leaf_220_clock _01378_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_25577_ _08952_ _09049_ VGND VGND VPWR VPWR _09053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13591_ _09955_ VGND VGND VPWR VPWR _09956_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_195_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22789_ _07289_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15330_ decode.regfile.registers_19\[1\] _11048_ _11215_ _11216_ _11325_ VGND VGND
+ VPWR VPWR _11326_ sky130_fd_sc_hd__o41a_1
X_24528_ _08445_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27316_ clknet_leaf_42_clock _00345_ VGND VGND VPWR VPWR decode.id_ex_ex_rd_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28296_ clknet_leaf_164_clock _00016_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15261_ _10657_ _11065_ _11061_ _10662_ VGND VGND VPWR VPWR _11257_ sky130_fd_sc_hd__or4b_4
X_24459_ _08087_ net1747 _08400_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__mux2_1
X_27247_ clknet_leaf_32_clock _00276_ VGND VGND VPWR VPWR decode.regfile.registers_30\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17000_ _12695_ _12957_ _12958_ _12959_ VGND VGND VPWR VPWR _12960_ sky130_fd_sc_hd__a31o_1
X_14212_ net805 _10376_ _10381_ _10369_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_10_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27178_ clknet_leaf_362_clock _00207_ VGND VGND VPWR VPWR decode.regfile.registers_27\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_15192_ _11132_ _11177_ _11188_ VGND VGND VPWR VPWR _11189_ sky130_fd_sc_hd__a21o_1
XFILLER_0_227_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26129_ _09263_ VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__clkbuf_4
X_14143_ _10008_ _10333_ VGND VGND VPWR VPWR _10341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14074_ net837 _10287_ _10301_ _10291_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_56_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18951_ _04209_ _03911_ _03989_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17902_ _12765_ net635 _13492_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__o21a_1
X_18882_ net335 _03701_ _03689_ decode.id_ex_rs1_data_reg\[14\] _04080_ VGND VGND
+ VPWR VPWR _04181_ sky130_fd_sc_hd__o221a_2
XFILLER_0_197_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17833_ decode.regfile.registers_2\[26\] _12835_ _12836_ _03233_ VGND VGND VPWR VPWR
+ _03234_ sky130_fd_sc_hd__a211o_1
X_29819_ clknet_leaf_315_clock _02832_ VGND VGND VPWR VPWR decode.regfile.registers_18\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17764_ decode.regfile.registers_15\[24\] _12667_ _12773_ _13011_ VGND VGND VPWR
+ VPWR _03167_ sky130_fd_sc_hd__o31a_1
XFILLER_0_221_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14976_ _10948_ _10954_ _10997_ net437 _10999_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__o311a_1
XFILLER_0_107_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19503_ _04786_ _04787_ net350 _04444_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__a31o_1
X_16715_ decode.regfile.registers_18\[0\] _12566_ _12573_ _12676_ _12679_ VGND VGND
+ VPWR VPWR _12680_ sky130_fd_sc_hd__o221a_1
X_13927_ _10042_ _10210_ VGND VGND VPWR VPWR _10216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17695_ _11014_ _13168_ decode.regfile.registers_23\[22\] _12995_ VGND VGND VPWR
+ VPWR _03100_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19434_ _04160_ _04164_ _04721_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_179_Right_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16646_ _12610_ VGND VGND VPWR VPWR _12611_ sky130_fd_sc_hd__clkbuf_4
X_13858_ _10131_ VGND VGND VPWR VPWR _10175_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_191_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19365_ _03972_ _03974_ _04007_ _04655_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16577_ _12541_ VGND VGND VPWR VPWR _12542_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_191_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13789_ memory.io_wb_reg_pc\[28\] _09946_ _09947_ _10125_ VGND VGND VPWR VPWR _10126_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18316_ _03623_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__clkbuf_1
X_15528_ decode.regfile.registers_21\[5\] _11060_ _11098_ _11227_ _11519_ VGND VGND
+ VPWR VPWR _11520_ sky130_fd_sc_hd__o311a_1
Xclkbuf_2_3_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_3_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19296_ net219 VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__buf_4
XFILLER_0_31_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18247_ _10910_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15459_ _11103_ VGND VGND VPWR VPWR _11452_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18178_ _10579_ decode.control.io_opcode\[5\] decode.control.io_opcode\[4\] _10580_
+ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__nand4_2
Xmax_cap200 _10101_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_4
XFILLER_0_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap211 _09963_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_4
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold503 decode.regfile.registers_8\[8\] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17129_ _12915_ decode.regfile.registers_25\[8\] _13045_ _12812_ VGND VGND VPWR VPWR
+ _13086_ sky130_fd_sc_hd__or4_1
Xhold514 decode.regfile.registers_30\[23\] VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 fetch.bht.bhtTable_target_pc\[1\]\[7\] VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold536 decode.regfile.registers_1\[8\] VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold547 decode.regfile.registers_28\[24\] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold558 fetch.bht.bhtTable_target_pc\[2\]\[11\] VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__dlygate4sd3_1
X_20140_ _05333_ _05346_ _05339_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__nand3_1
XFILLER_0_111_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold569 decode.regfile.registers_12\[10\] VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20071_ _00558_ _05228_ _05287_ _05231_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1203 fetch.bht.bhtTable_target_pc\[11\]\[14\] VGND VGND VPWR VPWR net1430 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 fetch.bht.bhtTable_target_pc\[12\]\[31\] VGND VGND VPWR VPWR net1441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 fetch.bht.bhtTable_target_pc\[5\]\[8\] VGND VGND VPWR VPWR net1452 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23830_ execute.io_target_pc\[12\] VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__buf_2
XFILLER_0_139_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1236 decode.regfile.registers_18\[14\] VGND VGND VPWR VPWR net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 fetch.bht.bhtTable_tag\[12\]\[1\] VGND VGND VPWR VPWR net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 fetch.bht.bhtTable_tag\[9\]\[13\] VGND VGND VPWR VPWR net1485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1269 fetch.bht.bhtTable_target_pc\[0\]\[2\] VGND VGND VPWR VPWR net1496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23761_ _08032_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__clkbuf_1
X_20973_ execute.io_reg_pc\[12\] _05965_ _05961_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__and3_1
XFILLER_0_174_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22712_ csr._mcycle_T_2\[30\] _07236_ VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__or2_1
X_25500_ _08978_ VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__clkbuf_4
X_26480_ net2253 _09578_ _09586_ _09582_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23692_ _07996_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25431_ _08964_ _08946_ VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_157_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22643_ _07199_ _07204_ _07205_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__nor3_1
XFILLER_0_220_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_362_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_362_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28150_ clknet_leaf_190_clock _01172_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_25362_ _08916_ _08907_ VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22574_ csr._minstret_T_3\[33\] csr.minstret\[30\] csr.minstret\[31\] _07151_ VGND
+ VGND VPWR VPWR _07158_ sky130_fd_sc_hd__and4_1
XFILLER_0_146_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24313_ _08332_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27101_ clknet_leaf_357_clock _00130_ VGND VGND VPWR VPWR decode.regfile.registers_25\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21525_ _06280_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__clkbuf_1
X_28081_ clknet_leaf_210_clock _01103_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25293_ _08869_ net2728 VGND VGND VPWR VPWR _08877_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27032_ clknet_leaf_332_clock _00061_ VGND VGND VPWR VPWR decode.regfile.registers_23\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24244_ _08072_ net1621 _08289_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21456_ _06147_ net1858 _06241_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20407_ csr.minstret\[0\] _05560_ _05566_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__a21o_1
X_24175_ _08261_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21387_ _06206_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_187_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23126_ _07557_ _07559_ _07097_ _07565_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_112_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20338_ _10790_ decode.id_ex_pc_reg\[26\] _10854_ _05494_ decode.id_ex_pc_reg\[28\]
+ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__a41o_1
X_28983_ clknet_leaf_125_clock _01996_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_300_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_300_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_183_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput67 net67 VGND VGND VPWR VPWR io_fetch_address[0] sky130_fd_sc_hd__clkbuf_4
X_27934_ clknet_leaf_165_clock _00005_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_23057_ execute.io_target_pc\[9\] _07346_ _07488_ _07500_ _07348_ VGND VGND VPWR
+ VPWR _07501_ sky130_fd_sc_hd__a2111o_1
Xoutput78 net78 VGND VGND VPWR VPWR io_fetch_address[1] sky130_fd_sc_hd__clkbuf_4
X_20269_ _05451_ _05452_ _05420_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__o21ai_1
Xoutput89 net89 VGND VGND VPWR VPWR io_fetch_address[2] sky130_fd_sc_hd__clkbuf_4
X_22008_ net2014 _06601_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_125_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27865_ clknet_leaf_317_clock _00894_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2460 execute.io_reg_pc\[3\] VGND VGND VPWR VPWR net2687 sky130_fd_sc_hd__dlygate4sd3_1
X_29604_ clknet_leaf_276_clock _02617_ VGND VGND VPWR VPWR decode.regfile.registers_11\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14830_ _10871_ _10872_ _10807_ _10763_ _10868_ VGND VGND VPWR VPWR _10873_ sky130_fd_sc_hd__a41o_1
Xhold2471 decode.regfile.registers_0\[27\] VGND VGND VPWR VPWR net2698 sky130_fd_sc_hd__dlygate4sd3_1
X_26816_ _09420_ _09776_ VGND VGND VPWR VPWR _09780_ sky130_fd_sc_hd__nand2_1
Xhold2482 decode.regfile.registers_14\[25\] VGND VGND VPWR VPWR net2709 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_315_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_315_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_208_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2493 decode.regfile.registers_13\[16\] VGND VGND VPWR VPWR net2720 sky130_fd_sc_hd__dlygate4sd3_1
X_27796_ clknet_leaf_305_clock _00825_ VGND VGND VPWR VPWR memory.io_wb_readdata\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1770 decode.regfile.registers_20\[19\] VGND VGND VPWR VPWR net1997 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29535_ clknet_leaf_312_clock _02548_ VGND VGND VPWR VPWR decode.regfile.registers_9\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ csr.io_mem_pc\[16\] _10764_ VGND VGND VPWR VPWR _10804_ sky130_fd_sc_hd__nand2_1
X_26747_ _09426_ _09733_ VGND VGND VPWR VPWR _09740_ sky130_fd_sc_hd__nand2_1
Xhold1781 decode.regfile.registers_20\[0\] VGND VGND VPWR VPWR net2008 sky130_fd_sc_hd__dlygate4sd3_1
X_23959_ net2029 execute.io_target_pc\[1\] _07983_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1792 csr.mscratch\[7\] VGND VGND VPWR VPWR net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16500_ decode.regfile.registers_8\[31\] _11284_ _11287_ decode.regfile.registers_9\[31\]
+ VGND VGND VPWR VPWR _12466_ sky130_fd_sc_hd__o22a_1
X_13712_ _10060_ _10021_ memory.io_wb_readdata\[16\] VGND VGND VPWR VPWR _10061_ sky130_fd_sc_hd__and3b_1
X_14692_ _10731_ execute.io_target_pc\[7\] decode.id_ex_pc_reg\[21\] _10717_ _10734_
+ VGND VGND VPWR VPWR _10735_ sky130_fd_sc_hd__o221a_1
X_29466_ clknet_leaf_250_clock _02479_ VGND VGND VPWR VPWR decode.regfile.registers_7\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_17480_ _13421_ _13427_ _12726_ VGND VGND VPWR VPWR _13428_ sky130_fd_sc_hd__nand3b_1
X_26678_ net2311 _09692_ _09699_ _09688_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28417_ clknet_leaf_39_clock _01430_ VGND VGND VPWR VPWR decode.immGen._imm_T_10\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16431_ _11047_ decode.regfile.registers_12\[29\] _10650_ _11053_ _10632_ VGND VGND
+ VPWR VPWR _12399_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25629_ _08929_ _09079_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__nand2_1
X_13643_ _09978_ VGND VGND VPWR VPWR _10001_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29397_ clknet_leaf_258_clock _02410_ VGND VGND VPWR VPWR decode.regfile.registers_4\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19150_ _04443_ _04273_ _04446_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__o21ai_1
X_28348_ clknet_leaf_201_clock _01361_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_16362_ _12329_ _12330_ _12331_ _11356_ VGND VGND VPWR VPWR _12332_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_45_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13574_ memory.io_wb_memtoreg\[1\] VGND VGND VPWR VPWR _09939_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_45_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18101_ _03469_ _03467_ _03474_ decode.io_id_pc\[8\] VGND VGND VPWR VPWR _03477_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15313_ decode.regfile.registers_7\[1\] _11308_ _11169_ decode.regfile.registers_6\[1\]
+ _11165_ VGND VGND VPWR VPWR _11309_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_147_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16293_ decode.regfile.registers_23\[25\] _11262_ _11089_ _11493_ _12264_ VGND VGND
+ VPWR VPWR _12265_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19081_ net286 _04181_ _04233_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__mux2_1
X_28279_ clknet_leaf_85_clock net2631 VGND VGND VPWR VPWR csr._csr_read_data_T_8\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18032_ _12670_ _03426_ _03427_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15244_ _11064_ net532 _11068_ _11240_ VGND VGND VPWR VPWR _11241_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15175_ _11136_ _11163_ _11166_ _11171_ VGND VGND VPWR VPWR _11172_ sky130_fd_sc_hd__a211o_1
X_14126_ _10330_ VGND VGND VPWR VPWR _10331_ sky130_fd_sc_hd__clkbuf_4
X_19983_ net408 _05217_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__nor2_1
X_14057_ net1295 _10287_ _10292_ _10291_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__o211a_1
X_18934_ _03988_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_185_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18865_ _03707_ decode.id_ex_imm_reg\[10\] _04161_ _04163_ VGND VGND VPWR VPWR _04164_
+ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_201_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17816_ _13407_ decode.regfile.registers_25\[25\] _13482_ _12811_ VGND VGND VPWR
+ VPWR _03218_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18796_ _04091_ _04094_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__xor2_4
XFILLER_0_221_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17747_ _11022_ _12568_ _12535_ _12674_ decode.regfile.registers_16\[24\] VGND VGND
+ VPWR VPWR _03150_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_193_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14959_ _10985_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17678_ decode.regfile.registers_7\[22\] _12882_ _13020_ _12622_ decode.regfile.registers_6\[22\]
+ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__a32o_1
XFILLER_0_159_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19417_ _04671_ _04704_ _04277_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16629_ _12593_ VGND VGND VPWR VPWR _12594_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19348_ _04130_ _04131_ _04637_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__or3_1
XFILLER_0_190_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19279_ _04280_ _04282_ _04368_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__or3b_2
XFILLER_0_116_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21310_ net980 _10871_ _06157_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22290_ _06687_ _06884_ _06641_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21241_ _09910_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__clkbuf_8
Xhold300 _01245_ VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold311 decode.regfile.registers_12\[5\] VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold322 decode.regfile.registers_13\[6\] VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold333 _01184_ VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold344 decode.regfile.registers_6\[10\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
X_21172_ _06080_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__clkbuf_1
Xhold355 decode.regfile.registers_31\[5\] VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__buf_1
XFILLER_0_229_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold366 decode.regfile.registers_7\[8\] VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold377 decode.regfile.registers_30\[2\] VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20123_ decode.id_ex_imm_reg\[18\] decode.id_ex_pc_reg\[18\] VGND VGND VPWR VPWR
+ _05332_ sky130_fd_sc_hd__nor2_1
Xhold388 decode.regfile.registers_19\[3\] VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 execute.csr_write_data_out_reg\[1\] VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25980_ _09930_ _10194_ _10240_ _08902_ VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_225_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_215_Right_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20054_ _05272_ _05273_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__nor2_1
X_24931_ csr._mcycle_T_3\[45\] csr._mcycle_T_3\[44\] csr._mcycle_T_3\[43\] _08662_
+ VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__and4_2
Xhold1000 fetch.bht.bhtTable_tag\[1\]\[12\] VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_0_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1011 fetch.bht.bhtTable_target_pc\[10\]\[7\] VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1022 fetch.bht.bhtTable_target_pc\[4\]\[10\] VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_37_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27650_ clknet_leaf_47_clock _00679_ VGND VGND VPWR VPWR execute.io_reg_pc\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1033 decode.regfile.registers_21\[18\] VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24862_ _06140_ net1021 _08388_ VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__mux2_1
Xhold1044 decode.regfile.registers_15\[30\] VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1055 fetch.bht.bhtTable_target_pc\[2\]\[6\] VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 fetch.bht.bhtTable_target_pc\[0\]\[27\] VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__dlygate4sd3_1
X_26601_ net2731 _09649_ _09655_ _09648_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__o211a_1
X_23813_ _08062_ net2614 _08058_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_159_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 decode.regfile.registers_15\[28\] VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24793_ _08087_ net2064 _08574_ VGND VGND VPWR VPWR _08583_ sky130_fd_sc_hd__mux2_1
X_27581_ clknet_leaf_171_clock _00610_ VGND VGND VPWR VPWR csr.io_mem_pc\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_1_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1088 decode.regfile.registers_5\[18\] VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1099 fetch.bht.bhtTable_tag\[3\]\[24\] VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29320_ clknet_leaf_228_clock _02333_ VGND VGND VPWR VPWR decode.regfile.registers_2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23744_ _08023_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__clkbuf_1
X_26532_ net1304 _09605_ _09615_ _09608_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20956_ _05959_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29251_ clknet_leaf_232_clock _02264_ VGND VGND VPWR VPWR decode.regfile.registers_0\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_23675_ _07986_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26463_ net1419 _09535_ _09575_ _09567_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20887_ _05922_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28202_ clknet_leaf_62_clock net1570 VGND VGND VPWR VPWR csr.mscratch\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22626_ csr._minstret_T_3\[56\] csr._minstret_T_3\[55\] _07190_ net1764 VGND VGND
+ VPWR VPWR _07194_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_165_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25414_ net574 _08951_ _08953_ _08950_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29182_ clknet_leaf_163_clock _02195_ VGND VGND VPWR VPWR fetch.btb.btbTable\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26394_ _09450_ _09535_ VGND VGND VPWR VPWR _09537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28133_ clknet_leaf_235_clock _01155_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_25345_ _08904_ VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__buf_2
XFILLER_0_118_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22557_ net2673 _07144_ _07145_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__o21a_1
XFILLER_0_180_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21508_ _06271_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28064_ clknet_leaf_190_clock _01086_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_25276_ _05856_ decode.regfile.registers_0\[0\] VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22488_ _07078_ _07079_ _07082_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24227_ _08055_ net1432 _06241_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27015_ clknet_leaf_342_clock _00044_ VGND VGND VPWR VPWR decode.regfile.registers_22\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_21439_ _06130_ net2025 _06230_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24158_ _08252_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23109_ net226 _07530_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__nand2_1
X_28966_ clknet_leaf_97_clock _01979_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_24089_ net1410 execute.io_target_pc\[0\] _06450_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__mux2_1
X_16980_ decode.regfile.registers_4\[5\] _12617_ _12619_ decode.regfile.registers_5\[5\]
+ _12622_ VGND VGND VPWR VPWR _12940_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_1323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27917_ clknet_leaf_66_clock _00946_ VGND VGND VPWR VPWR csr.io_csr_write_address\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_15931_ _10957_ decode.regfile.registers_22\[16\] _11450_ _10978_ _10990_ VGND VGND
+ VPWR VPWR _11912_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_55_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28897_ clknet_leaf_170_clock _01910_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_254_clock clknet_5_22__leaf_clock VGND VGND VPWR VPWR clknet_leaf_254_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _10086_ _03785_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__nand2_1
X_15862_ decode.regfile.registers_2\[14\] _11369_ _11152_ _11844_ VGND VGND VPWR VPWR
+ _11845_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27848_ clknet_leaf_324_clock _00877_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2290 csr.mscratch\[6\] VGND VGND VPWR VPWR net2517 sky130_fd_sc_hd__dlygate4sd3_1
X_17601_ _11017_ _12502_ _12509_ decode.regfile.registers_8\[20\] _12725_ VGND VGND
+ VPWR VPWR _03008_ sky130_fd_sc_hd__o32a_1
XFILLER_0_189_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14813_ _10772_ _10773_ _10774_ _10853_ decode.id_ex_pc_reg\[27\] VGND VGND VPWR
+ VPWR _10856_ sky130_fd_sc_hd__a311o_1
X_18581_ _03879_ _03759_ _10101_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__and3_1
X_15793_ _11765_ _11776_ _11777_ VGND VGND VPWR VPWR _11778_ sky130_fd_sc_hd__o21ai_1
X_27779_ clknet_leaf_35_clock _00808_ VGND VGND VPWR VPWR memory.io_wb_readdata\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17532_ decode.regfile.registers_22\[18\] _12528_ _13478_ _12687_ VGND VGND VPWR
+ VPWR _13479_ sky130_fd_sc_hd__a211o_1
X_29518_ clknet_leaf_266_clock _02531_ VGND VGND VPWR VPWR decode.regfile.registers_8\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14744_ csr.io_mem_pc\[22\] VGND VGND VPWR VPWR _10787_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_269_clock clknet_5_22__leaf_clock VGND VGND VPWR VPWR clknet_leaf_269_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17463_ _13215_ decode.regfile.registers_28\[16\] _13093_ VGND VGND VPWR VPWR _13412_
+ sky130_fd_sc_hd__o21a_1
X_29449_ clknet_leaf_262_clock _02462_ VGND VGND VPWR VPWR decode.regfile.registers_6\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14675_ _10690_ execute.io_target_pc\[4\] decode.id_ex_pc_reg\[21\] _10717_ VGND
+ VGND VPWR VPWR _10718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19202_ _04022_ _04023_ _04389_ _04398_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_0_104_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16414_ _11346_ decode.regfile.registers_30\[29\] _12095_ _12096_ _12097_ VGND VGND
+ VPWR VPWR _12382_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_7_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13626_ _09942_ VGND VGND VPWR VPWR _09986_ sky130_fd_sc_hd__buf_4
X_17394_ _12934_ _12616_ _12558_ decode.regfile.registers_0\[15\] VGND VGND VPWR VPWR
+ _13344_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19133_ _04045_ _04054_ _03971_ _04321_ _04307_ _04325_ VGND VGND VPWR VPWR _04430_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16345_ decode.regfile.registers_1\[27\] VGND VGND VPWR VPWR _12315_ sky130_fd_sc_hd__inv_2
X_13557_ csr.msie csr.msip csr.ie _09923_ VGND VGND VPWR VPWR _09924_ sky130_fd_sc_hd__a31o_1
XFILLER_0_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19064_ _04306_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16276_ _12245_ _12246_ _12247_ VGND VGND VPWR VPWR _12248_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18015_ _10616_ decode.regfile.registers_6\[31\] VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__and2b_1
XFILLER_0_129_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15227_ decode.regfile.registers_20\[0\] _11103_ _11214_ _11220_ _11223_ VGND VGND
+ VPWR VPWR _11224_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_207_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_207_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15158_ decode.immGen._imm_T_24\[1\] _11107_ _11041_ _11055_ VGND VGND VPWR VPWR
+ _11155_ sky130_fd_sc_hd__and4_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14109_ net2491 _10315_ _10321_ _10317_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__o211a_1
X_19966_ _05213_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15089_ _11060_ _11065_ _11049_ _11085_ VGND VGND VPWR VPWR _11086_ sky130_fd_sc_hd__or4_2
XFILLER_0_61_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18917_ _03835_ _03838_ _03844_ _03847_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__a211o_1
XFILLER_0_226_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19897_ _05160_ _05161_ _05165_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_207_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18848_ net102 _03664_ _04146_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_220_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clock clock VGND VGND VPWR VPWR clknet_0_clock sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_220_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18779_ _03658_ execute.csr_read_data_out_reg\[14\] execute.io_reg_pc\[14\] _03776_
+ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20810_ _05880_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21790_ _06457_ net217 _06458_ _06459_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__nand4b_2
XTAP_TAPCELL_ROW_19_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20741_ _05831_ _05813_ decode.id_ex_rs1_data_reg\[27\] _05841_ _00714_ VGND VGND
+ VPWR VPWR _00746_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23460_ _11012_ _07862_ _07859_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__or3b_1
X_20672_ _03585_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__buf_2
XFILLER_0_190_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22411_ net86 _07005_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__xor2_1
XFILLER_0_147_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23391_ _07064_ _07813_ _07814_ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__and3_1
XFILLER_0_174_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25130_ _08793_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__clkbuf_1
X_22342_ fetch.bht.bhtTable_tag\[8\]\[10\] fetch.bht.bhtTable_tag\[9\]\[10\] fetch.bht.bhtTable_tag\[10\]\[10\]
+ fetch.bht.bhtTable_tag\[11\]\[10\] _06878_ _06621_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__mux4_1
XFILLER_0_169_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25061_ _03555_ csr.mcycle\[24\] csr.mcycle\[23\] _08748_ VGND VGND VPWR VPWR _08754_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22273_ _06867_ _06623_ _06687_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_227_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24012_ _08177_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21224_ _06108_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold152 io_fetch_data[28] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 fetch.bht.bhtTable_valid\[0\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28820_ clknet_leaf_118_clock _01833_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_180_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold174 fetch.bht.bhtTable_valid\[15\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold185 fetch.btb.btbTable\[15\]\[0\] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21155_ _06071_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_180_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold196 fetch.btb.btbTable\[3\]\[0\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20106_ _05316_ _05317_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_6_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28751_ clknet_leaf_110_clock _01764_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25963_ _08960_ _09267_ VGND VGND VPWR VPWR _09275_ sky130_fd_sc_hd__nand2_1
X_21086_ execute.csr_read_data_out_reg\[31\] _06025_ _03583_ VGND VGND VPWR VPWR _06030_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27702_ clknet_leaf_20_clock _00731_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_20037_ _05257_ _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__nor2_1
X_24914_ csr._mcycle_T_3\[39\] csr._mcycle_T_3\[38\] _08654_ _06422_ VGND VGND VPWR
+ VPWR _08657_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28682_ clknet_leaf_96_clock _01695_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25894_ _09128_ VGND VGND VPWR VPWR _09235_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27633_ clknet_leaf_44_clock _00662_ VGND VGND VPWR VPWR execute.io_reg_pc\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_24845_ _08610_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__clkbuf_1
XINSDIODE1_20 _02984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_31 _08929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_198_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_42 _09392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_53 _10073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27564_ clknet_leaf_162_clock _00593_ VGND VGND VPWR VPWR csr.io_mem_pc\[5\] sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_64 _10127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24776_ _08562_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__clkbuf_8
X_21988_ csr._mcycle_T_2\[17\] _06587_ _06597_ _06592_ VGND VGND VPWR VPWR _01237_
+ sky130_fd_sc_hd__o211a_1
XINSDIODE1_75 _10240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_86 _10594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29303_ clknet_leaf_242_clock _02316_ VGND VGND VPWR VPWR decode.regfile.registers_1\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_97 _10610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_969 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26515_ net1994 _09605_ _09606_ _09595_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__o211a_1
X_23727_ net1624 _10760_ _08014_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__mux2_1
X_20939_ _05949_ _05945_ net54 VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27495_ clknet_leaf_30_clock _00524_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29234_ clknet_leaf_129_clock _02247_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_26446_ _09566_ VGND VGND VPWR VPWR _09567_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_42_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ net427 _10520_ _10524_ _10522_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__o211a_1
X_23658_ _07977_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29165_ clknet_leaf_202_clock _02178_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_22609_ csr._minstret_T_3\[50\] csr._minstret_T_3\[49\] _07178_ net1258 VGND VGND
+ VPWR VPWR _07183_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_10_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14391_ net678 _10477_ _10484_ _10481_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23589_ _07939_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26377_ net2223 _09518_ _09526_ _09525_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_137_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28116_ clknet_leaf_89_clock _01138_ VGND VGND VPWR VPWR csr.minstret\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_153_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16130_ decode.regfile.registers_3\[21\] _11614_ _11410_ _10636_ VGND VGND VPWR VPWR
+ _12106_ sky130_fd_sc_hd__o2bb2a_1
X_25328_ _08891_ net2695 VGND VGND VPWR VPWR _08895_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29096_ clknet_leaf_71_clock _02109_ VGND VGND VPWR VPWR csr._mcycle_T_3\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28047_ clknet_leaf_222_clock _01069_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16061_ decode.regfile.registers_17\[19\] _10988_ _11113_ _11119_ _12038_ VGND VGND
+ VPWR VPWR _12039_ sky130_fd_sc_hd__a41o_1
X_25259_ _08859_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15012_ _11021_ VGND VGND VPWR VPWR _11022_ sky130_fd_sc_hd__buf_2
XFILLER_0_110_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19820_ _04297_ _04261_ _04263_ _05091_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_193_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_193_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_166_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19751_ _04840_ _04212_ _04196_ _05025_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__a31o_4
X_28949_ clknet_leaf_141_clock _01962_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_16963_ _10931_ decode.regfile.registers_30\[5\] _12487_ VGND VGND VPWR VPWR _12923_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18702_ _03968_ _03995_ _03654_ _03649_ decode.id_ex_islui_reg VGND VGND VPWR VPWR
+ _04001_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_159_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15914_ _11879_ _11895_ _11054_ _11318_ VGND VGND VPWR VPWR _11896_ sky130_fd_sc_hd__o2bb2a_1
X_19682_ _04957_ _04959_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__nor2_1
X_16894_ decode.regfile.registers_18\[3\] _12826_ _12827_ _12855_ VGND VGND VPWR VPWR
+ _12856_ sky130_fd_sc_hd__o22a_1
XFILLER_0_200_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_1254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18633_ _10063_ _03785_ _03931_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__a21oi_2
X_15845_ _11679_ decode.regfile.registers_27\[13\] _11258_ VGND VGND VPWR VPWR _11829_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_95_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18564_ decode.id_ex_rs1_data_reg\[30\] _03817_ _03698_ _03858_ VGND VGND VPWR VPWR
+ _03863_ sky130_fd_sc_hd__o31a_4
X_15776_ _11243_ VGND VGND VPWR VPWR _11761_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17515_ decode.regfile.registers_7\[18\] _12645_ _12726_ VGND VGND VPWR VPWR _13462_
+ sky130_fd_sc_hd__o21ai_1
X_14727_ _10759_ csr.io_mem_pc\[28\] csr.io_mem_pc\[29\] _10769_ VGND VGND VPWR VPWR
+ _10770_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18495_ _03656_ _03793_ decode.id_ex_rs1_data_reg\[28\] _03689_ VGND VGND VPWR VPWR
+ _03794_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_131_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_131_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17446_ decode.regfile.registers_13\[16\] _12774_ _13393_ _13394_ _12662_ VGND VGND
+ VPWR VPWR _13395_ sky130_fd_sc_hd__a221o_1
X_14658_ decode.id_ex_pc_reg\[27\] _10687_ _10691_ _10700_ VGND VGND VPWR VPWR _10701_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13609_ net2490 _09938_ _09971_ _09957_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17377_ decode.regfile.registers_19\[14\] _12677_ _13306_ _13327_ _12543_ VGND VGND
+ VPWR VPWR _13328_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14589_ _10631_ VGND VGND VPWR VPWR _10632_ sky130_fd_sc_hd__buf_4
XFILLER_0_172_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19116_ _04273_ _04410_ _04412_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16328_ decode.regfile.registers_21\[26\] _11061_ _11099_ _11228_ _12298_ VGND VGND
+ VPWR VPWR _12299_ sky130_fd_sc_hd__o311a_1
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_146_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_146_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19047_ _04345_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16259_ _12230_ _11486_ _12231_ VGND VGND VPWR VPWR _12232_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_81_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_222_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_222_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19949_ _03581_ _05201_ net1020 VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__and3b_1
XFILLER_0_96_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22960_ _07406_ _07408_ _07085_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21911_ _06547_ _06543_ _06544_ _06548_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22891_ _07342_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24630_ net2108 execute.io_target_pc\[4\] _08497_ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__mux2_1
X_21842_ net512 _06497_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__or2_1
XFILLER_0_223_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24561_ _09896_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_172_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21773_ _06449_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26300_ _09432_ _09472_ VGND VGND VPWR VPWR _09482_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_173_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23512_ net2459 _07890_ _07887_ VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__or3b_1
XFILLER_0_19_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20724_ _05809_ decode.id_ex_rs1_data_reg\[20\] _05798_ VGND VGND VPWR VPWR _05832_
+ sky130_fd_sc_hd__a21oi_1
X_24492_ _08426_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27280_ clknet_leaf_328_clock _00309_ VGND VGND VPWR VPWR decode.regfile.registers_31\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23443_ net2 _07846_ _07856_ _07851_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__o211a_1
X_26231_ _10141_ VGND VGND VPWR VPWR _09441_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20655_ csr._minstret_T_3\[62\] _05556_ _05784_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__o21a_1
XFILLER_0_184_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23374_ _07797_ _07798_ _07081_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26162_ _09392_ _09390_ VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__nand2_1
X_20586_ csr._minstret_T_3\[52\] _05616_ _05622_ csr._csr_read_data_T_8\[20\] _05725_
+ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25113_ _06130_ net1963 _08778_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__mux2_1
X_22325_ _06917_ _06918_ _06675_ _06919_ _06686_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26093_ _08939_ _09340_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25044_ csr._mcycle_T_2\[19\] _08710_ _08742_ _03554_ VGND VGND VPWR VPWR _08743_
+ sky130_fd_sc_hd__a211oi_1
X_29921_ clknet_leaf_334_clock _02934_ VGND VGND VPWR VPWR decode.regfile.registers_21\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_22256_ fetch.bht.bhtTable_tag\[4\]\[17\] fetch.bht.bhtTable_tag\[5\]\[17\] _06643_
+ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21207_ _10613_ _05671_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29852_ clknet_leaf_306_clock _02865_ VGND VGND VPWR VPWR decode.regfile.registers_19\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_22187_ _06781_ _06661_ _06629_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__a21o_1
XFILLER_0_178_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28803_ clknet_leaf_131_clock _01816_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21138_ _05866_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_218_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29783_ clknet_leaf_295_clock _02796_ VGND VGND VPWR VPWR decode.regfile.registers_16\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_26995_ clknet_leaf_334_clock _00024_ VGND VGND VPWR VPWR decode.regfile.registers_22\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28734_ clknet_leaf_175_clock _01747_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13960_ net2549 _10226_ _10234_ _10232_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__o211a_1
X_25946_ net2380 _09256_ _09265_ _09264_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__o211a_1
X_21069_ execute.csr_read_data_out_reg\[23\] _06014_ _06010_ VGND VGND VPWR VPWR _06021_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_31_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28665_ clknet_leaf_122_clock _01678_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13891_ _10147_ _10152_ VGND VGND VPWR VPWR _10193_ sky130_fd_sc_hd__nand2_1
X_25877_ net2252 _09213_ _09225_ _09222_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__o211a_1
X_27616_ clknet_leaf_151_clock _00645_ VGND VGND VPWR VPWR execute.io_target_pc\[25\]
+ sky130_fd_sc_hd__dfxtp_4
X_15630_ _11614_ _11617_ _11618_ VGND VGND VPWR VPWR _11619_ sky130_fd_sc_hd__o21ai_1
X_24828_ _08601_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__clkbuf_1
X_28596_ clknet_leaf_119_clock _01609_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_307 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_318 execute.io_target_pc\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27547_ clknet_leaf_41_clock _00576_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfxtp_2
X_15561_ _10649_ _10632_ _11052_ _11551_ VGND VGND VPWR VPWR _11552_ sky130_fd_sc_hd__o31a_1
XFILLER_0_57_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24759_ _08565_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_329 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _12915_ decode.regfile.registers_25\[12\] _13045_ _12812_ VGND VGND VPWR
+ VPWR _13253_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14512_ _09888_ VGND VGND VPWR VPWR _10557_ sky130_fd_sc_hd__buf_4
X_18280_ _03604_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__clkbuf_1
X_27478_ clknet_leaf_65_clock net184 VGND VGND VPWR VPWR decode.csr_write_reg sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ decode.regfile.registers_25\[4\] _11483_ _11484_ decode.regfile.registers_24\[4\]
+ VGND VGND VPWR VPWR _11485_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_29_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29217_ clknet_leaf_88_clock _02230_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17231_ decode.regfile.registers_18\[11\] _10925_ _12569_ _11023_ _11008_ VGND VGND
+ VPWR VPWR _13185_ sky130_fd_sc_hd__o2111a_1
X_26429_ net1140 _09548_ _09556_ _09553_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14443_ net582 _10506_ _10514_ _10509_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_63_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_63_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29148_ clknet_leaf_165_clock _02161_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_17162_ decode.regfile.registers_13\[9\] _12775_ _13116_ _13117_ _12664_ VGND VGND
+ VPWR VPWR _13118_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14374_ _10015_ _10474_ VGND VGND VPWR VPWR _10475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16113_ _11260_ _12087_ _12088_ _12089_ VGND VGND VPWR VPWR _12090_ sky130_fd_sc_hd__a31o_1
X_29079_ clknet_leaf_192_clock _02092_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17093_ _10940_ _12706_ decode.regfile.registers_27\[7\] _13050_ VGND VGND VPWR VPWR
+ _13051_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_78_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_78_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16044_ decode.regfile.registers_1\[19\] _11116_ _11137_ _11157_ VGND VGND VPWR VPWR
+ _12022_ sky130_fd_sc_hd__nand4_1
XFILLER_0_33_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19803_ _05045_ _05031_ _05060_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17995_ _12499_ _12490_ _12511_ decode.regfile.registers_12\[30\] _12745_ VGND VGND
+ VPWR VPWR _03392_ sky130_fd_sc_hd__o32a_1
XFILLER_0_202_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19734_ _04349_ _04303_ _04816_ _05009_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__o31a_1
X_16946_ decode.regfile.registers_19\[4\] _11013_ _11012_ _12519_ _12906_ VGND VGND
+ VPWR VPWR _12907_ sky130_fd_sc_hd__o41a_1
XFILLER_0_208_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19665_ net190 _04234_ _04256_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__o21a_1
X_16877_ decode.regfile.registers_2\[3\] _12835_ _12836_ decode.regfile.registers_3\[3\]
+ _12838_ VGND VGND VPWR VPWR _12839_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_95_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18616_ _03659_ execute.csr_read_data_out_reg\[18\] execute.io_reg_pc\[18\] _03777_
+ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__o22a_1
X_15828_ decode.regfile.registers_9\[13\] _11547_ _11192_ _11131_ VGND VGND VPWR VPWR
+ _11812_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_16_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_16_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19596_ net309 net219 _03637_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__and3_1
XFILLER_0_189_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18547_ decode.id_ex_rs2_data_reg\[24\] _03747_ _03764_ _03842_ _03845_ VGND VGND
+ VPWR VPWR _03846_ sky130_fd_sc_hd__o221a_1
X_15759_ decode.regfile.registers_16\[11\] _11359_ _11727_ _11744_ _11127_ VGND VGND
+ VPWR VPWR _11745_ sky130_fd_sc_hd__o221a_1
XFILLER_0_220_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18478_ _03776_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_215_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17429_ decode.regfile.registers_20\[16\] _11024_ _12552_ _12823_ _12824_ VGND VGND
+ VPWR VPWR _13378_ sky130_fd_sc_hd__a41o_1
XFILLER_0_74_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20440_ csr._csr_read_data_T_8\[2\] _05593_ _05516_ _05528_ _05597_ VGND VGND VPWR
+ VPWR _05598_ sky130_fd_sc_hd__a41o_1
XFILLER_0_15_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20371_ csr.io_csr_address\[7\] VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22110_ fetch.bht.bhtTable_tag\[6\]\[3\] fetch.bht.bhtTable_tag\[7\]\[3\] _06700_
+ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23090_ _07391_ _07392_ _07530_ _07531_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_63_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22041_ _06635_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__buf_6
XFILLER_0_228_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25800_ _08948_ _09179_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_215_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26780_ net2153 _09752_ _09759_ _09758_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__o211a_1
X_23992_ _08167_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25731_ _09128_ VGND VGND VPWR VPWR _09142_ sky130_fd_sc_hd__clkbuf_4
X_22943_ net92 net89 VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__and2_1
XFILLER_0_223_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28450_ clknet_leaf_146_clock _01463_ VGND VGND VPWR VPWR decode.io_id_pc\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25662_ net2260 _09095_ _09101_ _09100_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__o211a_1
X_22874_ _07333_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27401_ clknet_leaf_29_clock _00430_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_24613_ net858 execute.io_target_pc\[28\] _09897_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28381_ clknet_leaf_170_clock _01394_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21825_ _06480_ csr._csr_read_data_T_9\[1\] _06486_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_65_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25593_ net2369 _09052_ _09061_ _09059_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_121_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27332_ clknet_leaf_46_clock _00361_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_24544_ _08453_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__clkbuf_1
X_21756_ net1195 _10803_ _06439_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20707_ decode.id_ex_funct3_reg\[0\] _05804_ _05821_ VGND VGND VPWR VPWR _05822_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27263_ clknet_leaf_1_clock _00292_ VGND VGND VPWR VPWR decode.regfile.registers_30\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_24475_ _08417_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__clkbuf_1
X_21687_ _06369_ _06380_ _06391_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_134_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29002_ clknet_leaf_98_clock _02015_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26214_ net2716 _09419_ _09429_ _09418_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20638_ csr.mcycle\[28\] _05587_ _05594_ csr.minstret\[28\] VGND VGND VPWR VPWR _05770_
+ sky130_fd_sc_hd__a22o_1
X_23426_ _10670_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27194_ clknet_leaf_360_clock _00223_ VGND VGND VPWR VPWR decode.regfile.registers_28\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23357_ _07782_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26145_ _09983_ VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__buf_4
X_20569_ csr.mcycle\[18\] _05551_ _05559_ csr.minstret\[18\] VGND VGND VPWR VPWR _05711_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22308_ fetch.bht.bhtTable_tag\[2\]\[0\] fetch.bht.bhtTable_tag\[3\]\[0\] _06644_
+ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14090_ net1796 _10302_ _10310_ _10304_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__o211a_1
X_23288_ _07089_ _07714_ _07715_ _07718_ VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26076_ _09328_ VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_225_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22239_ net80 _06833_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__nor2_1
X_25027_ net708 _08730_ _08731_ _06419_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__a211oi_1
X_29904_ clknet_leaf_301_clock _02917_ VGND VGND VPWR VPWR decode.regfile.registers_20\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_17__f_clock clknet_2_2_0_clock VGND VGND VPWR VPWR clknet_5_17__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_29835_ clknet_leaf_298_clock _02848_ VGND VGND VPWR VPWR decode.regfile.registers_18\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16800_ net539 _12709_ _12710_ _12763_ _12705_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__o221a_1
X_17780_ _12967_ _03180_ _03181_ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__a31o_1
X_29766_ clknet_leaf_293_clock _02779_ VGND VGND VPWR VPWR decode.regfile.registers_16\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14992_ _10944_ _11004_ _11006_ _11007_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__a31o_1
X_26978_ net2463 _09866_ _09872_ _09865_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__o211a_1
X_28717_ clknet_leaf_102_clock _01730_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16731_ decode.regfile.registers_27\[0\] _12507_ _12520_ _12695_ decode.regfile.registers_26\[0\]
+ VGND VGND VPWR VPWR _12696_ sky130_fd_sc_hd__o32a_1
X_13943_ _10081_ _10223_ VGND VGND VPWR VPWR _10225_ sky130_fd_sc_hd__nand2_1
X_25929_ net771 _09242_ _09255_ _09250_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29697_ clknet_leaf_291_clock _02710_ VGND VGND VPWR VPWR decode.regfile.registers_14\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19450_ _04736_ _04589_ _04346_ _04408_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__and4_1
X_28648_ clknet_leaf_96_clock _01661_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16662_ _10607_ _10614_ _12557_ _10591_ VGND VGND VPWR VPWR _12627_ sky130_fd_sc_hd__nand4_2
XFILLER_0_18_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13874_ _10102_ _10177_ VGND VGND VPWR VPWR _10184_ sky130_fd_sc_hd__nand2_1
X_18401_ _03699_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__buf_6
X_15613_ decode.regfile.registers_25\[7\] _11333_ _11336_ decode.regfile.registers_24\[7\]
+ VGND VGND VPWR VPWR _11603_ sky130_fd_sc_hd__o22a_1
XFILLER_0_202_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19381_ _04253_ _04137_ _04478_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__o21a_1
X_28579_ clknet_leaf_126_clock _01592_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_104 _10773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16593_ _12557_ VGND VGND VPWR VPWR _12558_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_115 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_126 _11167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_137 _11999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18332_ decode.id_ex_rs2_data_reg\[31\] _03627_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_148 _12512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15544_ decode.regfile.registers_7\[6\] _11533_ decode.regfile.registers_6\[6\] _11534_
+ _11174_ VGND VGND VPWR VPWR _11535_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_16_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_159 _13203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18263_ _03593_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15475_ _11136_ _11464_ _11467_ VGND VGND VPWR VPWR _11468_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17214_ _13081_ _13168_ decode.regfile.registers_23\[10\] _13041_ VGND VGND VPWR
+ VPWR _13169_ sky130_fd_sc_hd__or4_1
X_14426_ net498 _10464_ _10503_ _10494_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18194_ decode.control.io_opcode\[3\] _10585_ _03518_ _03531_ VGND VGND VPWR VPWR
+ _03532_ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17145_ decode.regfile.registers_15\[9\] _10612_ _10924_ _12589_ _12673_ VGND VGND
+ VPWR VPWR _13101_ sky130_fd_sc_hd__a41o_1
XFILLER_0_163_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14357_ net505 _10463_ _10465_ _10453_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold707 fetch.bht.bhtTable_tag\[12\]\[2\] VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold718 fetch.bht.bhtTable_tag\[8\]\[16\] VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold729 fetch.bht.bhtTable_tag\[4\]\[10\] VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17076_ decode.regfile.registers_16\[7\] _13011_ _12578_ _13033_ VGND VGND VPWR VPWR
+ _13034_ sky130_fd_sc_hd__o211a_1
X_14288_ _09984_ _10420_ VGND VGND VPWR VPWR _10425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_204_1226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16027_ decode.regfile.registers_19\[18\] _11453_ _11454_ _12005_ VGND VGND VPWR
+ VPWR _12006_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2108 decode.regfile.registers_2\[5\] VGND VGND VPWR VPWR net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2119 decode.regfile.registers_10\[28\] VGND VGND VPWR VPWR net2346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1407 fetch.bht.bhtTable_tag\[14\]\[23\] VGND VGND VPWR VPWR net1634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17978_ _10930_ decode.regfile.registers_28\[30\] _12698_ VGND VGND VPWR VPWR _03375_
+ sky130_fd_sc_hd__o21a_1
Xhold1418 decode.regfile.registers_28\[2\] VGND VGND VPWR VPWR net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1429 fetch.bht.bhtTable_tag\[6\]\[5\] VGND VGND VPWR VPWR net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16929_ decode.regfile.registers_7\[4\] _12612_ _12889_ VGND VGND VPWR VPWR _12890_
+ sky130_fd_sc_hd__a21oi_1
X_19717_ _03881_ _04991_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19648_ _04906_ _04927_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_217_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_217_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19579_ _04211_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21610_ csr._mcycle_T_2\[4\] _06325_ _06323_ _06333_ _05613_ VGND VGND VPWR VPWR
+ _06335_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_133_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_213_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22590_ csr._minstret_T_3\[44\] csr._minstret_T_3\[43\] _07166_ VGND VGND VPWR VPWR
+ _07170_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21541_ _06290_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24260_ _08305_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__clkbuf_1
X_21472_ _06101_ net1554 _06252_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23211_ _07642_ _07644_ _07645_ _07075_ _06637_ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__a221o_1
X_20423_ _05561_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__clkbuf_4
X_24191_ _08085_ net1679 _08266_ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23142_ _07097_ _07576_ _07578_ _07580_ _07368_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_168_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20354_ _03721_ _03737_ _03755_ _05516_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__and4_1
XFILLER_0_114_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23073_ _07513_ _07112_ _07122_ _07515_ VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__a211o_1
X_27950_ clknet_leaf_206_clock _00972_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_164_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20285_ _10694_ _10710_ decode.id_ex_pc_reg\[14\] _05452_ _10681_ VGND VGND VPWR
+ VPWR _05465_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_164_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22024_ _06618_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__buf_4
X_26901_ net2598 _09822_ _09828_ _09825_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__o211a_1
X_27881_ clknet_leaf_25_clock _00910_ VGND VGND VPWR VPWR csr._mcycle_T_2\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_220_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29620_ clknet_leaf_280_clock _02633_ VGND VGND VPWR VPWR decode.regfile.registers_11\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_26832_ net2462 _09779_ _09788_ _09784_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1930 decode.regfile.registers_21\[21\] VGND VGND VPWR VPWR net2157 sky130_fd_sc_hd__dlygate4sd3_1
X_29551_ clknet_leaf_274_clock _02564_ VGND VGND VPWR VPWR decode.regfile.registers_9\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1941 decode.regfile.registers_14\[28\] VGND VGND VPWR VPWR net2168 sky130_fd_sc_hd__dlygate4sd3_1
X_26763_ net1642 _09710_ _09748_ _09743_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23975_ _08158_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__clkbuf_1
Xhold1952 decode.regfile.registers_26\[13\] VGND VGND VPWR VPWR net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1963 decode.io_id_pc\[23\] VGND VGND VPWR VPWR net2190 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28502_ clknet_leaf_218_clock _01515_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1974 decode.regfile.registers_16\[18\] VGND VGND VPWR VPWR net2201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25714_ _08937_ _09122_ VGND VGND VPWR VPWR _09132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22926_ fetch.bht.bhtTable_target_pc\[8\]\[2\] fetch.bht.bhtTable_target_pc\[9\]\[2\]
+ fetch.bht.bhtTable_target_pc\[10\]\[2\] fetch.bht.bhtTable_target_pc\[11\]\[2\]
+ _07107_ _07114_ VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__mux4_1
Xhold1985 csr._minstret_T_3\[54\] VGND VGND VPWR VPWR net2212 sky130_fd_sc_hd__dlygate4sd3_1
X_29482_ clknet_leaf_263_clock _02495_ VGND VGND VPWR VPWR decode.regfile.registers_7\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1996 decode.regfile.registers_13\[26\] VGND VGND VPWR VPWR net2223 sky130_fd_sc_hd__dlygate4sd3_1
X_26694_ _09708_ VGND VGND VPWR VPWR _09710_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28433_ clknet_leaf_244_clock _01446_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_25645_ net2173 _09082_ _09091_ _09087_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__o211a_1
X_22857_ net947 _10807_ _07324_ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28364_ clknet_leaf_220_clock _01377_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21808_ net2533 _06467_ _06474_ _10546_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25576_ _09023_ VGND VGND VPWR VPWR _09052_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ _09954_ VGND VGND VPWR VPWR _09955_ sky130_fd_sc_hd__buf_4
X_22788_ net934 _10881_ _07286_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27315_ clknet_leaf_327_clock _00344_ VGND VGND VPWR VPWR decode.id_ex_ex_rd_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_24527_ _08087_ net1540 _08439_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21739_ net873 _10817_ _06428_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__mux2_1
X_28295_ clknet_leaf_164_clock _00017_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27246_ clknet_leaf_1_clock _00275_ VGND VGND VPWR VPWR decode.regfile.registers_29\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15260_ _10960_ decode.regfile.registers_28\[1\] _11067_ _11038_ _10994_ VGND VGND
+ VPWR VPWR _11256_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_97_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24458_ _08408_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14211_ _09975_ _10377_ VGND VGND VPWR VPWR _10381_ sky130_fd_sc_hd__nand2_1
X_23409_ net91 _07819_ _07830_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27177_ clknet_leaf_362_clock _00206_ VGND VGND VPWR VPWR decode.regfile.registers_27\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_15191_ decode.regfile.registers_11\[0\] _11181_ _11184_ decode.regfile.registers_10\[0\]
+ _11187_ VGND VGND VPWR VPWR _11188_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_229_Right_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24389_ net1477 execute.io_target_pc\[17\] _08367_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_9 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ net493 _10332_ _10340_ _10328_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__o211a_1
X_26128_ _08975_ _09328_ VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_1202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14073_ _10025_ _10299_ VGND VGND VPWR VPWR _10301_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_56_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26059_ _09025_ _09330_ VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__nand2_1
X_18950_ _04248_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__clkbuf_4
X_17901_ net518 _12872_ _03263_ _03300_ _03073_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__o221a_1
X_18881_ _04087_ _03701_ _03688_ decode.id_ex_rs1_data_reg\[15\] _04090_ VGND VGND
+ VPWR VPWR _04180_ sky130_fd_sc_hd__o221a_4
XFILLER_0_218_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17832_ decode.regfile.registers_1\[26\] _12631_ _12933_ _12508_ _03232_ VGND VGND
+ VPWR VPWR _03233_ sky130_fd_sc_hd__o221a_1
X_29818_ clknet_leaf_306_clock _02831_ VGND VGND VPWR VPWR decode.regfile.registers_18\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_17763_ decode.regfile.registers_14\[24\] _12670_ _03151_ _03165_ VGND VGND VPWR
+ VPWR _03166_ sky130_fd_sc_hd__o22a_1
X_14975_ _10998_ VGND VGND VPWR VPWR _10999_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29749_ clknet_leaf_285_clock _02762_ VGND VGND VPWR VPWR decode.regfile.registers_15\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16714_ _12678_ VGND VGND VPWR VPWR _12679_ sky130_fd_sc_hd__clkbuf_4
X_19502_ _04186_ _04785_ _04763_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__nand3_1
X_13926_ net1581 _10213_ _10215_ _10206_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17694_ decode.regfile.registers_22\[22\] _13100_ _03098_ _13289_ VGND VGND VPWR
+ VPWR _03099_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19433_ _04640_ _04719_ _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_187_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16645_ _12609_ VGND VGND VPWR VPWR _12610_ sky130_fd_sc_hd__clkbuf_4
X_13857_ _10064_ _10164_ VGND VGND VPWR VPWR _10174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19364_ _04270_ _04337_ _04343_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_191_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16576_ _12540_ VGND VGND VPWR VPWR _12541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13788_ _10060_ memory.io_wb_readdata\[28\] _10124_ VGND VGND VPWR VPWR _10125_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18315_ decode.id_ex_rs2_data_reg\[23\] _03616_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15527_ decode.regfile.registers_20\[5\] _11102_ _11221_ _11518_ VGND VGND VPWR VPWR
+ _11519_ sky130_fd_sc_hd__a211o_1
XFILLER_0_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19295_ _04580_ _04581_ _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18246_ _03567_ net2366 _03578_ _03580_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_199_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15458_ _11435_ decode.regfile.registers_22\[4\] _11450_ _10979_ _10991_ VGND VGND
+ VPWR VPWR _11451_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_167_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14409_ _10102_ _10487_ VGND VGND VPWR VPWR _10495_ sky130_fd_sc_hd__nand2_1
X_18177_ _10576_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15389_ decode.regfile.registers_10\[2\] _10639_ _11132_ _11364_ _11383_ VGND VGND
+ VPWR VPWR _11384_ sky130_fd_sc_hd__o311a_1
XFILLER_0_13_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap201 _10080_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_4
Xhold504 decode.regfile.registers_25\[11\] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ _12516_ _13080_ _13082_ _13084_ VGND VGND VPWR VPWR _13085_ sky130_fd_sc_hd__a31o_1
Xhold515 decode.regfile.registers_23\[16\] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold526 fetch.bht.bhtTable_target_pc\[8\]\[20\] VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold537 decode.regfile.registers_28\[10\] VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold548 decode.regfile.registers_31\[31\] VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17059_ decode.regfile.registers_4\[7\] _12617_ _12619_ decode.regfile.registers_5\[7\]
+ _12622_ VGND VGND VPWR VPWR _13017_ sky130_fd_sc_hd__a221o_1
Xhold559 execute.csr_write_data_out_reg\[19\] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_206_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_206_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20070_ _05284_ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1204 fetch.bht.bhtTable_target_pc\[6\]\[21\] VGND VGND VPWR VPWR net1431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 fetch.bht.bhtTable_target_pc\[8\]\[23\] VGND VGND VPWR VPWR net1442 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 fetch.bht.bhtTable_tag\[11\]\[20\] VGND VGND VPWR VPWR net1453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 fetch.bht.bhtTable_target_pc\[0\]\[26\] VGND VGND VPWR VPWR net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 fetch.bht.bhtTable_target_pc\[6\]\[12\] VGND VGND VPWR VPWR net1475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 fetch.bht.bhtTable_target_pc\[14\]\[27\] VGND VGND VPWR VPWR net1486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23760_ _06122_ net1575 _08030_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20972_ _05968_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22711_ net2757 _07235_ _07244_ _07234_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23691_ net789 _10817_ _07992_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25430_ net196 VGND VGND VPWR VPWR _08964_ sky130_fd_sc_hd__clkbuf_8
X_22642_ csr._minstret_T_3\[62\] csr._minstret_T_3\[61\] _07202_ VGND VGND VPWR VPWR
+ _07205_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22573_ csr.minstret\[28\] csr.minstret\[29\] _07156_ VGND VGND VPWR VPWR _07157_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25361_ _09992_ VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__buf_4
XFILLER_0_192_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27100_ clknet_leaf_348_clock _00129_ VGND VGND VPWR VPWR decode.regfile.registers_25\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_24312_ _08074_ net1827 _08323_ VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21524_ _06153_ net1373 _06274_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__mux2_1
X_28080_ clknet_leaf_196_clock _01102_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25292_ _08876_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27031_ clknet_leaf_332_clock _00060_ VGND VGND VPWR VPWR decode.regfile.registers_23\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_21455_ _06243_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__clkbuf_1
X_24243_ _08296_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20406_ csr.mcycle\[0\] _05561_ _05563_ csr._csr_read_data_T_9\[0\] _05565_ VGND
+ VGND VPWR VPWR _05566_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_92_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24174_ _08068_ net1989 _08255_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21386_ _06134_ net1275 _06199_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23125_ _07082_ _07560_ _07564_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_187_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20337_ _05420_ _05390_ _05504_ _05454_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__o211a_1
X_28982_ clknet_leaf_126_clock _01995_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27933_ clknet_leaf_165_clock _00006_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_23056_ _07368_ _07496_ _05246_ _07499_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_101_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput68 net68 VGND VGND VPWR VPWR io_fetch_address[10] sky130_fd_sc_hd__clkbuf_4
X_20268_ _10706_ decode.id_ex_pc_reg\[10\] _10689_ _05440_ VGND VGND VPWR VPWR _05452_
+ sky130_fd_sc_hd__and4_1
Xoutput79 net79 VGND VGND VPWR VPWR io_fetch_address[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_216_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22007_ net526 _06600_ _06608_ _06605_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_125_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27864_ clknet_leaf_320_clock _00893_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20199_ _05396_ _05397_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__or2b_1
Xhold2450 _01123_ VGND VGND VPWR VPWR net2677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2461 decode.regfile.registers_0\[23\] VGND VGND VPWR VPWR net2688 sky130_fd_sc_hd__dlygate4sd3_1
X_26815_ _09751_ VGND VGND VPWR VPWR _09779_ sky130_fd_sc_hd__buf_2
X_29603_ clknet_leaf_276_clock _02616_ VGND VGND VPWR VPWR decode.regfile.registers_11\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2472 csr.mcycle\[29\] VGND VGND VPWR VPWR net2699 sky130_fd_sc_hd__buf_1
XFILLER_0_157_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27795_ clknet_leaf_305_clock _00824_ VGND VGND VPWR VPWR memory.io_wb_readdata\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2483 decode.regfile.registers_17\[18\] VGND VGND VPWR VPWR net2710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2494 decode.regfile.registers_14\[27\] VGND VGND VPWR VPWR net2721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29534_ clknet_leaf_312_clock _02547_ VGND VGND VPWR VPWR decode.regfile.registers_9\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1760 decode.regfile.registers_5\[31\] VGND VGND VPWR VPWR net1987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1771 fetch.bht.bhtTable_tag\[10\]\[10\] VGND VGND VPWR VPWR net1998 sky130_fd_sc_hd__dlygate4sd3_1
X_14760_ csr.io_mem_pc\[17\] VGND VGND VPWR VPWR _10803_ sky130_fd_sc_hd__clkbuf_8
X_26746_ net1765 _09736_ _09739_ _09730_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_86_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1782 fetch.bht.bhtTable_target_pc\[0\]\[24\] VGND VGND VPWR VPWR net2009 sky130_fd_sc_hd__dlygate4sd3_1
X_23958_ _08149_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1793 _01227_ VGND VGND VPWR VPWR net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13711_ _10003_ VGND VGND VPWR VPWR _10060_ sky130_fd_sc_hd__clkbuf_4
X_22909_ net75 _06886_ _06862_ net222 VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__a2bb2o_1
X_29465_ clknet_leaf_249_clock _02478_ VGND VGND VPWR VPWR decode.regfile.registers_6\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14691_ _10732_ execute.io_target_pc\[23\] _10733_ execute.io_target_pc\[31\] VGND
+ VGND VPWR VPWR _10734_ sky130_fd_sc_hd__a22oi_1
X_26677_ _09432_ _09689_ VGND VGND VPWR VPWR _09699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23889_ _08113_ net1368 _07940_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28416_ clknet_leaf_52_clock _01429_ VGND VGND VPWR VPWR decode.control.io_opcode\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16430_ _11364_ _12396_ _12397_ VGND VGND VPWR VPWR _12398_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13642_ net1157 _09938_ _10000_ _09957_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__o211a_1
X_25628_ _09067_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_224_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29396_ clknet_leaf_259_clock _02409_ VGND VGND VPWR VPWR decode.regfile.registers_4\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28347_ clknet_leaf_197_clock _01360_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16361_ decode.regfile.registers_16\[27\] _11123_ VGND VGND VPWR VPWR _12331_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25559_ net1850 _09039_ _09042_ _09033_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_45_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13573_ _09937_ VGND VGND VPWR VPWR _09938_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18100_ _03476_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15312_ _11307_ VGND VGND VPWR VPWR _11308_ sky130_fd_sc_hd__clkbuf_2
X_19080_ _04375_ _04377_ _04324_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__mux2_1
X_28278_ clknet_leaf_59_clock _01300_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ decode.regfile.registers_22\[25\] _11096_ _11232_ _12263_ VGND VGND VPWR
+ VPWR _12264_ sky130_fd_sc_hd__a211o_1
XFILLER_0_227_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18031_ decode.regfile.registers_14\[31\] _10923_ _12876_ _12555_ VGND VGND VPWR
+ VPWR _03427_ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15243_ _11078_ _11081_ _11234_ _11239_ VGND VGND VPWR VPWR _11240_ sky130_fd_sc_hd__o31a_1
X_27229_ clknet_leaf_1_clock _00258_ VGND VGND VPWR VPWR decode.regfile.registers_29\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15174_ decode.regfile.registers_7\[0\] _11092_ _11167_ _11170_ decode.regfile.registers_6\[0\]
+ VGND VGND VPWR VPWR _11171_ sky130_fd_sc_hd__a32o_1
XFILLER_0_227_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14125_ _09930_ _10194_ _10149_ _10150_ VGND VGND VPWR VPWR _10330_ sky130_fd_sc_hd__and4b_1
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19982_ net462 _05217_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14056_ _09964_ _10288_ VGND VGND VPWR VPWR _10292_ sky130_fd_sc_hd__nand2_1
X_18933_ _04006_ _04228_ _04231_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__and3_1
XFILLER_0_197_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18864_ decode.id_ex_rs2_data_reg\[10\] _03796_ net204 _04162_ _03727_ VGND VGND
+ VPWR VPWR _04163_ sky130_fd_sc_hd__o311a_2
XFILLER_0_101_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_201_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17815_ _13339_ _03214_ _03215_ _03216_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__a31o_1
X_18795_ _03707_ decode.id_ex_imm_reg\[15\] _04093_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_94_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17746_ decode.regfile.registers_19\[24\] _12679_ _12906_ VGND VGND VPWR VPWR _03149_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_221_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14958_ _10974_ _10984_ VGND VGND VPWR VPWR _10985_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_193_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_193_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13909_ _10131_ VGND VGND VPWR VPWR _10206_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17677_ decode.regfile.registers_4\[22\] _12548_ _13145_ decode.regfile.registers_5\[22\]
+ _12625_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__a221o_1
X_14889_ _10925_ VGND VGND VPWR VPWR _10926_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_212_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16628_ _10609_ _10616_ _12592_ _10593_ VGND VGND VPWR VPWR _12593_ sky130_fd_sc_hd__and4_1
X_19416_ _04149_ _04166_ _03989_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16559_ _11021_ VGND VGND VPWR VPWR _12524_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19347_ _04637_ _04635_ _04452_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19278_ _03863_ _04338_ _04307_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18229_ csr.mcycle\[21\] csr.mcycle\[24\] csr.mcycle\[23\] _03563_ VGND VGND VPWR
+ VPWR _03564_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21240_ _10807_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__buf_2
XFILLER_0_131_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold301 decode.regfile.registers_21\[15\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 decode.regfile.registers_31\[1\] VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__buf_1
Xhold323 decode.regfile.registers_22\[10\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold334 decode.regfile.registers_27\[20\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21171_ _06074_ _06070_ net1956 VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_229_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold345 csr.meie VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold356 decode.regfile.registers_13\[1\] VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 decode.regfile.registers_22\[11\] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__dlygate4sd3_1
X_20122_ _00565_ _05226_ _05331_ _05239_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__o22a_1
Xhold378 decode.regfile.registers_31\[28\] VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__buf_1
Xhold389 decode.regfile.registers_5\[15\] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_225_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_225_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20053_ _05269_ _05270_ _05260_ _05265_ _05261_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__o221a_1
X_24930_ net468 _08665_ net2766 VGND VGND VPWR VPWR _08667_ sky130_fd_sc_hd__a21oi_1
Xhold1001 fetch.bht.bhtTable_tag\[3\]\[11\] VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 fetch.bht.bhtTable_tag\[10\]\[12\] VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__dlygate4sd3_1
X_24861_ _08618_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__clkbuf_1
Xhold1023 decode.regfile.registers_17\[17\] VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 fetch.bht.bhtTable_tag\[0\]\[15\] VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 fetch.bht.bhtTable_target_pc\[1\]\[16\] VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1056 fetch.bht.bhtTable_target_pc\[3\]\[24\] VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__dlygate4sd3_1
X_26600_ _09430_ _09645_ VGND VGND VPWR VPWR _09655_ sky130_fd_sc_hd__nand2_1
X_23812_ execute.io_target_pc\[6\] VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__buf_2
XFILLER_0_217_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1067 fetch.bht.bhtTable_target_pc\[9\]\[0\] VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27580_ clknet_leaf_171_clock _00609_ VGND VGND VPWR VPWR csr.io_mem_pc\[21\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_159_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24792_ _08582_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__clkbuf_1
Xhold1078 decode.regfile.registers_27\[15\] VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 fetch.bht.bhtTable_target_pc\[12\]\[27\] VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26531_ _09436_ _09577_ VGND VGND VPWR VPWR _09615_ sky130_fd_sc_hd__nand2_1
X_23743_ _06105_ net1886 _09907_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20955_ execute.io_reg_pc\[4\] _05915_ _05911_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29250_ clknet_leaf_233_clock _02263_ VGND VGND VPWR VPWR decode.regfile.registers_0\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26462_ _09443_ _09533_ VGND VGND VPWR VPWR _09575_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_81_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23674_ net1530 _10771_ _07983_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20886_ _05858_ _05921_ net60 VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__and3_1
XFILLER_0_177_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28201_ clknet_leaf_63_clock _01223_ VGND VGND VPWR VPWR csr.mscratch\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25413_ _08952_ _08946_ VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__nand2_1
X_22625_ _07192_ _07193_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__nor2_1
X_29181_ clknet_leaf_162_clock _02194_ VGND VGND VPWR VPWR fetch.btb.btbTable\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_1324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26393_ net1491 _09534_ _09536_ _09525_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28132_ clknet_leaf_222_clock _01154_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25344_ _10240_ _03672_ _08903_ VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__and3_1
XFILLER_0_192_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22556_ csr._minstret_T_3\[36\] _07144_ _06336_ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21507_ _06136_ net2147 _06263_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__mux2_1
X_28063_ clknet_leaf_190_clock _01085_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_25275_ _08867_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22487_ _07081_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_40_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27014_ clknet_leaf_342_clock _00043_ VGND VGND VPWR VPWR decode.regfile.registers_22\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_79_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24226_ _08287_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21438_ _06234_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24157_ _08051_ net1895 _06274_ VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__mux2_1
X_21369_ _06117_ net1665 _06188_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23108_ net69 net68 _06718_ _07472_ net226 VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__a41o_1
X_24088_ _08216_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__clkbuf_1
X_28965_ clknet_leaf_136_clock _01978_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold890 fetch.bht.bhtTable_target_pc\[11\]\[1\] VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15930_ _10959_ decode.regfile.registers_26\[16\] _11447_ _11348_ _10993_ VGND VGND
+ VPWR VPWR _11911_ sky130_fd_sc_hd__o2111a_1
X_23039_ _07473_ _07483_ _07368_ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__mux2_1
X_27916_ clknet_leaf_66_clock _00945_ VGND VGND VPWR VPWR csr.io_csr_write_address\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_88_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28896_ clknet_leaf_170_clock _01909_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_110_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_144_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15861_ _11842_ _11539_ _11843_ _11296_ VGND VGND VPWR VPWR _11844_ sky130_fd_sc_hd__o211ai_2
X_27847_ clknet_leaf_325_clock _00876_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2280 decode.regfile.registers_2\[25\] VGND VGND VPWR VPWR net2507 sky130_fd_sc_hd__dlygate4sd3_1
X_17600_ _03005_ _03006_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14812_ _10775_ _10853_ _10854_ VGND VGND VPWR VPWR _10855_ sky130_fd_sc_hd__o21ai_1
Xhold2291 decode.regfile.registers_16\[27\] VGND VGND VPWR VPWR net2518 sky130_fd_sc_hd__dlygate4sd3_1
X_18580_ _03874_ _03673_ _03877_ _03878_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__and4b_1
X_15792_ decode.regfile.registers_11\[12\] _11181_ _11690_ _10640_ VGND VGND VPWR
+ VPWR _11777_ sky130_fd_sc_hd__o2bb2a_1
X_27778_ clknet_leaf_34_clock _00807_ VGND VGND VPWR VPWR memory.io_wb_readdata\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1590 fetch.bht.bhtTable_target_pc\[13\]\[29\] VGND VGND VPWR VPWR net1817 sky130_fd_sc_hd__dlygate4sd3_1
X_17531_ _12682_ decode.regfile.registers_21\[18\] _12806_ _13477_ VGND VGND VPWR
+ VPWR _13478_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14743_ decode.id_ex_pc_reg\[23\] VGND VGND VPWR VPWR _10786_ sky130_fd_sc_hd__clkbuf_4
X_26729_ _09701_ VGND VGND VPWR VPWR _09730_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29517_ clknet_leaf_265_clock _02530_ VGND VGND VPWR VPWR decode.regfile.registers_8\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17462_ _13091_ _13176_ decode.regfile.registers_27\[16\] _13050_ VGND VGND VPWR
+ VPWR _13411_ sky130_fd_sc_hd__or4_1
X_29448_ clknet_leaf_254_clock _02461_ VGND VGND VPWR VPWR decode.regfile.registers_6\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14674_ execute.io_target_pc\[21\] VGND VGND VPWR VPWR _10717_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19201_ _04279_ _04019_ _04321_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16413_ _12133_ net605 _12346_ _12381_ _12132_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__o221a_1
XFILLER_0_200_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13625_ net2475 _09938_ _09985_ _09957_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__o211a_1
X_17393_ decode.regfile.registers_2\[15\] _10608_ _12636_ _12639_ VGND VGND VPWR VPWR
+ _13343_ sky130_fd_sc_hd__a31o_1
X_29379_ clknet_leaf_255_clock _02392_ VGND VGND VPWR VPWR decode.regfile.registers_4\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19132_ _04427_ _04428_ _04273_ _04349_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__and4b_1
X_16344_ decode.regfile.registers_3\[27\] _11110_ _11141_ _11145_ VGND VGND VPWR VPWR
+ _12314_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13556_ csr.meie csr.ie net33 VGND VGND VPWR VPWR _09923_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19063_ _04349_ _04357_ _04358_ _04360_ _04346_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__a2111o_1
X_16275_ decode.regfile.registers_4\[25\] _11178_ _11143_ _11091_ VGND VGND VPWR VPWR
+ _12247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18014_ decode.regfile.registers_7\[31\] _10617_ _13020_ _12888_ VGND VGND VPWR VPWR
+ _03410_ sky130_fd_sc_hd__a31o_1
X_15226_ _11222_ VGND VGND VPWR VPWR _11223_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15157_ _11153_ VGND VGND VPWR VPWR _11154_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14108_ _10107_ _10312_ VGND VGND VPWR VPWR _10321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19965_ _10689_ _03627_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15088_ _11084_ VGND VGND VPWR VPWR _11085_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_361_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_361_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14039_ net2499 _10271_ _10280_ _10275_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18916_ _03863_ _03861_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__or2_1
XFILLER_0_226_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19896_ _04452_ _05163_ _05164_ _04505_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_219_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18847_ _03658_ execute.csr_read_data_out_reg\[11\] execute.io_reg_pc\[11\] _03662_
+ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__o22a_1
XFILLER_0_207_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18778_ memory.csr_read_data_out_reg\[14\] _09986_ _10051_ VGND VGND VPWR VPWR _04077_
+ sky130_fd_sc_hd__o21ba_2
XFILLER_0_136_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17729_ _03113_ _03132_ _12566_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20740_ _05818_ decode.id_ex_rs1_data_reg\[27\] _03585_ VGND VGND VPWR VPWR _05841_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20671_ _05797_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22410_ _06699_ _06997_ _06999_ _07004_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__o2bb2a_1
X_23390_ _06795_ _07783_ net88 VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22341_ _06933_ _06678_ _06631_ _06935_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_314_clock clknet_5_18__leaf_clock VGND VGND VPWR VPWR clknet_leaf_314_clock
+ sky130_fd_sc_hd__clkbuf_8
X_25060_ net1787 _08751_ _08753_ _06327_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__a211oi_1
X_22272_ fetch.bht.bhtTable_tag\[14\]\[6\] fetch.bht.bhtTable_tag\[15\]\[6\] _06700_
+ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_227_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24011_ net1427 execute.io_target_pc\[26\] _07960_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__mux2_1
X_21223_ net984 _06107_ _09912_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_227_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold153 io_fetch_data[13] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold164 fetch.bht.bhtTable_valid\[12\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21154_ _06062_ _06070_ net2136 VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_180_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold175 decode.regfile.registers_30\[16\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_180_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold186 fetch.btb.btbTable\[0\]\[0\] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 fetch.btb.btbTable\[1\]\[0\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_329_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_329_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20105_ _05308_ _05312_ _05309_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__o21ai_1
X_28750_ clknet_leaf_110_clock _01763_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25962_ net2576 _09270_ _09274_ _09264_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__o211a_1
X_21085_ _06029_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27701_ clknet_leaf_22_clock _00730_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_20036_ _05254_ _05255_ _05256_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__and3_1
X_24913_ csr._mcycle_T_3\[38\] csr._mcycle_T_3\[37\] _08652_ VGND VGND VPWR VPWR _08656_
+ sky130_fd_sc_hd__and3_1
X_28681_ clknet_leaf_89_clock _01694_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25893_ _08966_ _09223_ VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27632_ clknet_leaf_44_clock _00661_ VGND VGND VPWR VPWR execute.io_reg_pc\[9\] sky130_fd_sc_hd__dfxtp_1
X_24844_ _06122_ net2130 _08607_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__mux2_1
XINSDIODE1_10 _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_21 _03064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_32 _08929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_43 _09932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27563_ clknet_leaf_162_clock _00592_ VGND VGND VPWR VPWR csr.io_mem_pc\[4\] sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_54 _10073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_217_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24775_ _08573_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_178_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_65 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21987_ net1417 _06588_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__or2_1
XINSDIODE1_76 _10240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29302_ clknet_leaf_231_clock _02315_ VGND VGND VPWR VPWR decode.regfile.registers_1\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26514_ _09420_ _09602_ VGND VGND VPWR VPWR _09606_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_87 _10594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23726_ _07990_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__clkbuf_8
XINSDIODE1_98 _10655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_205_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20938_ _05950_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__clkbuf_1
X_27494_ clknet_leaf_33_clock _00523_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_95_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29233_ clknet_leaf_128_clock _02246_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26445_ _10130_ VGND VGND VPWR VPWR _09566_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23657_ net1098 _10795_ _07972_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _05912_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_42_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29164_ clknet_leaf_200_clock _02177_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22608_ net2732 _07181_ _07182_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__o21ba_1
X_26376_ _09432_ _09515_ VGND VGND VPWR VPWR _09526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14390_ _10058_ _10474_ VGND VGND VPWR VPWR _10484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23588_ _06119_ net1959 _07930_ VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28115_ clknet_leaf_90_clock _01137_ VGND VGND VPWR VPWR csr.minstret\[20\] sky130_fd_sc_hd__dfxtp_1
X_25327_ _08894_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22539_ csr.io_mret_vector\[1\] VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__inv_2
X_29095_ clknet_leaf_70_clock _02108_ VGND VGND VPWR VPWR csr._mcycle_T_3\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28046_ clknet_leaf_236_clock _01068_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16060_ decode.regfile.registers_16\[19\] _11359_ _12017_ _12037_ _11127_ VGND VGND
+ VPWR VPWR _12038_ sky130_fd_sc_hd__o221a_1
X_25258_ _08097_ net1631 _09906_ VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15011_ _11020_ VGND VGND VPWR VPWR _11021_ sky130_fd_sc_hd__clkbuf_4
X_24209_ _08103_ net1312 _06251_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__mux2_1
X_25189_ _08823_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19750_ _04190_ _04195_ _03963_ _05021_ _05024_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__a311o_1
X_28948_ clknet_leaf_118_clock _01961_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16962_ _12872_ net429 _12873_ _12922_ _12705_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__o221a_1
XFILLER_0_198_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18701_ _03675_ _03685_ decode.id_ex_rs1_data_reg\[1\] VGND VGND VPWR VPWR _04000_
+ sky130_fd_sc_hd__o21bai_4
X_15913_ _11194_ decode.regfile.registers_12\[15\] _11196_ _11894_ VGND VGND VPWR
+ VPWR _11895_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_217_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16893_ decode.regfile.registers_16\[3\] _12576_ _12579_ _12854_ VGND VGND VPWR VPWR
+ _12855_ sky130_fd_sc_hd__o211a_1
X_19681_ _04191_ _03956_ _03959_ _04525_ _04958_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__a311o_1
X_28879_ clknet_leaf_111_clock _01892_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15844_ _11260_ _11825_ _11826_ _11827_ VGND VGND VPWR VPWR _11828_ sky130_fd_sc_hd__a31o_1
X_18632_ _03927_ _03797_ _03707_ _03930_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15775_ _11344_ net457 _11725_ _11759_ _11760_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__o221a_1
X_18563_ decode.id_ex_rs1_data_reg\[30\] _03689_ _03858_ _03861_ VGND VGND VPWR VPWR
+ _03862_ sky130_fd_sc_hd__o211a_4
XFILLER_0_204_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14726_ csr.io_mem_pc\[24\] csr.io_mem_pc\[25\] _10760_ _10768_ VGND VGND VPWR VPWR
+ _10769_ sky130_fd_sc_hd__and4_4
X_17514_ decode.regfile.registers_6\[18\] _12735_ _13459_ _13460_ VGND VGND VPWR VPWR
+ _13461_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_197_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18494_ execute.io_reg_pc\[28\] _03777_ _03666_ net120 _03792_ VGND VGND VPWR VPWR
+ _03793_ sky130_fd_sc_hd__o221a_1
X_17445_ _12498_ _12489_ _12511_ decode.regfile.registers_12\[16\] _12590_ VGND VGND
+ VPWR VPWR _13394_ sky130_fd_sc_hd__o32a_1
XFILLER_0_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14657_ _10692_ execute.io_target_pc\[19\] _10693_ execute.io_target_pc\[24\] _10699_
+ VGND VGND VPWR VPWR _10700_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13608_ _09970_ _09951_ VGND VGND VPWR VPWR _09971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17376_ decode.regfile.registers_17\[14\] _12578_ _13307_ _13326_ _12564_ VGND VGND
+ VPWR VPWR _13327_ sky130_fd_sc_hd__o221a_1
X_14588_ _10630_ VGND VGND VPWR VPWR _10631_ sky130_fd_sc_hd__buf_4
XFILLER_0_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19115_ _04280_ _04282_ _04411_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__or3_2
X_16327_ decode.regfile.registers_20\[26\] _11103_ _12296_ _12297_ _11222_ VGND VGND
+ VPWR VPWR _12298_ sky130_fd_sc_hd__a221o_1
X_13539_ _09885_ VGND VGND VPWR VPWR _09914_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19046_ _04056_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__clkbuf_4
X_16258_ _10959_ decode.regfile.registers_26\[24\] _11349_ _10980_ _11347_ VGND VGND
+ VPWR VPWR _12231_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_113_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15209_ _10631_ _11035_ _11044_ _11058_ VGND VGND VPWR VPWR _11206_ sky130_fd_sc_hd__and4_2
X_16189_ decode.regfile.registers_25\[22\] _11483_ _11484_ decode.regfile.registers_24\[22\]
+ VGND VGND VPWR VPWR _12164_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_222_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_206_Left_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_222_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19948_ _05208_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19879_ _03789_ _03790_ _03803_ _05127_ _03802_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21910_ csr._mcycle_T_2\[21\] _06545_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__or2_1
X_22890_ net1317 csr.io_mem_pc\[31\] _07335_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21841_ csr.io_mret_vector\[1\] csr.io_mem_pc\[1\] _06040_ VGND VGND VPWR VPWR _06499_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24560_ _08461_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_215_Left_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21772_ net1459 _10773_ _06439_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23511_ net227 _07889_ _07896_ _07893_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_173_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20723_ _05792_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__buf_2
X_24491_ _08051_ net1686 _07276_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26230_ net1965 _09419_ _09439_ _09440_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23442_ decode.immGen._imm_T_10\[3\] _07847_ _05206_ VGND VGND VPWR VPWR _07856_
+ sky130_fd_sc_hd__or3b_1
X_20654_ csr._csr_read_data_T_8\[30\] _05617_ _05781_ _05783_ _05646_ VGND VGND VPWR
+ VPWR _05784_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26161_ _10024_ VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_253_clock clknet_5_19__leaf_clock VGND VGND VPWR VPWR clknet_leaf_253_clock
+ sky130_fd_sc_hd__clkbuf_8
X_23373_ fetch.bht.bhtTable_target_pc\[0\]\[28\] fetch.bht.bhtTable_target_pc\[1\]\[28\]
+ fetch.bht.bhtTable_target_pc\[2\]\[28\] fetch.bht.bhtTable_target_pc\[3\]\[28\]
+ _07384_ _07386_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__mux4_1
X_20585_ csr.mcycle\[20\] _05587_ _05575_ csr.minstret\[20\] VGND VGND VPWR VPWR _05725_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25112_ _08784_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_76_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22324_ fetch.bht.bhtTable_tag\[8\]\[8\] fetch.bht.bhtTable_tag\[9\]\[8\] _06616_
+ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26092_ net1774 _09343_ _09349_ _09346_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_132_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25043_ csr.mcycle\[8\] _08628_ _08635_ VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29920_ clknet_leaf_335_clock _02933_ VGND VGND VPWR VPWR decode.regfile.registers_21\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_22255_ fetch.bht.bhtTable_tag\[0\]\[17\] fetch.bht.bhtTable_tag\[1\]\[17\] fetch.bht.bhtTable_tag\[2\]\[17\]
+ fetch.bht.bhtTable_tag\[3\]\[17\] _06691_ _06677_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_72_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_224_Left_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21206_ _06098_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__clkbuf_1
X_22186_ fetch.bht.bhtTable_tag\[14\]\[25\] fetch.bht.bhtTable_tag\[15\]\[25\] _06646_
+ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__mux2_1
X_29851_ clknet_leaf_306_clock _02864_ VGND VGND VPWR VPWR decode.regfile.registers_19\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28802_ clknet_leaf_134_clock _01815_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21137_ _06061_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29782_ clknet_leaf_295_clock _02795_ VGND VGND VPWR VPWR decode.regfile.registers_16\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_26994_ clknet_leaf_333_clock _00023_ VGND VGND VPWR VPWR decode.regfile.registers_22\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_28733_ clknet_leaf_179_clock _01746_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_25945_ _08941_ _09253_ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__nand2_1
X_21068_ _06020_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20019_ decode.id_ex_imm_reg\[1\] decode.id_ex_pc_reg\[1\] _10834_ decode.id_ex_imm_reg\[2\]
+ _05234_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_31_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28664_ clknet_leaf_121_clock _01677_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_13890_ net1482 _10154_ _10192_ _10188_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__o211a_1
X_25876_ _08948_ _09223_ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27615_ clknet_leaf_151_clock _00644_ VGND VGND VPWR VPWR execute.io_target_pc\[24\]
+ sky130_fd_sc_hd__dfxtp_4
X_24827_ _06105_ net1969 _08422_ VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28595_ clknet_leaf_139_clock _01608_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_206_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_206_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27546_ clknet_leaf_44_clock _00575_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_2
X_15560_ decode.regfile.registers_11\[6\] _11070_ _11470_ _11549_ _11550_ VGND VGND
+ VPWR VPWR _11551_ sky130_fd_sc_hd__a32o_1
X_24758_ _08051_ net1389 _08563_ VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__mux2_1
XINSDIODE1_308 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_319 execute.io_target_pc\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14511_ _09891_ VGND VGND VPWR VPWR _10556_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_139_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23709_ _08005_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27477_ clknet_leaf_53_clock _00506_ VGND VGND VPWR VPWR csr.io_csr_address\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_15491_ _11335_ VGND VGND VPWR VPWR _11484_ sky130_fd_sc_hd__buf_2
X_24689_ _08051_ net1588 _06306_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ decode.regfile.registers_20\[11\] _11024_ _12553_ _12823_ _12824_ VGND VGND
+ VPWR VPWR _13184_ sky130_fd_sc_hd__a41o_1
X_29216_ clknet_leaf_99_clock _02229_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26428_ _09408_ _09545_ VGND VGND VPWR VPWR _09556_ sky130_fd_sc_hd__nand2_1
X_14442_ _09993_ _10507_ VGND VGND VPWR VPWR _10514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29147_ clknet_leaf_72_clock _02160_ VGND VGND VPWR VPWR csr.mcycle\[31\] sky130_fd_sc_hd__dfxtp_2
X_17161_ _12499_ _12490_ _12511_ decode.regfile.registers_12\[9\] _12745_ VGND VGND
+ VPWR VPWR _13117_ sky130_fd_sc_hd__o32a_1
XFILLER_0_52_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26359_ net2148 _09505_ _09516_ _09512_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__o211a_1
X_14373_ _10462_ VGND VGND VPWR VPWR _10474_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16112_ _11436_ decode.regfile.registers_26\[20\] _11676_ _11338_ _11564_ VGND VGND
+ VPWR VPWR _12089_ sky130_fd_sc_hd__o2111a_1
X_29078_ clknet_leaf_192_clock _02091_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_17092_ _12506_ VGND VGND VPWR VPWR _13050_ sky130_fd_sc_hd__buf_2
XFILLER_0_165_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28029_ clknet_leaf_194_clock _01051_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16043_ decode.regfile.registers_3\[19\] _11109_ _11141_ _11145_ VGND VGND VPWR VPWR
+ _12021_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19802_ _04618_ _05069_ _04589_ _04492_ _05074_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__a311o_1
XFILLER_0_62_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17994_ decode.regfile.registers_11\[30\] _12499_ _12504_ _12650_ _03390_ VGND VGND
+ VPWR VPWR _03391_ sky130_fd_sc_hd__o41a_1
XFILLER_0_97_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19733_ net313 _04537_ _04301_ _05008_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__or4b_1
XFILLER_0_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16945_ _12543_ VGND VGND VPWR VPWR _12906_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19664_ _03959_ _04425_ net190 VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16876_ _12837_ VGND VGND VPWR VPWR _12838_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18615_ _03699_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__clkbuf_8
X_15827_ decode.regfile.registers_8\[13\] _11284_ _11801_ _11810_ VGND VGND VPWR VPWR
+ _11811_ sky130_fd_sc_hd__o22ai_2
X_19595_ _04769_ _04876_ _04272_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15758_ _10650_ _10625_ _11053_ _11742_ _11743_ VGND VGND VPWR VPWR _11744_ sky130_fd_sc_hd__o32a_1
X_18546_ _03715_ _03725_ _03841_ _03727_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14709_ _10746_ _10749_ _10750_ _10751_ VGND VGND VPWR VPWR _10752_ sky130_fd_sc_hd__and4b_1
XFILLER_0_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15689_ _11436_ decode.regfile.registers_26\[9\] _11676_ _10980_ _11564_ VGND VGND
+ VPWR VPWR _11677_ sky130_fd_sc_hd__o2111a_1
X_18477_ _03662_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17428_ _13055_ net402 _13097_ VGND VGND VPWR VPWR _13377_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17359_ decode.regfile.registers_8\[14\] _10593_ _12549_ _12592_ _12605_ VGND VGND
+ VPWR VPWR _13310_ sky130_fd_sc_hd__a41o_1
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20370_ decode.csr_write_reg _05531_ _05532_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19029_ _04320_ _04070_ _04327_ _04249_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22040_ _00003_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_162_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23991_ net1766 execute.io_target_pc\[16\] _08164_ VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_162_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25730_ _08954_ _09136_ VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22942_ _07366_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25661_ _08960_ _09092_ VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22873_ net2292 csr.io_mem_pc\[23\] _07324_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27400_ clknet_leaf_28_clock _00429_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_4
X_24612_ _08488_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28380_ clknet_leaf_189_clock _01393_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_21824_ _06481_ csr.io_ecause\[1\] _06316_ _06470_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25592_ _08966_ _09049_ VGND VGND VPWR VPWR _09061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27331_ clknet_leaf_43_clock _00360_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_4
X_24543_ _08103_ net1057 _09902_ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21755_ _06440_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27262_ clknet_leaf_4_clock _00291_ VGND VGND VPWR VPWR decode.regfile.registers_30\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_20706_ _03728_ decode.id_ex_rs1_data_reg\[13\] VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__nand2_1
X_24474_ _08101_ net1614 _08411_ VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_192_clock clknet_5_25__leaf_clock VGND VGND VPWR VPWR clknet_leaf_192_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_163_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21686_ csr.minstret\[21\] csr.minstret\[22\] csr.minstret\[23\] csr.minstret\[24\]
+ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29001_ clknet_leaf_96_clock _02014_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26213_ _09428_ _09413_ VGND VGND VPWR VPWR _09429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23425_ _03546_ VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20637_ _05766_ _05769_ _05630_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__o21a_2
X_27193_ clknet_leaf_355_clock _00222_ VGND VGND VPWR VPWR decode.regfile.registers_28\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26144_ net564 _09373_ _09380_ _09370_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23356_ net86 net85 net220 _07740_ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20568_ _05710_ _05671_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__nor2_1
XFILLER_0_225_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22307_ _06645_ fetch.bht.bhtTable_tag\[6\]\[0\] _06690_ _06901_ VGND VGND VPWR VPWR
+ _06902_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26075_ net1844 _09329_ _09339_ _09333_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_95_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23287_ net223 _07716_ _07717_ _07064_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20499_ _05645_ _05650_ _03595_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__o21a_2
XFILLER_0_30_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25026_ net2770 _08710_ _08730_ csr.mcycle\[13\] VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__a211oi_1
X_29903_ clknet_leaf_300_clock _02916_ VGND VGND VPWR VPWR decode.regfile.registers_20\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_22238_ _06636_ _06824_ _06826_ _06830_ _06832_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__a32o_2
X_29834_ clknet_leaf_298_clock _02847_ VGND VGND VPWR VPWR decode.regfile.registers_18\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_130_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_130_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22169_ _06763_ _06678_ _06627_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14991_ _10941_ _11004_ _11006_ _11007_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__a31o_1
X_29765_ clknet_leaf_293_clock _02778_ VGND VGND VPWR VPWR decode.regfile.registers_16\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26977_ net192 _09862_ VGND VGND VPWR VPWR _09872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28716_ clknet_leaf_87_clock _01729_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13942_ net2218 _10213_ _10224_ _10219_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__o211a_1
X_16730_ _12694_ VGND VGND VPWR VPWR _12695_ sky130_fd_sc_hd__buf_2
XFILLER_0_57_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25928_ _08925_ _09253_ VGND VGND VPWR VPWR _09255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29696_ clknet_leaf_290_clock _02709_ VGND VGND VPWR VPWR decode.regfile.registers_14\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_145_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_145_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16661_ _12625_ VGND VGND VPWR VPWR _12626_ sky130_fd_sc_hd__buf_4
XFILLER_0_202_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28647_ clknet_leaf_114_clock _01660_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13873_ net2443 _10180_ _10183_ _10175_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__o211a_1
X_25859_ net761 _09213_ _09215_ _09209_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15612_ _10992_ _11066_ _11261_ _11601_ VGND VGND VPWR VPWR _11602_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18400_ net354 net228 VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__nand2_8
XFILLER_0_97_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16592_ _12556_ VGND VGND VPWR VPWR _12557_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19380_ _04376_ _04141_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__or2_1
X_28578_ clknet_leaf_133_clock _01591_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_105 _10935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_116 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_127 _11167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18331_ _03631_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__clkbuf_1
X_15543_ _10646_ _10624_ _10635_ _11082_ VGND VGND VPWR VPWR _11534_ sky130_fd_sc_hd__or4_4
X_27529_ clknet_leaf_45_clock _00558_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_2
XINSDIODE1_138 _12049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_149 _12512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18262_ fetch.bht.bhtTable_tag_MPORT_en _10907_ _03590_ _03592_ _09953_ VGND VGND
+ VPWR VPWR _03593_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15474_ decode.regfile.registers_7\[4\] _11465_ _11466_ decode.regfile.registers_6\[4\]
+ _11281_ VGND VGND VPWR VPWR _11467_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17213_ _10936_ VGND VGND VPWR VPWR _13168_ sky130_fd_sc_hd__clkbuf_2
X_14425_ _10147_ _10462_ VGND VGND VPWR VPWR _10503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18193_ decode.control.io_funct7\[5\] decode.control.io_funct7\[2\] _03523_ _03530_
+ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__o31a_1
XFILLER_0_128_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17144_ _12527_ VGND VGND VPWR VPWR _13100_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14356_ _09950_ _10464_ VGND VGND VPWR VPWR _10465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold708 decode.regfile.registers_29\[24\] VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold719 decode.regfile.registers_2\[9\] VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__dlygate4sd3_1
X_17075_ _13030_ _13032_ VGND VGND VPWR VPWR _13033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14287_ net566 _10419_ _10424_ _10411_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16026_ decode.regfile.registers_18\[18\] _11455_ _11456_ _12004_ VGND VGND VPWR
+ VPWR _12005_ sky130_fd_sc_hd__a211o_1
XFILLER_0_204_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_139_Left_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2109 fetch.bht.bhtTable_target_pc\[7\]\[11\] VGND VGND VPWR VPWR net2336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1408 fetch.bht.bhtTable_target_pc\[9\]\[21\] VGND VGND VPWR VPWR net1635 sky130_fd_sc_hd__dlygate4sd3_1
X_17977_ _10931_ decode.regfile.registers_30\[30\] _12487_ VGND VGND VPWR VPWR _03374_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_204_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1419 fetch.bht.bhtTable_tag\[12\]\[24\] VGND VGND VPWR VPWR net1646 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19716_ _04991_ _03881_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16928_ _12888_ VGND VGND VPWR VPWR _12889_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_215_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19647_ _04386_ _04476_ _04907_ _04917_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__o221a_1
XFILLER_0_205_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16859_ _10931_ net553 _12487_ VGND VGND VPWR VPWR _12821_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_217_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_217_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19578_ _04197_ _04198_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_148_Left_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_213_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18529_ _03826_ _03827_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__or2b_1
XFILLER_0_87_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21540_ _06111_ net2145 _06284_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21471_ _06251_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23210_ fetch.bht.bhtTable_target_pc\[12\]\[18\] fetch.bht.bhtTable_target_pc\[13\]\[18\]
+ fetch.bht.bhtTable_target_pc\[14\]\[18\] fetch.bht.bhtTable_target_pc\[15\]\[18\]
+ _07098_ _07100_ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20422_ _05522_ _03737_ _03721_ _05525_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__and4b_4
XFILLER_0_114_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24190_ _08269_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23141_ _07122_ _07579_ _07084_ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_168_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20353_ csr.io_csr_address\[2\] VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_157_Left_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23072_ _07072_ _07514_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__and2b_1
X_20284_ _10702_ _10682_ _05458_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__or3b_1
XFILLER_0_140_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_164_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22023_ _06617_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__buf_4
X_26900_ _09428_ _09819_ VGND VGND VPWR VPWR _09828_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_90_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27880_ clknet_leaf_25_clock _00909_ VGND VGND VPWR VPWR csr._mcycle_T_2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26831_ _09434_ _09776_ VGND VGND VPWR VPWR _09788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_215_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_62_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_215_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1920 fetch.bht.bhtTable_tag\[5\]\[17\] VGND VGND VPWR VPWR net2147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1931 csr._mcycle_T_2\[28\] VGND VGND VPWR VPWR net2158 sky130_fd_sc_hd__buf_1
X_26762_ _09441_ _09708_ VGND VGND VPWR VPWR _09748_ sky130_fd_sc_hd__nand2_1
X_29550_ clknet_leaf_274_clock _02563_ VGND VGND VPWR VPWR decode.regfile.registers_9\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_23974_ net1262 execute.io_target_pc\[8\] _08153_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__mux2_1
Xhold1942 decode.regfile.registers_25\[18\] VGND VGND VPWR VPWR net2169 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1953 decode.regfile.registers_15\[0\] VGND VGND VPWR VPWR net2180 sky130_fd_sc_hd__dlygate4sd3_1
X_28501_ clknet_leaf_233_clock _01514_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1964 decode.regfile.registers_2\[7\] VGND VGND VPWR VPWR net2191 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25713_ net1773 _09125_ _09131_ _09129_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__o211a_1
X_22925_ _07375_ _07101_ _07081_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__a21o_1
Xhold1975 fetch.bht.bhtTable_tag\[6\]\[11\] VGND VGND VPWR VPWR net2202 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1986 decode.io_id_pc\[4\] VGND VGND VPWR VPWR net2213 sky130_fd_sc_hd__dlygate4sd3_1
X_26693_ _09708_ VGND VGND VPWR VPWR _09709_ sky130_fd_sc_hd__clkbuf_4
X_29481_ clknet_leaf_263_clock _02494_ VGND VGND VPWR VPWR decode.regfile.registers_7\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1997 fetch.bht.bhtTable_tag\[0\]\[17\] VGND VGND VPWR VPWR net2224 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_166_Left_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28432_ clknet_leaf_246_clock _01445_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_25644_ _08943_ _09079_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__nand2_1
X_22856_ _09896_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_77_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_77_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28363_ clknet_leaf_165_clock _01376_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_21807_ csr._mcycle_T_2\[3\] _06467_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25575_ net2361 _09039_ _09051_ _09046_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22787_ _07288_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_26_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27314_ clknet_leaf_42_clock _00343_ VGND VGND VPWR VPWR decode.id_ex_ex_rd_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_24526_ _08444_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28294_ clknet_leaf_238_clock _00018_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_21738_ _06431_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27245_ clknet_leaf_4_clock _00274_ VGND VGND VPWR VPWR decode.regfile.registers_29\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24457_ _08085_ net1415 _08400_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21669_ csr.minstret\[17\] csr.minstret\[18\] csr.minstret\[19\] _06369_ VGND VGND
+ VPWR VPWR _06378_ sky130_fd_sc_hd__and4_1
XFILLER_0_163_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14210_ net1645 _10376_ _10380_ _10369_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_193_Right_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23408_ net91 _07819_ _07087_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_948 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27176_ clknet_leaf_362_clock _00205_ VGND VGND VPWR VPWR decode.regfile.registers_27\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15190_ _11186_ VGND VGND VPWR VPWR _11187_ sky130_fd_sc_hd__buf_4
X_24388_ _08371_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14141_ _09999_ _10333_ VGND VGND VPWR VPWR _10340_ sky130_fd_sc_hd__nand2_1
X_26127_ net1651 _09330_ _09368_ _09359_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__o211a_1
X_23339_ fetch.bht.bhtTable_target_pc\[0\]\[26\] fetch.bht.bhtTable_target_pc\[1\]\[26\]
+ fetch.bht.bhtTable_target_pc\[2\]\[26\] fetch.bht.bhtTable_target_pc\[3\]\[26\]
+ _07669_ _07656_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_15_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14072_ net497 _10287_ _10300_ _10291_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__o211a_1
X_26058_ _09328_ VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25009_ net2483 _08704_ _08719_ VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__a21oi_1
X_17900_ _02997_ _12767_ _12965_ decode.regfile.registers_29\[27\] _03299_ VGND VGND
+ VPWR VPWR _03300_ sky130_fd_sc_hd__o221a_1
X_18880_ _04153_ _04176_ _04178_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_218_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17831_ _12530_ _10591_ _12557_ decode.regfile.registers_0\[26\] VGND VGND VPWR VPWR
+ _03232_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29817_ clknet_leaf_313_clock _02830_ VGND VGND VPWR VPWR decode.regfile.registers_17\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17762_ decode.regfile.registers_12\[24\] _12542_ _12723_ _12659_ _03164_ VGND VGND
+ VPWR VPWR _03165_ sky130_fd_sc_hd__o311a_1
X_29748_ clknet_leaf_285_clock _02761_ VGND VGND VPWR VPWR decode.regfile.registers_15\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_14974_ _10973_ VGND VGND VPWR VPWR _10998_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19501_ _04785_ _04763_ _04186_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__a21o_1
X_16713_ _12677_ VGND VGND VPWR VPWR _12678_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13925_ _10036_ _10210_ VGND VGND VPWR VPWR _10215_ sky130_fd_sc_hd__nand2_1
X_17693_ _12822_ decode.regfile.registers_21\[22\] _13164_ _03097_ VGND VGND VPWR
+ VPWR _03098_ sky130_fd_sc_hd__o211a_1
X_29679_ clknet_leaf_283_clock _02692_ VGND VGND VPWR VPWR decode.regfile.registers_13\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19432_ _04376_ _04141_ _04645_ _04144_ _04165_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_202_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13856_ net565 _10167_ _10173_ _10162_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16644_ _10607_ _10614_ _12522_ _10591_ VGND VGND VPWR VPWR _12609_ sky130_fd_sc_hd__and4_1
XFILLER_0_186_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19363_ _04546_ _04653_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_191_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13787_ _10060_ memory.io_wb_aluresult\[28\] _10021_ VGND VGND VPWR VPWR _10124_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16575_ _12539_ VGND VGND VPWR VPWR _12540_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18314_ _03622_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15526_ decode.regfile.registers_19\[5\] _11354_ _11218_ _11517_ VGND VGND VPWR VPWR
+ _11518_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19294_ _04496_ _04583_ _04584_ _04586_ _04445_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18245_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__buf_6
X_15457_ _11404_ VGND VGND VPWR VPWR _11450_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14408_ net450 _10490_ _10493_ _10494_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18176_ _12553_ _12569_ _10940_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__and3_2
X_15388_ _11366_ _11380_ _11382_ VGND VGND VPWR VPWR _11383_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap202 _03815_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
X_17127_ _10927_ decode.regfile.registers_24\[8\] _10933_ _13083_ _12862_ VGND VGND
+ VPWR VPWR _13084_ sky130_fd_sc_hd__o2111a_1
X_14339_ net721 _10447_ _10454_ _10453_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold505 decode.regfile.registers_27\[0\] VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold516 decode.regfile.registers_14\[6\] VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 _08375_ VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 fetch.bht.bhtTable_tag\[2\]\[4\] VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17058_ decode.regfile.registers_3\[7\] _12628_ _13013_ _13015_ VGND VGND VPWR VPWR
+ _13016_ sky130_fd_sc_hd__o22a_1
Xhold549 csr._mcycle_T_3\[37\] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_206_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16009_ decode.regfile.registers_7\[18\] _11465_ _11466_ decode.regfile.registers_6\[18\]
+ _11281_ VGND VGND VPWR VPWR _11988_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_206_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_198_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 fetch.bht.bhtTable_target_pc\[6\]\[3\] VGND VGND VPWR VPWR net1432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_198_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1216 csr.minstret\[11\] VGND VGND VPWR VPWR net1443 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 fetch.bht.bhtTable_target_pc\[4\]\[5\] VGND VGND VPWR VPWR net1454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1238 fetch.bht.bhtTable_target_pc\[12\]\[25\] VGND VGND VPWR VPWR net1465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1249 execute.csr_write_address_out_reg\[1\] VGND VGND VPWR VPWR net1476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20971_ execute.io_reg_pc\[11\] _05965_ _05961_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22710_ csr._mcycle_T_2\[29\] _07236_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23690_ _07995_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22641_ csr._minstret_T_3\[61\] _07202_ net2460 VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_157_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25360_ net1842 _08906_ _08915_ _07247_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__o211a_1
X_22572_ _07155_ _06399_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24311_ _08331_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21523_ _06279_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25291_ _08869_ decode.regfile.registers_0\[7\] VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__and2_1
XFILLER_0_185_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27030_ clknet_leaf_331_clock _00059_ VGND VGND VPWR VPWR decode.regfile.registers_23\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_24242_ _08070_ net1901 _08289_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21454_ _06145_ net1910 _06241_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20405_ _05564_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_92_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24173_ _08260_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21385_ _06205_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23124_ _07561_ _07072_ _07075_ _07563_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_187_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20336_ _05502_ _05503_ _05416_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28981_ clknet_leaf_115_clock _01994_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_187_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1091 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27932_ clknet_leaf_162_clock _00007_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_23055_ _07497_ _07498_ _07368_ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__a21oi_1
Xoutput69 net69 VGND VGND VPWR VPWR io_fetch_address[11] sky130_fd_sc_hd__clkbuf_4
X_20267_ _10689_ _05449_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22006_ csr.mscratch\[25\] _06601_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__or2_1
X_20198_ decode.id_ex_imm_reg\[27\] _10854_ _05395_ _05392_ VGND VGND VPWR VPWR _05397_
+ sky130_fd_sc_hd__o211ai_1
X_27863_ clknet_leaf_321_clock _00892_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2440 decode.regfile.registers_11\[26\] VGND VGND VPWR VPWR net2667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2451 decode.regfile.registers_0\[30\] VGND VGND VPWR VPWR net2678 sky130_fd_sc_hd__dlygate4sd3_1
X_29602_ clknet_leaf_276_clock _02615_ VGND VGND VPWR VPWR decode.regfile.registers_11\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26814_ net1341 _09766_ _09778_ _09771_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__o211a_1
Xhold2462 csr._csr_read_data_T_8\[28\] VGND VGND VPWR VPWR net2689 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2473 decode.regfile.registers_12\[25\] VGND VGND VPWR VPWR net2700 sky130_fd_sc_hd__dlygate4sd3_1
X_27794_ clknet_leaf_316_clock _00823_ VGND VGND VPWR VPWR memory.io_wb_readdata\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2484 _10733_ VGND VGND VPWR VPWR net2711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1750 fetch.bht.bhtTable_target_pc\[12\]\[28\] VGND VGND VPWR VPWR net1977 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_174_Left_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2495 _10743_ VGND VGND VPWR VPWR net2722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1761 decode.regfile.registers_17\[9\] VGND VGND VPWR VPWR net1988 sky130_fd_sc_hd__dlygate4sd3_1
X_29533_ clknet_leaf_251_clock _02546_ VGND VGND VPWR VPWR decode.regfile.registers_9\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23957_ net917 execute.io_target_pc\[0\] _07983_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__mux2_1
X_26745_ _09424_ _09733_ VGND VGND VPWR VPWR _09739_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1772 decode.id_ex_rs1_data_reg\[6\] VGND VGND VPWR VPWR net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1783 fetch.bht.bhtTable_target_pc\[9\]\[31\] VGND VGND VPWR VPWR net2010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ net1637 _10027_ _10059_ _10020_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__o211a_1
Xhold1794 decode.regfile.registers_24\[3\] VGND VGND VPWR VPWR net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22908_ _06671_ _07356_ _07357_ _07358_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__and4b_1
X_14690_ decode.id_ex_pc_reg\[31\] VGND VGND VPWR VPWR _10733_ sky130_fd_sc_hd__inv_2
X_26676_ net2577 _09692_ _09698_ _09688_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29464_ clknet_leaf_249_clock _02477_ VGND VGND VPWR VPWR decode.regfile.registers_6\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_23888_ execute.io_target_pc\[31\] VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28415_ clknet_leaf_39_clock _01428_ VGND VGND VPWR VPWR decode.control.io_opcode\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_13641_ _09999_ _09951_ VGND VGND VPWR VPWR _10000_ sky130_fd_sc_hd__nand2_1
X_22839_ _07315_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25627_ net849 _09068_ _09081_ _09074_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29395_ clknet_leaf_258_clock _02408_ VGND VGND VPWR VPWR decode.regfile.registers_4\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16360_ decode.regfile.registers_14\[27\] _11360_ _11274_ decode.regfile.registers_15\[27\]
+ _11361_ VGND VGND VPWR VPWR _12330_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_15_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28346_ clknet_leaf_194_clock _01359_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25558_ _08933_ _09036_ VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__nand2_1
X_13572_ _09936_ VGND VGND VPWR VPWR _09937_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15311_ _10627_ decode.immGen._imm_T_24\[11\] _11091_ _11056_ VGND VGND VPWR VPWR
+ _11307_ sky130_fd_sc_hd__and4_2
XFILLER_0_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24509_ _08435_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__clkbuf_1
X_28277_ clknet_leaf_59_clock _01299_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_16291_ decode.regfile.registers_21\[25\] _11060_ _11098_ _11227_ _12262_ VGND VGND
+ VPWR VPWR _12263_ sky130_fd_sc_hd__o311a_1
XFILLER_0_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25489_ net2397 _08995_ _09001_ _08991_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_183_Left_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18030_ decode.regfile.registers_13\[31\] _12927_ _12588_ _03424_ _03425_ VGND VGND
+ VPWR VPWR _03426_ sky130_fd_sc_hd__a32o_1
X_15242_ decode.regfile.registers_26\[0\] _11236_ _11237_ decode.regfile.registers_27\[0\]
+ _11238_ VGND VGND VPWR VPWR _11239_ sky130_fd_sc_hd__o221a_1
X_27228_ clknet_leaf_4_clock _00257_ VGND VGND VPWR VPWR decode.regfile.registers_29\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27159_ clknet_leaf_356_clock _00188_ VGND VGND VPWR VPWR decode.regfile.registers_27\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15173_ _11169_ VGND VGND VPWR VPWR _11170_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14124_ net1709 _10288_ _10329_ _10328_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__o211a_1
X_19981_ _05218_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14055_ net897 _10287_ _10289_ _10291_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__o211a_1
X_18932_ _03670_ net261 _04230_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18863_ net308 _04158_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_201_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_192_Left_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17814_ _12712_ decode.regfile.registers_24\[25\] _12997_ _12998_ _13367_ VGND VGND
+ VPWR VPWR _03216_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_59_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18794_ decode.id_ex_rs2_data_reg\[15\] net199 _04087_ _04046_ _04092_ VGND VGND
+ VPWR VPWR _04093_ sky130_fd_sc_hd__o221a_1
XFILLER_0_98_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17745_ decode.regfile.registers_20\[24\] _12525_ _12552_ _12823_ _12824_ VGND VGND
+ VPWR VPWR _03148_ sky130_fd_sc_hd__a41o_1
X_14957_ decode.immGen._imm_T_10\[2\] _10667_ _10975_ _10657_ VGND VGND VPWR VPWR
+ _10984_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_193_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13908_ _09984_ _10200_ VGND VGND VPWR VPWR _10205_ sky130_fd_sc_hd__nand2_1
X_17676_ _03078_ _03079_ _03080_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14888_ _10924_ VGND VGND VPWR VPWR _10925_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19415_ _04334_ net278 VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16627_ decode.immGen._imm_T_24\[17\] _10605_ VGND VGND VPWR VPWR _12592_ sky130_fd_sc_hd__nor2_4
X_13839_ _10152_ VGND VGND VPWR VPWR _10164_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19346_ _04582_ _04172_ _04075_ _04227_ _04174_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_58_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16558_ _12522_ VGND VGND VPWR VPWR _12523_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15509_ decode.regfile.registers_3\[5\] _11292_ _11293_ _10635_ VGND VGND VPWR VPWR
+ _11501_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_57_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19277_ _04243_ _04570_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16489_ decode.regfile.registers_13\[31\] _11276_ _11407_ decode.regfile.registers_12\[31\]
+ VGND VGND VPWR VPWR _12455_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18228_ csr.mcycle\[20\] _03554_ _03555_ _03562_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18159_ _03463_ _03464_ _03465_ _10662_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_14_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold302 decode.regfile.registers_17\[11\] VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold313 decode.regfile.registers_20\[10\] VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold324 decode.regfile.registers_9\[10\] VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_229_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21170_ _06079_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__clkbuf_1
Xhold335 decode.regfile.registers_12\[1\] VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_229_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold346 decode.regfile.registers_28\[0\] VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 csr.minstret\[27\] VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20121_ _05329_ _05330_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold368 decode.regfile.registers_19\[15\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold379 csr.minstret\[10\] VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20052_ _05261_ _05268_ _05271_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_225_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 fetch.bht.bhtTable_target_pc\[14\]\[14\] VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__dlygate4sd3_1
X_24860_ _06138_ net1893 _08388_ VGND VGND VPWR VPWR _08618_ sky130_fd_sc_hd__mux2_1
Xhold1013 fetch.bht.bhtTable_tag\[3\]\[9\] VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 csr.mscratch\[30\] VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 fetch.bht.bhtTable_target_pc\[2\]\[8\] VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1046 fetch.bht.bhtTable_tag\[10\]\[19\] VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__dlygate4sd3_1
X_23811_ _08061_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__clkbuf_1
Xhold1057 fetch.bht.bhtTable_tag\[1\]\[9\] VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24791_ _08085_ net1880 _08574_ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1068 decode.regfile.registers_26\[1\] VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1079 decode.regfile.registers_23\[1\] VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26530_ net2424 _09605_ _09614_ _09608_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__o211a_1
X_23742_ _08022_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20954_ _05958_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26461_ net1054 _09535_ _09574_ _09567_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_81_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _07985_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_81_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20885_ _09955_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28200_ clknet_leaf_63_clock net1914 VGND VGND VPWR VPWR csr.mscratch\[2\] sky130_fd_sc_hd__dfxtp_1
X_25412_ net198 VGND VGND VPWR VPWR _08952_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22624_ csr._minstret_T_3\[56\] csr._minstret_T_3\[55\] _07190_ _07148_ VGND VGND
+ VPWR VPWR _07193_ sky130_fd_sc_hd__a31o_1
X_29180_ clknet_leaf_157_clock _02193_ VGND VGND VPWR VPWR fetch.btb.btbTable\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26392_ _10245_ _09535_ VGND VGND VPWR VPWR _09536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28131_ clknet_leaf_236_clock _01153_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25343_ _08902_ VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__buf_2
XFILLER_0_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22555_ _06377_ _07142_ _07144_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__nor3_1
XFILLER_0_180_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21506_ _06270_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__clkbuf_1
X_28062_ clknet_leaf_195_clock _01084_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25274_ _08113_ net2010 _09906_ VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22486_ _07080_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27013_ clknet_leaf_342_clock _00042_ VGND VGND VPWR VPWR decode.regfile.registers_22\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_40_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24225_ _08053_ net1867 _06241_ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21437_ _06128_ net1882 _06230_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24156_ _08251_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__clkbuf_1
X_21368_ _06196_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23107_ _07541_ _07085_ _07547_ VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__a21oi_2
X_20319_ _10864_ _05482_ _10786_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__a21oi_1
X_28964_ clknet_leaf_128_clock _01977_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24087_ net1308 execute.io_target_pc\[31\] _07991_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__mux2_1
Xhold880 _08513_ VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__dlygate4sd3_1
X_21299_ _06159_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold891 fetch.bht.bhtTable_target_pc\[11\]\[10\] VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__dlygate4sd3_1
X_23038_ _07475_ _07479_ _07097_ _07482_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__o22a_2
X_27915_ clknet_leaf_69_clock _00944_ VGND VGND VPWR VPWR csr.io_csr_write_address\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28895_ clknet_leaf_182_clock _01908_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15860_ decode.regfile.registers_1\[14\] _11539_ VGND VGND VPWR VPWR _11843_ sky130_fd_sc_hd__nand2_1
X_27846_ clknet_leaf_320_clock _00875_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2270 decode.regfile.registers_19\[0\] VGND VGND VPWR VPWR net2497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14811_ decode.id_ex_pc_reg\[27\] VGND VGND VPWR VPWR _10854_ sky130_fd_sc_hd__clkbuf_4
Xhold2281 decode.regfile.registers_8\[21\] VGND VGND VPWR VPWR net2508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2292 decode.regfile.registers_11\[22\] VGND VGND VPWR VPWR net2519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15791_ _11058_ _10632_ _10640_ _11071_ _11775_ VGND VGND VPWR VPWR _11776_ sky130_fd_sc_hd__a41o_1
X_27777_ clknet_leaf_328_clock _00806_ VGND VGND VPWR VPWR memory.io_wb_readdata\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_24989_ net512 _08704_ _08705_ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__a21oi_1
Xhold1580 fetch.bht.bhtTable_target_pc\[13\]\[15\] VGND VGND VPWR VPWR net1807 sky130_fd_sc_hd__dlygate4sd3_1
X_17530_ decode.regfile.registers_20\[18\] _12770_ _13475_ _13476_ _12537_ VGND VGND
+ VPWR VPWR _13477_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29516_ clknet_leaf_265_clock _02529_ VGND VGND VPWR VPWR decode.regfile.registers_8\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1591 fetch.bht.bhtTable_target_pc\[11\]\[25\] VGND VGND VPWR VPWR net1818 sky130_fd_sc_hd__dlygate4sd3_1
X_14742_ _10697_ _10776_ _10783_ _10784_ VGND VGND VPWR VPWR _10785_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_153_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26728_ _09406_ _09720_ VGND VGND VPWR VPWR _09729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14673_ decode.id_ex_pc_reg\[20\] VGND VGND VPWR VPWR _10716_ sky130_fd_sc_hd__inv_2
X_17461_ _13183_ _13406_ _13408_ _13409_ VGND VGND VPWR VPWR _13410_ sky130_fd_sc_hd__a31o_1
X_29447_ clknet_leaf_269_clock _02460_ VGND VGND VPWR VPWR decode.regfile.registers_6\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26659_ _09664_ VGND VGND VPWR VPWR _09689_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_103_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19200_ net212 VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_103_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13624_ _09984_ _09951_ VGND VGND VPWR VPWR _09985_ sky130_fd_sc_hd__nand2_1
X_16412_ _10961_ _11834_ _11944_ decode.regfile.registers_29\[28\] _12380_ VGND VGND
+ VPWR VPWR _12381_ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17392_ decode.regfile.registers_4\[15\] _12618_ _12620_ decode.regfile.registers_5\[15\]
+ _12622_ VGND VGND VPWR VPWR _13342_ sky130_fd_sc_hd__a221o_1
X_29378_ clknet_leaf_256_clock _02391_ VGND VGND VPWR VPWR decode.regfile.registers_4\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19131_ _04392_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28329_ clknet_leaf_170_clock _01342_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_13555_ net100 net111 net132 execute.io_mem_memwrite VGND VGND VPWR VPWR _09922_
+ sky130_fd_sc_hd__o22a_1
X_16343_ decode.regfile.registers_17\[27\] _11356_ VGND VGND VPWR VPWR _12313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19062_ _04242_ _04359_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__nand2_4
X_16274_ net343 decode.regfile.registers_3\[25\] _11121_ _11178_ _11367_ VGND VGND
+ VPWR VPWR _12246_ sky130_fd_sc_hd__o32a_1
XFILLER_0_82_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15225_ _11221_ VGND VGND VPWR VPWR _11222_ sky130_fd_sc_hd__clkbuf_4
X_18013_ _12765_ net498 _12486_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15156_ _11107_ _10623_ _11055_ decode.immGen._imm_T_24\[11\] VGND VGND VPWR VPWR
+ _11153_ sky130_fd_sc_hd__nand4_4
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14107_ net2467 _10315_ _10320_ _10317_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19964_ net1630 _03599_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__nor2_1
X_15087_ _11083_ VGND VGND VPWR VPWR _11084_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_1196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14038_ _10122_ _10268_ VGND VGND VPWR VPWR _10280_ sky130_fd_sc_hd__nand2_1
X_18915_ _04175_ _04188_ _03867_ _04213_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__a211o_1
X_19895_ _03790_ _05162_ _03865_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18846_ memory.csr_read_data_out_reg\[11\] _10010_ _10033_ _10034_ VGND VGND VPWR
+ VPWR _04145_ sky130_fd_sc_hd__o22a_2
XFILLER_0_101_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_220_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18777_ _04045_ _04049_ _04062_ _04065_ _04075_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__o221a_1
XFILLER_0_175_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15989_ decode.regfile.registers_17\[17\] _11094_ _11114_ _11119_ _11968_ VGND VGND
+ VPWR VPWR _11969_ sky130_fd_sc_hd__a41o_1
XFILLER_0_37_1310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17728_ decode.regfile.registers_16\[23\] _13011_ _03114_ _03131_ _12579_ VGND VGND
+ VPWR VPWR _03132_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17659_ _13407_ decode.regfile.registers_25\[21\] _13482_ _13294_ VGND VGND VPWR
+ VPWR _03065_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_154_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20670_ _05795_ _05792_ _05796_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19329_ _04065_ _04062_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__or2b_1
XFILLER_0_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22340_ _06730_ _06934_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_171_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22271_ _06651_ _06865_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24010_ _08176_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_227_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21222_ _10817_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_115_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_148_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold154 io_fetch_data[0] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold165 fetch.bht.bhtTable_valid\[2\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21153_ _09955_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_180_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold176 execute.csr_write_address_out_reg\[7\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_180_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold187 fetch.btb.btbTable\[10\]\[0\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 fetch.btb.btbTable\[4\]\[0\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
X_20104_ _05314_ _05315_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25961_ _08958_ _09267_ VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_70_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21084_ execute.csr_read_data_out_reg\[30\] _06025_ _03583_ VGND VGND VPWR VPWR _06029_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_10_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27700_ clknet_leaf_24_clock _00729_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20035_ _05254_ _05255_ _05256_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__a21oi_1
X_24912_ net2057 _08654_ _08655_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28680_ clknet_leaf_96_clock _01693_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25892_ net2521 _09226_ _09233_ _09222_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27631_ clknet_leaf_44_clock _00660_ VGND VGND VPWR VPWR execute.io_reg_pc\[8\] sky130_fd_sc_hd__dfxtp_1
X_24843_ _08609_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_11 _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_22 _03142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_33 _08929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_44 _09932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24774_ _08068_ net991 _08563_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_178_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27562_ clknet_leaf_157_clock _00591_ VGND VGND VPWR VPWR csr.io_mem_pc\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_178_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ csr._mcycle_T_2\[16\] _06587_ _06596_ _06592_ VGND VGND VPWR VPWR _01236_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_55 _10073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_66 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_217_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29301_ clknet_leaf_225_clock _02314_ VGND VGND VPWR VPWR decode.regfile.registers_1\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_77 _10240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23725_ _08013_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__clkbuf_1
X_26513_ _09577_ VGND VGND VPWR VPWR _09605_ sky130_fd_sc_hd__buf_2
XINSDIODE1_88 _10594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_99 _10655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20937_ _05949_ _05945_ net53 VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27493_ clknet_leaf_27_clock _00522_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dfxtp_1
X_29232_ clknet_leaf_122_clock _02245_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23656_ _07976_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26444_ _09426_ _09558_ VGND VGND VPWR VPWR _09565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20868_ net120 _05903_ _05911_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22607_ csr._minstret_T_3\[50\] csr._minstret_T_3\[49\] _07178_ _06422_ VGND VGND
+ VPWR VPWR _07182_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_42_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29163_ clknet_leaf_195_clock _02176_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_26375_ net2683 _09518_ _09524_ _09525_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23587_ _07938_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20799_ execute.io_mem_regwrite _05867_ _05868_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28114_ clknet_leaf_81_clock _01136_ VGND VGND VPWR VPWR csr.minstret\[19\] sky130_fd_sc_hd__dfxtp_2
X_25326_ _08891_ net2666 VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22538_ _07129_ _07091_ net280 _07131_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__o31a_1
XFILLER_0_10_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29094_ clknet_leaf_70_clock _02107_ VGND VGND VPWR VPWR csr._mcycle_T_3\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25257_ _08858_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__clkbuf_1
X_28045_ clknet_leaf_222_clock _01067_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22469_ _07063_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15010_ _11019_ VGND VGND VPWR VPWR _11020_ sky130_fd_sc_hd__clkbuf_4
X_24208_ _08278_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25188_ _10572_ fetch.btb.btbTable\[5\]\[1\] _08822_ VGND VGND VPWR VPWR _08823_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24139_ net1001 execute.io_target_pc\[24\] _06427_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28947_ clknet_leaf_140_clock _01960_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16961_ _12765_ _12768_ _12493_ decode.regfile.registers_29\[4\] _12921_ VGND VGND
+ VPWR VPWR _12922_ sky130_fd_sc_hd__o221a_1
XFILLER_0_159_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18700_ _03768_ _03769_ _03770_ _09963_ net234 VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__o311a_1
X_15912_ decode.regfile.registers_11\[15\] _11181_ _11892_ _11893_ _11407_ VGND VGND
+ VPWR VPWR _11894_ sky130_fd_sc_hd__a221o_1
XFILLER_0_200_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19680_ _03956_ _03959_ _04932_ _04192_ _04191_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__a221oi_1
X_28878_ clknet_leaf_111_clock _01891_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_16892_ decode.regfile.registers_15\[3\] _12584_ _12673_ _12853_ VGND VGND VPWR VPWR
+ _12854_ sky130_fd_sc_hd__a211o_1
X_18631_ decode.id_ex_rs2_data_reg\[16\] _03746_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_216_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15843_ _11436_ decode.regfile.registers_26\[13\] _11676_ _11338_ _11564_ VGND VGND
+ VPWR VPWR _11827_ sky130_fd_sc_hd__o2111a_1
X_27829_ clknet_leaf_325_clock _00858_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18562_ _03709_ decode.id_ex_imm_reg\[30\] _03859_ _03860_ VGND VGND VPWR VPWR _03861_
+ sky130_fd_sc_hd__a22oi_4
X_15774_ _11248_ VGND VGND VPWR VPWR _11760_ sky130_fd_sc_hd__buf_2
XFILLER_0_86_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17513_ decode.regfile.registers_4\[18\] _12618_ _12620_ decode.regfile.registers_5\[18\]
+ _12737_ VGND VGND VPWR VPWR _13460_ sky130_fd_sc_hd__a221o_1
X_14725_ csr.io_mem_pc\[22\] csr.io_mem_pc\[23\] _10767_ VGND VGND VPWR VPWR _10768_
+ sky130_fd_sc_hd__and3_4
XFILLER_0_169_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18493_ execute.csr_read_data_out_reg\[28\] _03661_ _03660_ VGND VGND VPWR VPWR _03792_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_129_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17444_ _12540_ _12722_ _12724_ _13391_ _13392_ VGND VGND VPWR VPWR _13393_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_196_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14656_ _10695_ _10696_ _10697_ _10698_ VGND VGND VPWR VPWR _10699_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_5_8__f_clock clknet_2_1_0_clock VGND VGND VPWR VPWR clknet_5_8__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13607_ _09969_ VGND VGND VPWR VPWR _09970_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17375_ _12584_ _13324_ _13325_ VGND VGND VPWR VPWR _13326_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14587_ _10629_ VGND VGND VPWR VPWR _10630_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_188_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19114_ _04275_ _04284_ _04352_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16326_ decode.regfile.registers_19\[26\] _11048_ _11215_ _11217_ _11219_ VGND VGND
+ VPWR VPWR _12297_ sky130_fd_sc_hd__o41a_1
X_13538_ _09913_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19045_ _04281_ _04337_ _04283_ _04244_ _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__o311a_1
XFILLER_0_3_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16257_ _11076_ _11090_ decode.regfile.registers_25\[24\] _12203_ _12229_ VGND VGND
+ VPWR VPWR _12230_ sky130_fd_sc_hd__o32a_1
XFILLER_0_207_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15208_ _11204_ VGND VGND VPWR VPWR _11205_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16188_ decode.regfile.registers_23\[22\] _11087_ _12136_ _12162_ VGND VGND VPWR
+ VPWR _12163_ sky130_fd_sc_hd__o22a_1
XFILLER_0_112_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15139_ _11135_ VGND VGND VPWR VPWR _11136_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_222_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_222_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19947_ _03581_ _05201_ net1983 VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__and3b_1
XFILLER_0_103_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19878_ _03791_ _03803_ _05123_ _05147_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__a31o_1
XFILLER_0_177_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18829_ decode.id_ex_rs2_data_reg\[8\] _03746_ _03764_ _04122_ VGND VGND VPWR VPWR
+ _04128_ sky130_fd_sc_hd__o22a_1
X_21840_ _06491_ _06494_ _06495_ _06498_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21771_ _06448_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23510_ net2024 _07890_ _07887_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__or3b_1
XFILLER_0_114_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20722_ _00514_ _05723_ _05830_ net182 net2730 VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__a32o_1
X_24490_ _08425_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_173_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23441_ net32 _07846_ _07855_ _07851_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20653_ csr.minstret\[30\] _05572_ _05582_ csr.mcycle\[30\] _05782_ VGND VGND VPWR
+ VPWR _05783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_870 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26160_ net2585 _09373_ _09391_ _09370_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__o211a_1
X_23372_ fetch.bht.bhtTable_target_pc\[4\]\[28\] fetch.bht.bhtTable_target_pc\[5\]\[28\]
+ fetch.bht.bhtTable_target_pc\[6\]\[28\] fetch.bht.bhtTable_target_pc\[7\]\[28\]
+ _07384_ _07386_ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__mux4_1
XFILLER_0_190_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20584_ _05724_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25111_ _06128_ net1815 _08778_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22323_ _06691_ fetch.bht.bhtTable_tag\[10\]\[8\] VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_76_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26091_ _08937_ _09340_ VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25042_ _08701_ _03562_ _06327_ _08741_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_132_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22254_ _06642_ _06838_ _06842_ _06848_ net220 VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__o311a_1
XFILLER_0_42_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21205_ decode.id_ex_ex_rd_reg\[0\] _05214_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29850_ clknet_leaf_306_clock _02863_ VGND VGND VPWR VPWR decode.regfile.registers_19\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_22185_ _06624_ _06779_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28801_ clknet_leaf_175_clock _01814_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21136_ _06050_ _06058_ net1404 VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_109_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29781_ clknet_leaf_294_clock _02794_ VGND VGND VPWR VPWR decode.regfile.registers_16\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_26993_ clknet_leaf_334_clock _00022_ VGND VGND VPWR VPWR decode.regfile.registers_22\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28732_ clknet_leaf_185_clock _01745_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_25944_ net1198 _09256_ _09262_ _09264_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__o211a_1
X_21067_ execute.csr_read_data_out_reg\[22\] _06014_ _06010_ VGND VGND VPWR VPWR _06020_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_214_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20018_ _05240_ _05241_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28663_ clknet_leaf_117_clock _01676_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25875_ net2266 _09213_ _09224_ _09222_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__o211a_1
X_27614_ clknet_leaf_150_clock _00643_ VGND VGND VPWR VPWR execute.io_target_pc\[23\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_119_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24826_ _08600_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__clkbuf_1
X_28594_ clknet_leaf_102_clock _01607_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27545_ clknet_leaf_44_clock _00574_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfxtp_4
X_24757_ _08564_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__clkbuf_1
X_21969_ csr._mcycle_T_2\[9\] _06572_ _06586_ _06579_ VGND VGND VPWR VPWR _01229_
+ sky130_fd_sc_hd__o211a_1
XINSDIODE1_309 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14510_ fetch.btb.btbTable\[0\]\[0\] fetch.btb.btbTable\[1\]\[0\] fetch.btb.btbTable\[2\]\[0\]
+ fetch.btb.btbTable\[3\]\[0\] _09891_ _09888_ VGND VGND VPWR VPWR _10555_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_139_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23708_ net1228 _10803_ _08003_ VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _11333_ VGND VGND VPWR VPWR _11483_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24688_ _08527_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27476_ clknet_leaf_53_clock _00505_ VGND VGND VPWR VPWR csr.io_csr_address\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29215_ clknet_leaf_114_clock _02228_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_23639_ _07967_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__clkbuf_1
X_26427_ net1332 _09548_ _09555_ _09553_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_29_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ net429 _10506_ _10513_ _10509_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_360_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_360_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29146_ clknet_leaf_78_clock _02159_ VGND VGND VPWR VPWR csr.mcycle\[30\] sky130_fd_sc_hd__dfxtp_2
X_17160_ _13114_ _13115_ VGND VGND VPWR VPWR _13116_ sky130_fd_sc_hd__nand2_1
X_14372_ net467 _10463_ _10473_ _10468_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26358_ _09412_ _09515_ VGND VGND VPWR VPWR _09516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16111_ _11050_ decode.regfile.registers_25\[20\] _11089_ VGND VGND VPWR VPWR _12088_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_88_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25309_ _08880_ net2694 VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29077_ clknet_leaf_191_clock _02090_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26289_ net2543 _09475_ _09476_ _09471_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__o211a_1
X_17091_ _12695_ _13044_ _13046_ _13048_ VGND VGND VPWR VPWR _13049_ sky130_fd_sc_hd__a31o_1
XFILLER_0_162_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28028_ clknet_leaf_205_clock _01050_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16042_ decode.regfile.registers_7\[19\] _11092_ _11142_ _11166_ VGND VGND VPWR VPWR
+ _12020_ sky130_fd_sc_hd__a31o_1
XFILLER_0_161_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19801_ _04330_ _04984_ _05073_ _04302_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_209_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17993_ decode.regfile.registers_10\[30\] _12599_ _12594_ _03389_ VGND VGND VPWR
+ VPWR _03390_ sky130_fd_sc_hd__a211o_1
X_19732_ _05007_ _04919_ _04269_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__mux2_1
X_16944_ decode.regfile.registers_18\[4\] _12572_ _12903_ _12904_ _12562_ VGND VGND
+ VPWR VPWR _12905_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19663_ _04446_ _04934_ _04940_ _04941_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__o31a_1
X_16875_ _12522_ _10601_ _10591_ VGND VGND VPWR VPWR _12837_ sky130_fd_sc_hd__and3_2
X_18614_ _10072_ _10071_ _09986_ memory.csr_read_data_out_reg\[18\] VGND VGND VPWR
+ VPWR _03913_ sky130_fd_sc_hd__o2bb2a_2
X_15826_ _10647_ _10624_ _11462_ _11802_ _11809_ VGND VGND VPWR VPWR _11810_ sky130_fd_sc_hd__o32a_2
XFILLER_0_56_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_313_clock clknet_5_18__leaf_clock VGND VGND VPWR VPWR clknet_leaf_313_clock
+ sky130_fd_sc_hd__clkbuf_8
X_19594_ _04812_ _04875_ _04277_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18545_ _03656_ _03841_ _03670_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__o211a_4
X_15757_ decode.regfile.registers_13\[11\] _10639_ _11187_ VGND VGND VPWR VPWR _11743_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_172_1287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14708_ _10713_ execute.io_target_pc\[18\] VGND VGND VPWR VPWR _10751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18476_ _03774_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_157_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15688_ _11080_ VGND VGND VPWR VPWR _11676_ sky130_fd_sc_hd__buf_2
XFILLER_0_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_215_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17427_ net438 _12709_ _13338_ _13376_ _13219_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_328_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_328_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14639_ _10681_ VGND VGND VPWR VPWR _10682_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_211_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17358_ decode.regfile.registers_11\[14\] _12594_ _12582_ _12550_ VGND VGND VPWR
+ VPWR _13309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16309_ _11371_ decode.regfile.registers_0\[26\] _11156_ _12279_ VGND VGND VPWR VPWR
+ _12280_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17289_ decode.regfile.registers_16\[12\] _12674_ _12901_ _13241_ VGND VGND VPWR
+ VPWR _13242_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19028_ _03986_ _03985_ _03984_ _03987_ _04062_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__a311o_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23990_ _08166_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_162_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22941_ net186 VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22872_ _07332_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__clkbuf_1
X_25660_ net2328 _09095_ _09099_ _09100_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24611_ net1241 execute.io_target_pc\[27\] _09897_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21823_ _06479_ net559 _06396_ _06485_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_65_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25591_ net2302 _09052_ _09060_ _09059_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24542_ _08452_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_174_Right_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27330_ clknet_leaf_41_clock _00359_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_66_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21754_ net956 _10868_ _06439_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20705_ _05801_ _05808_ decode.id_ex_rs1_data_reg\[12\] _05820_ _00699_ VGND VGND
+ VPWR VPWR _00731_ sky130_fd_sc_hd__a32o_1
X_24473_ _08416_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__clkbuf_1
X_27261_ clknet_leaf_5_clock _00290_ VGND VGND VPWR VPWR decode.regfile.registers_30\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_21685_ csr._mcycle_T_2\[24\] _06329_ _06389_ csr.minstret\[24\] VGND VGND VPWR VPWR
+ _06390_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_163_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29000_ clknet_leaf_103_clock _02013_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23424_ net91 _07706_ _07707_ _07845_ _05856_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_134_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26212_ net197 VGND VGND VPWR VPWR _09428_ sky130_fd_sc_hd__buf_4
X_20636_ csr.mscratch\[27\] _05593_ _05625_ _05767_ _05768_ VGND VGND VPWR VPWR _05769_
+ sky130_fd_sc_hd__o32a_1
X_27192_ clknet_leaf_355_clock _00221_ VGND VGND VPWR VPWR decode.regfile.registers_28\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26143_ _09379_ _09374_ VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__nand2_1
X_23355_ execute.io_target_pc\[27\] _10757_ _10970_ _06037_ VGND VGND VPWR VPWR _07781_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_190_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20567_ _05705_ _05707_ _05709_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22306_ fetch.bht.bhtTable_tag\[7\]\[0\] _06674_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26074_ _08920_ _09330_ VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_95_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23286_ net223 _07716_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20498_ _05556_ csr._minstret_T_3\[40\] _05647_ _05649_ VGND VGND VPWR VPWR _05650_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25025_ _08729_ _08727_ _06327_ _08730_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__a211oi_1
X_29902_ clknet_leaf_301_clock _02915_ VGND VGND VPWR VPWR decode.regfile.registers_20\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_22237_ _06831_ _06628_ _06635_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29833_ clknet_leaf_298_clock _02846_ VGND VGND VPWR VPWR decode.regfile.registers_18\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_22168_ fetch.bht.bhtTable_tag\[14\]\[13\] fetch.bht.bhtTable_tag\[15\]\[13\] _06644_
+ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__mux2_1
X_21119_ _06050_ _06046_ net1785 VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29764_ clknet_leaf_293_clock _02777_ VGND VGND VPWR VPWR decode.regfile.registers_16\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_22099_ fetch.bht.bhtTable_tag\[14\]\[7\] fetch.bht.bhtTable_tag\[15\]\[7\] _06680_
+ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__mux2_1
X_14990_ _10948_ _10950_ _10952_ _10998_ decode.control.io_funct7\[6\] VGND VGND VPWR
+ VPWR _11007_ sky130_fd_sc_hd__o311a_2
XFILLER_0_22_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26976_ net2309 _09866_ _09871_ _09865_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_54_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28715_ clknet_leaf_95_clock _01728_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13941_ _10074_ _10223_ VGND VGND VPWR VPWR _10224_ sky130_fd_sc_hd__nand2_1
X_25927_ net730 _09242_ _09254_ _09250_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__o211a_1
X_29695_ clknet_leaf_289_clock _02708_ VGND VGND VPWR VPWR decode.regfile.registers_14\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28646_ clknet_leaf_96_clock _01659_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16660_ _12613_ VGND VGND VPWR VPWR _12625_ sky130_fd_sc_hd__clkbuf_4
X_13872_ _10097_ _10177_ VGND VGND VPWR VPWR _10183_ sky130_fd_sc_hd__nand2_1
X_25858_ _08931_ _09210_ VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15611_ decode.regfile.registers_23\[7\] _11087_ _11573_ _11600_ VGND VGND VPWR VPWR
+ _11601_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24809_ _08591_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28577_ clknet_leaf_185_clock _01590_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_16591_ _10597_ decode.immGen._imm_T_24\[17\] VGND VGND VPWR VPWR _12556_ sky130_fd_sc_hd__nor2_1
X_25789_ _08937_ _09166_ VGND VGND VPWR VPWR _09175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_106 _10935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_26__f_clock clknet_2_3_0_clock VGND VGND VPWR VPWR clknet_5_26__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_117 _11054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18330_ decode.id_ex_rs2_data_reg\[30\] _03627_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27528_ clknet_leaf_44_clock _00557_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_128 _11192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15542_ _11503_ _10624_ _11043_ _11083_ VGND VGND VPWR VPWR _11533_ sky130_fd_sc_hd__or4_2
XFILLER_0_167_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_139 _12377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18261_ _03591_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27459_ clknet_leaf_137_clock _00488_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15473_ _11169_ VGND VGND VPWR VPWR _11466_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_194_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17212_ decode.regfile.registers_22\[10\] _12528_ _13166_ _12687_ VGND VGND VPWR
+ VPWR _13167_ sky130_fd_sc_hd__a211o_1
X_14424_ net1571 _10464_ _10502_ _10494_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__o211a_1
X_18192_ decode.control.io_funct7\[6\] _03529_ decode.control.io_funct7\[5\] decode.control.io_funct7\[3\]
+ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__or4b_1
XFILLER_0_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29129_ clknet_leaf_76_clock _02142_ VGND VGND VPWR VPWR csr.mcycle\[13\] sky130_fd_sc_hd__dfxtp_2
X_17143_ _10930_ VGND VGND VPWR VPWR _13099_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14355_ _10462_ VGND VGND VPWR VPWR _10464_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17074_ decode.regfile.registers_15\[7\] _12584_ _13031_ VGND VGND VPWR VPWR _13032_
+ sky130_fd_sc_hd__a21oi_1
X_14286_ _09975_ _10420_ VGND VGND VPWR VPWR _10424_ sky130_fd_sc_hd__nand2_1
Xhold709 decode.regfile.registers_30\[20\] VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16025_ _10955_ _11215_ _11216_ _12003_ VGND VGND VPWR VPWR _12004_ sky130_fd_sc_hd__o31a_1
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17976_ _12708_ net445 _03336_ _03373_ _03073_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__o221a_1
Xhold1409 fetch.bht.bhtTable_tag\[12\]\[25\] VGND VGND VPWR VPWR net1636 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_204_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19715_ _03868_ _03701_ _03689_ decode.id_ex_rs1_data_reg\[23\] _03871_ VGND VGND
+ VPWR VPWR _04991_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_204_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16927_ _12843_ VGND VGND VPWR VPWR _12888_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_252_clock clknet_5_18__leaf_clock VGND VGND VPWR VPWR clknet_leaf_252_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19646_ _04922_ _04923_ _04925_ _04515_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__and4_1
X_16858_ net801 _12709_ _12764_ _12820_ _12705_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__o221a_1
XFILLER_0_215_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_217_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15809_ _11489_ decode.regfile.registers_28\[12\] decode.regfile.registers_29\[12\]
+ _11255_ _11246_ VGND VGND VPWR VPWR _11794_ sky130_fd_sc_hd__o221a_1
X_19577_ _03639_ _04620_ _04197_ _04858_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__o22a_1
XFILLER_0_215_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16789_ decode.regfile.registers_17\[1\] _12719_ _12565_ _12752_ VGND VGND VPWR VPWR
+ _12753_ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18528_ net188 _03825_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_267_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_267_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18459_ _03751_ _03752_ _03757_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__nand3_4
XFILLER_0_29_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21470_ _06250_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20421_ _03721_ _05554_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23140_ fetch.bht.bhtTable_target_pc\[12\]\[14\] fetch.bht.bhtTable_target_pc\[13\]\[14\]
+ fetch.bht.bhtTable_target_pc\[14\]\[14\] fetch.bht.bhtTable_target_pc\[15\]\[14\]
+ _07069_ _07111_ VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_168_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20352_ _05513_ _05515_ _05410_ _05412_ _03588_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_168_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23071_ fetch.bht.bhtTable_target_pc\[8\]\[10\] fetch.bht.bhtTable_target_pc\[9\]\[10\]
+ _07119_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_205_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_205_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20283_ _05417_ _05313_ _05463_ _05454_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22022_ _06616_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_90_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26830_ net2619 _09779_ _09787_ _09784_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1910 fetch.bht.bhtTable_target_pc\[0\]\[10\] VGND VGND VPWR VPWR net2137 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1921 decode.regfile.registers_13\[18\] VGND VGND VPWR VPWR net2148 sky130_fd_sc_hd__dlygate4sd3_1
X_26761_ net2682 _09736_ _09747_ _09743_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__o211a_1
Xhold1932 _01248_ VGND VGND VPWR VPWR net2159 sky130_fd_sc_hd__dlygate4sd3_1
X_23973_ _08157_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1943 decode.regfile.registers_11\[1\] VGND VGND VPWR VPWR net2170 sky130_fd_sc_hd__dlygate4sd3_1
X_28500_ clknet_leaf_214_clock _01513_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_123_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1954 decode.id_ex_ex_rd_reg\[3\] VGND VGND VPWR VPWR net2181 sky130_fd_sc_hd__buf_1
XFILLER_0_98_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1965 decode.regfile.registers_9\[8\] VGND VGND VPWR VPWR net2192 sky130_fd_sc_hd__dlygate4sd3_1
X_25712_ _08935_ _09122_ VGND VGND VPWR VPWR _09131_ sky130_fd_sc_hd__nand2_1
X_22924_ fetch.bht.bhtTable_target_pc\[14\]\[2\] fetch.bht.bhtTable_target_pc\[15\]\[2\]
+ _07119_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29480_ clknet_leaf_254_clock _02493_ VGND VGND VPWR VPWR decode.regfile.registers_7\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_123_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1976 decode.regfile.registers_15\[31\] VGND VGND VPWR VPWR net2203 sky130_fd_sc_hd__dlygate4sd3_1
X_26692_ _09707_ VGND VGND VPWR VPWR _09708_ sky130_fd_sc_hd__clkbuf_4
Xhold1987 decode.regfile.registers_12\[12\] VGND VGND VPWR VPWR net2214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1998 fetch.bht.bhtTable_tag\[13\]\[16\] VGND VGND VPWR VPWR net2225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28431_ clknet_leaf_246_clock _01444_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[1\]
+ sky130_fd_sc_hd__dfxtp_4
X_25643_ net1133 _09082_ _09090_ _09087_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__o211a_1
X_22855_ _07323_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28362_ clknet_leaf_238_clock _01375_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_21806_ net2613 _06471_ _06473_ _10546_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__o211a_1
X_22786_ net1474 _10821_ _07286_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__mux2_1
X_25574_ _08948_ _09049_ VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27313_ clknet_leaf_34_clock _00342_ VGND VGND VPWR VPWR decode.id_ex_ex_use_rs1_reg
+ sky130_fd_sc_hd__dfxtp_1
X_24525_ _08085_ net1832 _08439_ VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21737_ net2000 _10881_ _06428_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__mux2_1
X_28293_ clknet_leaf_60_clock _01315_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27244_ clknet_leaf_2_clock _00273_ VGND VGND VPWR VPWR decode.regfile.registers_29\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24456_ _08407_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__clkbuf_1
X_21668_ _03579_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_97_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23407_ net90 _07706_ _07707_ _07829_ _07705_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__o311a_1
X_20619_ csr.mscratch\[25\] _05592_ _05611_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__or3_1
XFILLER_0_123_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24387_ net1219 execute.io_target_pc\[16\] _08367_ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__mux2_1
X_27175_ clknet_leaf_362_clock _00204_ VGND VGND VPWR VPWR decode.regfile.registers_27\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_21599_ _10576_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_10_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14140_ net460 _10332_ _10339_ _10328_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23338_ fetch.bht.bhtTable_target_pc\[4\]\[26\] fetch.bht.bhtTable_target_pc\[5\]\[26\]
+ fetch.bht.bhtTable_target_pc\[6\]\[26\] fetch.bht.bhtTable_target_pc\[7\]\[26\]
+ _07669_ _07656_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26126_ _08973_ _09328_ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14071_ _10015_ _10299_ VGND VGND VPWR VPWR _10300_ sky130_fd_sc_hd__nand2_1
X_23269_ _07692_ _07697_ _07127_ _07700_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__a2bb2o_1
X_26057_ _09328_ VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_56_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25008_ _08701_ _03558_ csr.mcycle\[6\] csr.mcycle\[7\] VGND VGND VPWR VPWR _08719_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29816_ clknet_leaf_313_clock _02829_ VGND VGND VPWR VPWR decode.regfile.registers_17\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17830_ decode.regfile.registers_4\[26\] _12618_ _12620_ decode.regfile.registers_5\[26\]
+ _12737_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__a221o_1
XFILLER_0_218_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_210_Right_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29747_ clknet_leaf_284_clock _02760_ VGND VGND VPWR VPWR decode.regfile.registers_15\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_17761_ decode.regfile.registers_11\[24\] _12595_ _03162_ _03163_ _12794_ VGND VGND
+ VPWR VPWR _03164_ sky130_fd_sc_hd__a221o_1
X_14973_ _10967_ VGND VGND VPWR VPWR _10997_ sky130_fd_sc_hd__clkbuf_4
X_26959_ net1222 _09853_ _09861_ _09852_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19500_ _03708_ decode.id_ex_imm_reg\[13\] _04101_ _04102_ _04100_ VGND VGND VPWR
+ VPWR _04785_ sky130_fd_sc_hd__a221o_2
X_16712_ _10598_ _10588_ _12666_ _10594_ VGND VGND VPWR VPWR _12677_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13924_ net904 _10213_ _10214_ _10206_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17692_ decode.regfile.registers_20\[22\] _12771_ _03096_ _12537_ VGND VGND VPWR
+ VPWR _03097_ sky130_fd_sc_hd__a211o_1
X_29678_ clknet_leaf_283_clock _02691_ VGND VGND VPWR VPWR decode.regfile.registers_13\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19431_ _04130_ _04131_ _04142_ _04143_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__o22a_1
X_28629_ clknet_leaf_116_clock _01642_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_16643_ decode.regfile.registers_8\[0\] _10594_ _12550_ _12604_ _12607_ VGND VGND
+ VPWR VPWR _12608_ sky130_fd_sc_hd__a41o_1
XFILLER_0_201_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13855_ _10058_ _10164_ VGND VGND VPWR VPWR _10173_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19362_ _04273_ _04278_ _04288_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__a21oi_1
X_16574_ _10608_ _12508_ VGND VGND VPWR VPWR _12539_ sky130_fd_sc_hd__or2_4
X_13786_ net2482 _10083_ _10123_ _10077_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_191_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18313_ decode.id_ex_rs2_data_reg\[22\] _03616_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15525_ decode.regfile.registers_18\[5\] _11268_ _11271_ _11516_ VGND VGND VPWR VPWR
+ _11517_ sky130_fd_sc_hd__a211o_1
X_19293_ _04075_ _04172_ _04585_ _04553_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18244_ _10575_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__buf_4
XFILLER_0_72_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15456_ _11446_ decode.regfile.registers_26\[4\] _11447_ _10981_ _11448_ VGND VGND
+ VPWR VPWR _11449_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_154_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14407_ _10426_ VGND VGND VPWR VPWR _10494_ sky130_fd_sc_hd__clkbuf_4
X_18175_ _03515_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15387_ _11381_ VGND VGND VPWR VPWR _11382_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17126_ _12690_ VGND VGND VPWR VPWR _13083_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_150_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14338_ _10112_ _10444_ VGND VGND VPWR VPWR _10454_ sky130_fd_sc_hd__nand2_1
Xmax_cap203 net204 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_4
Xmax_cap214 _03521_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_1
Xhold506 decode.regfile.registers_18\[5\] VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold517 decode.regfile.registers_26\[7\] VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_1342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold528 decode.regfile.registers_3\[16\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17057_ decode.regfile.registers_1\[7\] _12631_ _12933_ _12508_ _13014_ VGND VGND
+ VPWR VPWR _13015_ sky130_fd_sc_hd__o221a_1
Xhold539 decode.regfile.registers_13\[3\] VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14269_ net1421 _10403_ _10413_ _10411_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16008_ decode.regfile.registers_11\[18\] _11180_ _11509_ decode.regfile.registers_10\[18\]
+ _11186_ VGND VGND VPWR VPWR _11987_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_206_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_191_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_191_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1206 fetch.bht.bhtTable_target_pc\[2\]\[27\] VGND VGND VPWR VPWR net1433 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 fetch.bht.bhtTable_tag\[6\]\[17\] VGND VGND VPWR VPWR net1444 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 decode.regfile.registers_2\[10\] VGND VGND VPWR VPWR net1455 sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ _11020_ _12491_ _12650_ decode.regfile.registers_14\[29\] _12669_ VGND VGND
+ VPWR VPWR _03357_ sky130_fd_sc_hd__o32a_1
Xhold1239 fetch.bht.bhtTable_target_pc\[12\]\[29\] VGND VGND VPWR VPWR net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_213_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20970_ _05967_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19629_ _03638_ _04207_ _04887_ _04899_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_177_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22640_ csr._minstret_T_3\[61\] _07202_ _07203_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_157_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22571_ csr.minstret\[27\] VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24310_ _08072_ net2336 _08323_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__mux2_1
X_21522_ _06151_ net1313 _06274_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25290_ _08875_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24241_ _08295_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_21_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21453_ _06242_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20404_ _05522_ _03755_ _03741_ _03737_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_116_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24172_ _08066_ net1452 _08255_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21384_ _06132_ net1600 _06199_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_144_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_144_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23123_ _07071_ _07562_ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20335_ _10854_ _05500_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28980_ clknet_leaf_118_clock _01993_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_187_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27931_ clknet_leaf_162_clock _00008_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_23054_ net97 net96 net227 _07427_ _06718_ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__a41o_1
X_20266_ _05417_ _05287_ _05450_ _05414_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22005_ net2142 _06600_ _06607_ _06605_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27862_ clknet_leaf_325_clock _00891_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_159_clock clknet_5_24__leaf_clock VGND VGND VPWR VPWR clknet_leaf_159_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20197_ _05385_ _05392_ _05395_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_51_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29601_ clknet_leaf_271_clock _02614_ VGND VGND VPWR VPWR decode.regfile.registers_11\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2430 execute.csr_write_data_out_reg\[31\] VGND VGND VPWR VPWR net2657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2441 decode.regfile.registers_2\[28\] VGND VGND VPWR VPWR net2668 sky130_fd_sc_hd__dlygate4sd3_1
X_26813_ _09415_ _09776_ VGND VGND VPWR VPWR _09778_ sky130_fd_sc_hd__nand2_1
Xhold2452 csr.minstret\[29\] VGND VGND VPWR VPWR net2679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2463 fetch.btb.btbTable\[7\]\[1\] VGND VGND VPWR VPWR net2690 sky130_fd_sc_hd__dlygate4sd3_1
X_27793_ clknet_leaf_305_clock _00822_ VGND VGND VPWR VPWR memory.io_wb_readdata\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2474 decode.regfile.registers_0\[10\] VGND VGND VPWR VPWR net2701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1740 fetch.bht.bhtTable_target_pc\[0\]\[23\] VGND VGND VPWR VPWR net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2485 csr._minstret_T_3\[41\] VGND VGND VPWR VPWR net2712 sky130_fd_sc_hd__dlygate4sd3_1
X_29532_ clknet_leaf_314_clock _02545_ VGND VGND VPWR VPWR decode.regfile.registers_9\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1751 csr._minstret_T_3\[48\] VGND VGND VPWR VPWR net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2496 decode.regfile.registers_27\[29\] VGND VGND VPWR VPWR net2723 sky130_fd_sc_hd__dlygate4sd3_1
X_26744_ net2282 _09736_ _09738_ _09730_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23956_ _08148_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__clkbuf_1
Xhold1762 fetch.bht.bhtTable_target_pc\[5\]\[9\] VGND VGND VPWR VPWR net1989 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_86_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1773 fetch.bht.bhtTable_tag\[4\]\[2\] VGND VGND VPWR VPWR net2000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1784 fetch.bht.bhtTable_target_pc\[7\]\[14\] VGND VGND VPWR VPWR net2011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1795 fetch.bht.bhtTable_tag\[9\]\[20\] VGND VGND VPWR VPWR net2022 sky130_fd_sc_hd__dlygate4sd3_1
X_22907_ net68 _06739_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__or2_1
X_29463_ clknet_leaf_254_clock _02476_ VGND VGND VPWR VPWR decode.regfile.registers_6\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_26675_ _09430_ _09689_ VGND VGND VPWR VPWR _09698_ sky130_fd_sc_hd__nand2_1
X_23887_ _08112_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28414_ clknet_leaf_54_clock _01427_ VGND VGND VPWR VPWR decode.control.io_opcode\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_13640_ _09998_ VGND VGND VPWR VPWR _09999_ sky130_fd_sc_hd__buf_4
X_25626_ _08925_ _09079_ VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22838_ net1396 _10820_ _09898_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__mux2_1
X_29394_ clknet_leaf_258_clock _02407_ VGND VGND VPWR VPWR decode.regfile.registers_4\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28345_ clknet_leaf_209_clock _01358_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_25557_ net667 _09039_ _09041_ _09033_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__o211a_1
X_13571_ _09930_ _09932_ _09933_ _09935_ VGND VGND VPWR VPWR _09936_ sky130_fd_sc_hd__and4_1
X_22769_ _06143_ net1321 _07276_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15310_ decode.regfile.registers_5\[1\] _11291_ _11304_ _11305_ VGND VGND VPWR VPWR
+ _11306_ sky130_fd_sc_hd__a22oi_2
X_24508_ _08068_ net1838 _08428_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28276_ clknet_leaf_60_clock _01298_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_16290_ decode.regfile.registers_20\[25\] _11101_ _11221_ _12261_ VGND VGND VPWR
+ VPWR _12262_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25488_ _08939_ _08992_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15241_ _10979_ _10958_ _11054_ _11062_ VGND VGND VPWR VPWR _11238_ sky130_fd_sc_hd__or4_2
XFILLER_0_35_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27227_ clknet_leaf_3_clock _00256_ VGND VGND VPWR VPWR decode.regfile.registers_29\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_24439_ _08398_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27158_ clknet_leaf_355_clock _00187_ VGND VGND VPWR VPWR decode.regfile.registers_27\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_15172_ _11168_ VGND VGND VPWR VPWR _11169_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_969 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26109_ decode.regfile.registers_10\[21\] _09356_ _09358_ _09359_ VGND VGND VPWR
+ VPWR _02596_ sky130_fd_sc_hd__o211a_1
X_14123_ _10147_ _10286_ VGND VGND VPWR VPWR _10329_ sky130_fd_sc_hd__nand2_1
X_19980_ _10798_ _05214_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27089_ clknet_leaf_352_clock _00118_ VGND VGND VPWR VPWR decode.regfile.registers_25\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18931_ _03984_ _03985_ _03986_ _03987_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__a31o_2
XFILLER_0_120_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14054_ _10290_ VGND VGND VPWR VPWR _10291_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18862_ _03751_ net306 _03757_ net238 _04156_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__a311o_2
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17813_ _11014_ _10936_ decode.regfile.registers_23\[25\] _12995_ VGND VGND VPWR
+ VPWR _03215_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_201_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18793_ _03796_ _04089_ _03706_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17744_ _13451_ net543 _13492_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__o21a_1
XFILLER_0_206_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14956_ _10983_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_193_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13907_ net2021 _10199_ _10204_ _10188_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17675_ decode.regfile.registers_2\[22\] _12835_ _12639_ decode.regfile.registers_3\[22\]
+ _12838_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_202_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14887_ _10923_ VGND VGND VPWR VPWR _10924_ sky130_fd_sc_hd__clkbuf_4
X_19414_ _04699_ _04702_ _03587_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_134_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16626_ _12590_ VGND VGND VPWR VPWR _12591_ sky130_fd_sc_hd__clkbuf_4
X_13838_ net563 _10153_ _10163_ _10162_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19345_ _04618_ _04129_ _04446_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_186_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16557_ _10597_ decode.immGen._imm_T_24\[17\] VGND VGND VPWR VPWR _12522_ sky130_fd_sc_hd__nor2b_4
X_13769_ _10060_ memory.io_wb_aluresult\[25\] _10004_ memory.io_wb_readdata\[25\]
+ VGND VGND VPWR VPWR _10109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15508_ decode.regfile.registers_2\[5\] _11369_ _11297_ _11121_ _11499_ VGND VGND
+ VPWR VPWR _11500_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_72_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19276_ _04365_ _04353_ _04272_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16488_ decode.regfile.registers_14\[31\] _11207_ _11273_ decode.regfile.registers_15\[31\]
+ _11361_ VGND VGND VPWR VPWR _12454_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18227_ csr.mcycle\[18\] _03556_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_61_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15439_ _10992_ _11066_ _11261_ _11432_ VGND VGND VPWR VPWR _11433_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18158_ _03507_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold303 io_fetch_data[8] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17109_ decode.regfile.registers_10\[8\] _10617_ _10594_ _10611_ _12690_ VGND VGND
+ VPWR VPWR _13066_ sky130_fd_sc_hd__o2111a_1
Xhold314 decode.regfile.registers_29\[7\] VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold325 _09983_ VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18089_ _03470_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold336 decode.regfile.registers_23\[7\] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_229_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold347 decode.regfile.registers_1\[20\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20120_ _05319_ _05325_ _05320_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__o21ai_1
Xhold358 decode.regfile.registers_13\[7\] VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_76_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_76_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold369 _10711_ VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_225_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20051_ _05269_ _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_182_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1003 fetch.bht.bhtTable_target_pc\[2\]\[23\] VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1014 fetch.bht.bhtTable_target_pc\[11\]\[27\] VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1025 fetch.bht.bhtTable_tag\[1\]\[24\] VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1036 decode.regfile.registers_5\[8\] VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 fetch.bht.bhtTable_tag\[12\]\[22\] VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__dlygate4sd3_1
X_23810_ _08060_ net1857 _08058_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__mux2_1
Xhold1058 fetch.bht.bhtTable_target_pc\[14\]\[22\] VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__dlygate4sd3_1
X_24790_ _08581_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_159_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1069 fetch.bht.bhtTable_target_pc\[1\]\[15\] VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23741_ _06103_ net1786 _09907_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__mux2_1
X_20953_ net2687 _05915_ _05911_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26460_ _09441_ _09533_ VGND VGND VPWR VPWR _09574_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_14_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_14_clock
+ sky130_fd_sc_hd__clkbuf_8
X_23672_ net2251 _10759_ _07983_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20884_ _05920_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_81_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25411_ _08905_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__clkbuf_4
X_22623_ net2795 _07190_ net2481 VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26391_ _09533_ VGND VGND VPWR VPWR _09535_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28130_ clknet_leaf_223_clock _01152_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22554_ _07143_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_118_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25342_ decode.io_wb_rd\[4\] decode.io_wb_regwrite VGND VGND VPWR VPWR _08902_ sky130_fd_sc_hd__and2b_4
XFILLER_0_146_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21505_ _06134_ net2245 _06263_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_29_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_29_clock
+ sky130_fd_sc_hd__clkbuf_8
X_28061_ clknet_leaf_198_clock _01083_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22485_ _06629_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__clkbuf_8
X_25273_ _08866_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27012_ clknet_leaf_342_clock _00041_ VGND VGND VPWR VPWR decode.regfile.registers_22\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24224_ _08286_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__clkbuf_1
X_21436_ _06233_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24155_ _08049_ net1378 _06274_ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21367_ _06115_ net2230 _06188_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23106_ _07122_ _07542_ _07544_ _07546_ _07127_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__o221a_1
X_20318_ _10864_ _10786_ _05482_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__and3_1
X_28963_ clknet_leaf_132_clock _01976_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_24086_ _08215_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold870 fetch.bht.bhtTable_target_pc\[4\]\[23\] VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__dlygate4sd3_1
X_21298_ net1053 _10821_ _06157_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold881 fetch.bht.bhtTable_tag\[1\]\[22\] VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__dlygate4sd3_1
X_23037_ _07480_ _07481_ _07082_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__mux2_1
Xhold892 fetch.bht.bhtTable_target_pc\[1\]\[26\] VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__dlygate4sd3_1
X_27914_ clknet_leaf_23_clock _00943_ VGND VGND VPWR VPWR csr.io_csr_write_address\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20249_ _10730_ _05433_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_229_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28894_ clknet_leaf_174_clock _01907_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_27845_ clknet_leaf_36_clock _00874_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2260 csr.mcycle\[17\] VGND VGND VPWR VPWR net2487 sky130_fd_sc_hd__dlygate4sd3_1
X_14810_ csr.io_mem_pc\[27\] _10769_ VGND VGND VPWR VPWR _10853_ sky130_fd_sc_hd__nor2_1
Xhold2271 decode.regfile.registers_8\[1\] VGND VGND VPWR VPWR net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2282 decode.regfile.registers_23\[5\] VGND VGND VPWR VPWR net2509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2293 decode.regfile.registers_25\[28\] VGND VGND VPWR VPWR net2520 sky130_fd_sc_hd__dlygate4sd3_1
X_27776_ clknet_leaf_327_clock _00805_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15790_ decode.regfile.registers_9\[12\] _11547_ _11773_ _11774_ _11184_ VGND VGND
+ VPWR VPWR _11775_ sky130_fd_sc_hd__a221oi_2
X_24988_ net340 csr.mcycle\[0\] csr.mcycle\[1\] VGND VGND VPWR VPWR _08705_ sky130_fd_sc_hd__a21o_1
Xhold1570 fetch.bht.bhtTable_target_pc\[5\]\[2\] VGND VGND VPWR VPWR net1797 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_24_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29515_ clknet_leaf_267_clock _02528_ VGND VGND VPWR VPWR decode.regfile.registers_8\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1581 fetch.bht.bhtTable_target_pc\[0\]\[21\] VGND VGND VPWR VPWR net1808 sky130_fd_sc_hd__dlygate4sd3_1
X_14741_ _10771_ _10775_ _10782_ decode.id_ex_pc_reg\[28\] VGND VGND VPWR VPWR _10784_
+ sky130_fd_sc_hd__a211oi_1
X_26727_ net1463 _09723_ _09728_ _09717_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__o211a_1
Xhold1592 fetch.bht.bhtTable_target_pc\[7\]\[24\] VGND VGND VPWR VPWR net1819 sky130_fd_sc_hd__dlygate4sd3_1
X_23939_ net862 _08097_ _08130_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17460_ _13087_ decode.regfile.registers_26\[16\] _13254_ _13047_ _13088_ VGND VGND
+ VPWR VPWR _13409_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_47_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29446_ clknet_leaf_262_clock _02459_ VGND VGND VPWR VPWR decode.regfile.registers_6\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14672_ decode.id_ex_pc_reg\[0\] _10703_ _10708_ _10712_ _10714_ VGND VGND VPWR VPWR
+ _10715_ sky130_fd_sc_hd__o2111ai_2
X_26658_ net1250 _09679_ _09687_ _09688_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16411_ _11396_ _12377_ _12378_ _12379_ VGND VGND VPWR VPWR _12380_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_103_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ _09983_ VGND VGND VPWR VPWR _09984_ sky130_fd_sc_hd__buf_4
XFILLER_0_67_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25609_ net803 _09068_ _09071_ _09059_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__o211a_1
X_17391_ decode.regfile.registers_9\[15\] _12776_ _12604_ _12532_ _12599_ VGND VGND
+ VPWR VPWR _13341_ sky130_fd_sc_hd__a41o_1
XFILLER_0_89_1209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29377_ clknet_leaf_256_clock _02390_ VGND VGND VPWR VPWR decode.regfile.registers_4\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26589_ _09621_ VGND VGND VPWR VPWR _09649_ sky130_fd_sc_hd__buf_2
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19130_ _03983_ _04234_ _04277_ _04318_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__o32a_1
XFILLER_0_67_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28328_ clknet_leaf_189_clock _01341_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_16342_ _11263_ decode.regfile.registers_22\[27\] _11404_ _11264_ _11265_ VGND VGND
+ VPWR VPWR _12312_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_137_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13554_ _09918_ _09919_ _09920_ VGND VGND VPWR VPWR _09921_ sky130_fd_sc_hd__nand3_4
XFILLER_0_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19061_ _04299_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28259_ clknet_leaf_92_clock _01281_ VGND VGND VPWR VPWR csr._minstret_T_3\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_16273_ _11156_ _12243_ _12244_ VGND VGND VPWR VPWR _12245_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18012_ _03374_ _03407_ _12704_ _03408_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__o211a_1
X_15224_ _10988_ _11118_ _11093_ VGND VGND VPWR VPWR _11221_ sky130_fd_sc_hd__and3_2
XFILLER_0_120_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15155_ _11151_ VGND VGND VPWR VPWR _11152_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14106_ _10102_ _10312_ VGND VGND VPWR VPWR _10320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_974 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19963_ _10707_ _03599_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__nor2_1
X_15086_ _11082_ VGND VGND VPWR VPWR _11083_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14037_ net2215 _10271_ _10279_ _10275_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__o211a_1
X_18914_ _04196_ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__nand2_1
X_19894_ _03781_ _03788_ _03865_ _05162_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_207_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18845_ _04142_ _04143_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__nor2_4
XFILLER_0_101_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_220_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_220_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_220_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18776_ _04074_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15988_ _11124_ decode.regfile.registers_16\[17\] _11127_ _11967_ VGND VGND VPWR
+ VPWR _11968_ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17727_ decode.regfile.registers_14\[23\] _12984_ _03115_ _03130_ _12874_ VGND VGND
+ VPWR VPWR _03131_ sky130_fd_sc_hd__o221a_1
XFILLER_0_171_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14939_ _10579_ decode.control.io_opcode\[3\] decode.control.io_opcode\[4\] _10584_
+ VGND VGND VPWR VPWR _10968_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_37_1322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17658_ _13339_ _03061_ _03062_ _03063_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16609_ _10594_ _10598_ _10588_ _12540_ VGND VGND VPWR VPWR _12574_ sky130_fd_sc_hd__or4_1
XFILLER_0_159_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17589_ _13451_ decode.regfile.registers_30\[20\] _13492_ VGND VGND VPWR VPWR _02996_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19328_ _04424_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__buf_4
XFILLER_0_156_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19259_ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_171_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22270_ fetch.bht.bhtTable_tag\[12\]\[6\] fetch.bht.bhtTable_tag\[13\]\[6\] _06617_
+ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21221_ _06106_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_184_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_184_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21152_ _06069_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold155 io_fetch_data[10] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold166 fetch.bht.bhtTable_valid\[14\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold177 fetch.btb.btbTable\[6\]\[0\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold188 fetch.btb.btbTable\[5\]\[0\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
X_20103_ decode.id_ex_imm_reg\[15\] _10681_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__or2_1
XFILLER_0_217_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold199 _10725_ VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
X_25960_ net2284 _09270_ _09273_ _09264_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__o211a_1
X_21083_ _06028_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20034_ _05248_ _05252_ _05249_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__o21ai_1
X_24911_ csr._mcycle_T_3\[38\] _08654_ _07179_ VGND VGND VPWR VPWR _08655_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_60_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25891_ _08964_ _09223_ VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__nand2_1
X_27630_ clknet_leaf_44_clock _00659_ VGND VGND VPWR VPWR execute.io_reg_pc\[7\] sky130_fd_sc_hd__dfxtp_1
X_24842_ _06119_ net1627 _08607_ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_12 _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_23 _03314_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27561_ clknet_leaf_157_clock _00590_ VGND VGND VPWR VPWR csr.io_mem_pc\[2\] sky130_fd_sc_hd__dfxtp_2
XINSDIODE1_34 _08929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24773_ _08572_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_45 _09949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ net1609 _06588_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__or2_1
XINSDIODE1_56 _10073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_205_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29300_ clknet_leaf_232_clock _02313_ VGND VGND VPWR VPWR decode.regfile.registers_1\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_67 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26512_ net1529 _09592_ _09604_ _09595_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23724_ net1557 _10773_ _08003_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__mux2_1
XINSDIODE1_78 _10240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_89 _10595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20936_ _05857_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__buf_2
X_27492_ clknet_leaf_34_clock _00521_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29231_ clknet_leaf_124_clock _02244_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_26443_ net2406 _09561_ _09564_ _09553_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__o211a_1
X_23655_ net1163 _10800_ _07972_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__mux2_1
X_20867_ _03582_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_42_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29162_ clknet_leaf_205_clock _02175_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_22606_ csr._minstret_T_3\[49\] csr._minstret_T_3\[48\] csr._minstret_T_3\[47\] _07174_
+ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26374_ _09417_ VGND VGND VPWR VPWR _09525_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_42_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23586_ _06117_ net1741 _07930_ VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20798_ _05873_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__clkbuf_1
X_28113_ clknet_leaf_81_clock net2649 VGND VGND VPWR VPWR csr.minstret\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25325_ _08893_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22537_ execute.io_target_pc\[1\] _07091_ _06041_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29093_ clknet_leaf_70_clock _02106_ VGND VGND VPWR VPWR csr._mcycle_T_3\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28044_ clknet_leaf_216_clock _01066_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25256_ _08095_ net1351 _08848_ VGND VGND VPWR VPWR _08858_ sky130_fd_sc_hd__mux2_1
X_22468_ _06720_ _06769_ _06822_ _07062_ _03591_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__o41a_4
XFILLER_0_106_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24207_ _08101_ net1788 _06251_ VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__mux2_1
X_21419_ _06224_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__clkbuf_1
X_22399_ _06650_ _06993_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__and2b_1
X_25187_ net415 _08822_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24138_ _08242_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16960_ _12496_ _12918_ _12919_ _12920_ VGND VGND VPWR VPWR _12921_ sky130_fd_sc_hd__a31o_1
X_24069_ net1503 execute.io_target_pc\[22\] _08198_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__mux2_1
X_28946_ clknet_leaf_106_clock _01959_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15911_ _11070_ _11470_ decode.regfile.registers_10\[15\] _11381_ VGND VGND VPWR
+ VPWR _11893_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_120_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28877_ clknet_leaf_101_clock _01890_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16891_ decode.regfile.registers_14\[3\] _12669_ _12828_ _12851_ _12852_ VGND VGND
+ VPWR VPWR _12853_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_188_Right_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18630_ _03925_ _03700_ _03688_ decode.id_ex_rs1_data_reg\[16\] _03928_ VGND VGND
+ VPWR VPWR _03929_ sky130_fd_sc_hd__o221a_4
XFILLER_0_216_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15842_ decode.regfile.registers_25\[13\] _11333_ _11336_ decode.regfile.registers_24\[13\]
+ VGND VGND VPWR VPWR _11826_ sky130_fd_sc_hd__o22a_1
X_27828_ clknet_leaf_317_clock _00857_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2090 execute.csr_write_data_out_reg\[18\] VGND VGND VPWR VPWR net2317 sky130_fd_sc_hd__dlygate4sd3_1
X_18561_ decode.id_ex_rs2_data_reg\[30\] _03747_ _03764_ _03857_ VGND VGND VPWR VPWR
+ _03860_ sky130_fd_sc_hd__o22a_1
X_15773_ _11646_ _11253_ _11064_ decode.regfile.registers_29\[11\] _11758_ VGND VGND
+ VPWR VPWR _11759_ sky130_fd_sc_hd__o221a_1
X_27759_ clknet_leaf_316_clock _00788_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_17512_ _13456_ _13457_ _13458_ VGND VGND VPWR VPWR _13459_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14724_ _10766_ VGND VGND VPWR VPWR _10767_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_185_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18492_ _03789_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17443_ _11018_ _12977_ _12637_ decode.regfile.registers_11\[16\] VGND VGND VPWR
+ VPWR _13392_ sky130_fd_sc_hd__or4b_1
XFILLER_0_68_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29429_ clknet_leaf_260_clock _02442_ VGND VGND VPWR VPWR decode.regfile.registers_5\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14655_ execute.io_target_pc\[29\] VGND VGND VPWR VPWR _10698_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13606_ memory.csr_read_data_out_reg\[2\] _09942_ _09967_ _09968_ VGND VGND VPWR
+ VPWR _09969_ sky130_fd_sc_hd__a2bb2o_4
X_17374_ decode.regfile.registers_15\[14\] _12650_ _12723_ _12574_ VGND VGND VPWR
+ VPWR _13325_ sky130_fd_sc_hd__o31a_1
XFILLER_0_83_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14586_ _10628_ VGND VGND VPWR VPWR _10629_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_188_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_188_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19113_ _03863_ _04255_ _04338_ _04286_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__o211a_2
X_16325_ decode.regfile.registers_18\[26\] _11455_ _11456_ _12295_ VGND VGND VPWR
+ VPWR _12296_ sky130_fd_sc_hd__a211o_1
X_13537_ net576 _09912_ VGND VGND VPWR VPWR _09913_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19044_ _04281_ _04283_ _04342_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__o21ai_1
X_16256_ decode.regfile.registers_23\[24\] _11262_ _12204_ _12228_ _11335_ VGND VGND
+ VPWR VPWR _12229_ sky130_fd_sc_hd__o221a_1
XFILLER_0_152_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15207_ _11167_ VGND VGND VPWR VPWR _11204_ sky130_fd_sc_hd__clkbuf_4
X_16187_ decode.regfile.registers_21\[22\] _11061_ _11099_ _11229_ _12161_ VGND VGND
+ VPWR VPWR _12162_ sky130_fd_sc_hd__o311a_1
XFILLER_0_11_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15138_ _10645_ _10623_ _11082_ VGND VGND VPWR VPWR _11135_ sky130_fd_sc_hd__or3_2
XFILLER_0_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_1202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19946_ _05207_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__clkbuf_1
X_15069_ _11065_ VGND VGND VPWR VPWR _11066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19877_ _04525_ _05146_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18828_ _03797_ _04124_ _03890_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_207_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18759_ execute.csr_read_data_out_reg\[7\] _03661_ _03660_ VGND VGND VPWR VPWR _04058_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_223_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21770_ net1445 _10772_ _06439_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20721_ _05809_ decode.id_ex_rs1_data_reg\[19\] VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20652_ _05540_ csr.io_mret_vector\[30\] _05565_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__o21a_1
X_23440_ decode.immGen._imm_T_10\[2\] _07847_ _05206_ VGND VGND VPWR VPWR _07855_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23371_ _07793_ _07794_ _07795_ _07072_ _07371_ VGND VGND VPWR VPWR _07796_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_144_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20583_ _05439_ _05723_ _03449_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__and3b_1
XFILLER_0_74_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25110_ _08783_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22322_ _06707_ fetch.bht.bhtTable_tag\[11\]\[8\] _06649_ VGND VGND VPWR VPWR _06917_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26090_ net2166 _09343_ _09348_ _09346_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_76_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22253_ _06631_ _06843_ _06845_ _06847_ _06640_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__o221ai_4
X_25041_ net2658 _08704_ _08740_ csr.mcycle\[18\] VGND VGND VPWR VPWR _08741_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_132_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21204_ _06097_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__clkbuf_1
X_22184_ fetch.bht.bhtTable_tag\[12\]\[25\] fetch.bht.bhtTable_tag\[13\]\[25\] _06646_
+ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28800_ clknet_leaf_171_clock _01813_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_21135_ _06060_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__clkbuf_1
X_29780_ clknet_leaf_295_clock _02793_ VGND VGND VPWR VPWR decode.regfile.registers_16\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26992_ clknet_leaf_333_clock _00021_ VGND VGND VPWR VPWR decode.regfile.registers_22\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28731_ clknet_leaf_172_clock _01744_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_25943_ _09263_ VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__clkbuf_4
X_21066_ _06019_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20017_ decode.id_ex_imm_reg\[3\] decode.id_ex_pc_reg\[3\] VGND VGND VPWR VPWR _05241_
+ sky130_fd_sc_hd__nand2_1
X_28662_ clknet_leaf_124_clock _01675_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25874_ _08945_ _09223_ VGND VGND VPWR VPWR _09224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27613_ clknet_leaf_152_clock _00642_ VGND VGND VPWR VPWR execute.io_target_pc\[22\]
+ sky130_fd_sc_hd__dfxtp_4
X_24825_ _06103_ net1215 _08422_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__mux2_1
X_28593_ clknet_leaf_103_clock _01606_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_1264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27544_ clknet_leaf_44_clock _00573_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_96_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24756_ _08049_ net1458 _08563_ VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21968_ net884 _06574_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _08004_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_139_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27475_ clknet_leaf_52_clock _00504_ VGND VGND VPWR VPWR csr.io_csr_address\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_20919_ _05937_ _05933_ net44 VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24687_ _08049_ net1728 _06306_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21899_ _06039_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__clkbuf_4
X_29214_ clknet_leaf_97_clock _02227_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26426_ _09406_ _09545_ VGND VGND VPWR VPWR _09555_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_29_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _09984_ _10507_ VGND VGND VPWR VPWR _10513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23638_ net1472 _10812_ _07961_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29145_ clknet_leaf_92_clock _02158_ VGND VGND VPWR VPWR csr.mcycle\[29\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_61_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26357_ _09490_ VGND VGND VPWR VPWR _09515_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_61_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ _10008_ _10464_ VGND VGND VPWR VPWR _10473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23569_ _09900_ _06281_ _09894_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__or3b_4
XFILLER_0_153_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16110_ _12055_ _12085_ _12086_ VGND VGND VPWR VPWR _12087_ sky130_fd_sc_hd__o21ai_2
X_25308_ _08884_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__clkbuf_1
X_29076_ clknet_leaf_198_clock _02089_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17090_ _10928_ decode.regfile.registers_26\[7\] _12814_ _13047_ _11027_ VGND VGND
+ VPWR VPWR _13048_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26288_ _09420_ _09472_ VGND VGND VPWR VPWR _09476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28027_ clknet_leaf_204_clock _01049_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16041_ decode.regfile.registers_9\[19\] _11280_ _11134_ _11509_ VGND VGND VPWR VPWR
+ _12019_ sky130_fd_sc_hd__a31o_1
X_25239_ _08849_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19800_ _04304_ _05072_ _04537_ _04898_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__a2bb2o_1
X_17992_ _12602_ decode.regfile.registers_9\[30\] _12652_ _03388_ VGND VGND VPWR VPWR
+ _03389_ sky130_fd_sc_hd__o211a_1
X_19731_ _05006_ _04964_ _04352_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16943_ decode.regfile.registers_17\[4\] _12719_ _12826_ VGND VGND VPWR VPWR _12904_
+ sky130_fd_sc_hd__o21a_1
X_28929_ clknet_leaf_175_clock _01942_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16874_ _12638_ VGND VGND VPWR VPWR _12836_ sky130_fd_sc_hd__clkbuf_4
X_19662_ _03959_ _03639_ _04667_ _04192_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15825_ _11803_ _11807_ _11808_ VGND VGND VPWR VPWR _11809_ sky130_fd_sc_hd__o21a_1
X_18613_ _03708_ decode.id_ex_imm_reg\[17\] _03906_ _03907_ _03911_ VGND VGND VPWR
+ VPWR _03912_ sky130_fd_sc_hd__a221o_2
X_19593_ _03934_ _04253_ _04380_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15756_ _11728_ _11740_ _11741_ VGND VGND VPWR VPWR _11742_ sky130_fd_sc_hd__o21a_1
X_18544_ decode.id_ex_rs1_data_reg\[24\] _03688_ _03842_ _03701_ VGND VGND VPWR VPWR
+ _03843_ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14707_ _10748_ execute.io_target_pc\[3\] _10677_ execute.io_target_pc\[22\] VGND
+ VGND VPWR VPWR _10750_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18475_ net353 VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__buf_4
X_15687_ _11050_ decode.regfile.registers_25\[9\] _11090_ VGND VGND VPWR VPWR _11675_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_213_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_215_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17426_ _13099_ _13262_ _13182_ decode.regfile.registers_29\[15\] _13375_ VGND VGND
+ VPWR VPWR _13376_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_215_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14638_ decode.id_ex_pc_reg\[15\] VGND VGND VPWR VPWR _10681_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17357_ decode.regfile.registers_13\[14\] _12533_ _12587_ _12662_ VGND VGND VPWR
+ VPWR _13308_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14569_ _10611_ VGND VGND VPWR VPWR _10612_ sky130_fd_sc_hd__buf_4
XFILLER_0_172_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16308_ decode.regfile.registers_1\[26\] _11116_ _11056_ _11108_ VGND VGND VPWR VPWR
+ _12279_ sky130_fd_sc_hd__and4_1
X_17288_ _12585_ _13223_ _13239_ _13240_ VGND VGND VPWR VPWR _13241_ sky130_fd_sc_hd__o31a_1
XFILLER_0_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19027_ _04045_ _04054_ _04307_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__mux2_1
X_16239_ decode.regfile.registers_4\[24\] _11410_ _12208_ _12211_ VGND VGND VPWR VPWR
+ _12212_ sky130_fd_sc_hd__a2bb2oi_1
XPHY_EDGE_ROW_224_Right_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19929_ _05192_ _05194_ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22940_ _07385_ _07387_ _07388_ _07389_ _07080_ _06637_ VGND VGND VPWR VPWR _07390_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_177_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22871_ net747 _10787_ _07324_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24610_ _08487_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_175_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21822_ _06480_ csr._csr_read_data_T_9\[0\] _06484_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__a21o_1
XFILLER_0_195_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25590_ _08964_ _09049_ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24541_ _08101_ net1567 _09902_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21753_ _06427_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27260_ clknet_leaf_12_clock _00289_ VGND VGND VPWR VPWR decode.regfile.registers_30\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_20704_ _05809_ decode.id_ex_rs1_data_reg\[12\] _05798_ VGND VGND VPWR VPWR _05820_
+ sky130_fd_sc_hd__a21oi_1
X_24472_ _08099_ net2009 _08411_ VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21684_ csr.minstret\[21\] csr.minstret\[22\] csr.minstret\[23\] _06383_ VGND VGND
+ VPWR VPWR _06389_ sky130_fd_sc_hd__and4_1
XFILLER_0_175_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26211_ net2618 _09419_ _09427_ _09418_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__o211a_1
X_23423_ _05857_ _07345_ _10672_ _07844_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20635_ _05627_ csr.io_mret_vector\[27\] _05603_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__o21a_1
X_27191_ clknet_leaf_355_clock _00220_ VGND VGND VPWR VPWR decode.regfile.registers_28\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26142_ net210 VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__buf_4
X_23354_ _07776_ _07777_ _07778_ _07779_ _07371_ _07084_ VGND VGND VPWR VPWR _07780_
+ sky130_fd_sc_hd__mux4_2
X_20566_ csr.mcycle\[17\] _05588_ _05618_ csr._csr_read_data_T_8\[17\] _05708_ VGND
+ VGND VPWR VPWR _05709_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22305_ _06690_ _06899_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26073_ net2439 _09329_ _09338_ _09333_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23285_ net80 net79 _07651_ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__and3_1
X_20497_ csr.io_mret_vector\[8\] _05580_ _05581_ csr.mscratch\[8\] _05648_ VGND VGND
+ VPWR VPWR _05649_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25024_ csr.mcycle\[12\] csr.mcycle\[11\] _08725_ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__and3_1
X_29901_ clknet_leaf_301_clock _02914_ VGND VGND VPWR VPWR decode.regfile.registers_20\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22236_ fetch.bht.bhtTable_tag\[8\]\[15\] fetch.bht.bhtTable_tag\[9\]\[15\] fetch.bht.bhtTable_tag\[10\]\[15\]
+ fetch.bht.bhtTable_tag\[11\]\[15\] _06754_ _06675_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__mux4_1
XFILLER_0_225_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22167_ _06690_ _06761_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__and2b_1
X_29832_ clknet_5_16__leaf_clock _02845_ VGND VGND VPWR VPWR decode.regfile.registers_18\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21118_ _06051_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22098_ _06690_ _06692_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__and2b_1
X_26975_ net197 _09862_ VGND VGND VPWR VPWR _09871_ sky130_fd_sc_hd__nand2_1
X_29763_ clknet_leaf_291_clock _02776_ VGND VGND VPWR VPWR decode.regfile.registers_16\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28714_ clknet_leaf_98_clock _01727_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13940_ _10198_ VGND VGND VPWR VPWR _10223_ sky130_fd_sc_hd__buf_2
X_25926_ _08922_ _09253_ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__nand2_1
X_21049_ _09954_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__buf_2
XFILLER_0_227_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29694_ clknet_leaf_311_clock _02707_ VGND VGND VPWR VPWR decode.regfile.registers_14\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28645_ clknet_leaf_137_clock _01658_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13871_ net783 _10180_ _10182_ _10175_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__o211a_1
X_25857_ net681 _09213_ _09214_ _09209_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15610_ decode.regfile.registers_21\[7\] _11267_ _11099_ _11228_ _11599_ VGND VGND
+ VPWR VPWR _11600_ sky130_fd_sc_hd__o311a_1
XFILLER_0_198_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24808_ _08101_ net1633 _08585_ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28576_ clknet_leaf_169_clock _01589_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_16590_ _10611_ VGND VGND VPWR VPWR _12555_ sky130_fd_sc_hd__clkbuf_4
X_25788_ net523 _09170_ _09174_ _09169_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_1094 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_107 _10935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27527_ clknet_leaf_46_clock _00556_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dfxtp_2
X_15541_ decode.regfile.registers_13\[6\] _11275_ _11278_ decode.regfile.registers_12\[6\]
+ VGND VGND VPWR VPWR _11532_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24739_ _08101_ net1562 _06283_ VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_118 _11054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_129 _11217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18260_ _10756_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27458_ clknet_leaf_137_clock _00487_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[24\]
+ sky130_fd_sc_hd__dfxtp_4
X_15472_ _11308_ VGND VGND VPWR VPWR _11465_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_167_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17211_ _13139_ _13163_ _13164_ _13165_ VGND VGND VPWR VPWR _13166_ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26409_ _09533_ VGND VGND VPWR VPWR _09545_ sky130_fd_sc_hd__clkbuf_4
X_14423_ _10142_ _10462_ VGND VGND VPWR VPWR _10502_ sky130_fd_sc_hd__nand2_1
X_18191_ decode.control.io_funct7\[2\] decode.control.io_funct7\[1\] decode.control.io_funct7\[0\]
+ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27389_ clknet_leaf_9_clock _00418_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29128_ clknet_leaf_76_clock net2644 VGND VGND VPWR VPWR csr.mcycle\[12\] sky130_fd_sc_hd__dfxtp_2
X_17142_ _13055_ net458 _13097_ VGND VGND VPWR VPWR _13098_ sky130_fd_sc_hd__o21a_1
X_14354_ _10462_ VGND VGND VPWR VPWR _10463_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29059_ clknet_leaf_217_clock _02072_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_17073_ _12672_ VGND VGND VPWR VPWR _13031_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14285_ net617 _10419_ _10423_ _10411_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16024_ decode.regfile.registers_17\[18\] _10652_ _11112_ _11118_ _12002_ VGND VGND
+ VPWR VPWR _12003_ sky130_fd_sc_hd__a41o_1
XFILLER_0_122_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17975_ _02997_ _12767_ _12965_ decode.regfile.registers_29\[29\] _03372_ VGND VGND
+ VPWR VPWR _03373_ sky130_fd_sc_hd__o221a_1
XFILLER_0_224_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19714_ _04981_ _04989_ _04883_ _04990_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__o22a_2
X_16926_ decode.regfile.registers_6\[4\] _12880_ _12881_ _12886_ VGND VGND VPWR VPWR
+ _12887_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_204_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19645_ _04537_ _04270_ _04924_ _04463_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__or4_1
X_16857_ _12765_ _12768_ _12493_ decode.regfile.registers_29\[2\] _12819_ VGND VGND
+ VPWR VPWR _12820_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_217_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_196_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15808_ _11251_ _11259_ decode.regfile.registers_27\[12\] _11763_ _11792_ VGND VGND
+ VPWR VPWR _11793_ sky130_fd_sc_hd__o32a_1
XFILLER_0_88_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_217_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16788_ _11022_ _12567_ _12586_ _12751_ VGND VGND VPWR VPWR _12752_ sky130_fd_sc_hd__a31o_1
X_19576_ _04198_ _04359_ _04504_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15739_ _11571_ decode.regfile.registers_30\[11\] _11722_ _11723_ _11724_ VGND VGND
+ VPWR VPWR _11725_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18527_ net188 _03825_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18458_ _03753_ _03754_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_173_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17409_ _12719_ _13358_ VGND VGND VPWR VPWR _13359_ sky130_fd_sc_hd__nand2_1
X_18389_ _03687_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20420_ csr._minstret_T_3\[33\] _05577_ _05578_ _05563_ csr._csr_read_data_T_9\[1\]
+ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20351_ _10733_ _05514_ _05416_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_168_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23070_ fetch.bht.bhtTable_target_pc\[10\]\[10\] fetch.bht.bhtTable_target_pc\[11\]\[10\]
+ _07069_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__mux2_1
X_20282_ _05461_ _05462_ _05420_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22021_ net301 VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1900 decode.regfile.registers_8\[14\] VGND VGND VPWR VPWR net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1911 decode.io_id_pc\[24\] VGND VGND VPWR VPWR net2138 sky130_fd_sc_hd__dlygate4sd3_1
X_26760_ _09438_ _09708_ VGND VGND VPWR VPWR _09747_ sky130_fd_sc_hd__nand2_1
X_23972_ net1423 execute.io_target_pc\[7\] _08153_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__mux2_1
Xhold1922 decode.regfile.registers_23\[18\] VGND VGND VPWR VPWR net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1933 decode.regfile.registers_26\[18\] VGND VGND VPWR VPWR net2160 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1944 decode.io_id_pc\[22\] VGND VGND VPWR VPWR net2171 sky130_fd_sc_hd__dlygate4sd3_1
X_25711_ net820 _09125_ _09130_ _09129_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__o211a_1
X_22923_ _07103_ _07373_ VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__and2b_1
Xhold1955 fetch.bht.bhtTable_tag\[7\]\[20\] VGND VGND VPWR VPWR net2182 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1966 fetch.bht.bhtTable_tag\[5\]\[3\] VGND VGND VPWR VPWR net2193 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26691_ _09932_ _10149_ _03672_ VGND VGND VPWR VPWR _09707_ sky130_fd_sc_hd__and3_1
XFILLER_0_224_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1977 fetch.bht.bhtTable_tag\[15\]\[21\] VGND VGND VPWR VPWR net2204 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1988 decode.regfile.registers_25\[26\] VGND VGND VPWR VPWR net2215 sky130_fd_sc_hd__dlygate4sd3_1
X_28430_ clknet_leaf_246_clock _01443_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[11\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_79_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1999 fetch.bht.bhtTable_target_pc\[9\]\[18\] VGND VGND VPWR VPWR net2226 sky130_fd_sc_hd__dlygate4sd3_1
X_25642_ _08941_ _09079_ VGND VGND VPWR VPWR _09090_ sky130_fd_sc_hd__nand2_1
X_22854_ net1615 _10872_ _09898_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28361_ clknet_leaf_219_clock _01374_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_21805_ csr._mcycle_T_2\[3\] _06457_ _06466_ _06472_ VGND VGND VPWR VPWR _06473_
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_196_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25573_ net2589 _09039_ _09050_ _09046_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22785_ _07287_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27312_ clknet_leaf_238_clock _00341_ VGND VGND VPWR VPWR fetch.btb.btbTable\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_24524_ _08443_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28292_ clknet_leaf_85_clock _01314_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_21736_ _06430_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27243_ clknet_leaf_0_clock _00272_ VGND VGND VPWR VPWR decode.regfile.registers_29\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24455_ _08083_ net1414 _08400_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21667_ net567 _06375_ _06376_ _06352_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_35_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23406_ _05857_ _07345_ _10672_ _07828_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20618_ _05750_ _05753_ _05630_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__o21a_2
XFILLER_0_149_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27174_ clknet_leaf_362_clock _00203_ VGND VGND VPWR VPWR decode.regfile.registers_27\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_24386_ _08370_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21598_ net512 _06325_ _06323_ csr.minstret\[0\] csr.minstret\[1\] VGND VGND VPWR
+ VPWR _06326_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_10_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26125_ net701 _09356_ _09367_ _09359_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__o211a_1
X_23337_ _07762_ _07763_ _07075_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20549_ csr._minstret_T_3\[47\] _05555_ _05581_ csr.mscratch\[15\] _05559_ VGND VGND
+ VPWR VPWR _05694_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_312_clock clknet_5_18__leaf_clock VGND VGND VPWR VPWR clknet_leaf_312_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14070_ _10286_ VGND VGND VPWR VPWR _10299_ sky130_fd_sc_hd__clkbuf_4
X_26056_ _09327_ VGND VGND VPWR VPWR _09328_ sky130_fd_sc_hd__buf_4
X_23268_ _07698_ _07699_ _07081_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25007_ net777 _08701_ net1256 _05856_ _08718_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_56_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22219_ fetch.bht.bhtTable_tag\[8\]\[20\] fetch.bht.bhtTable_tag\[9\]\[20\] _06616_
+ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23199_ csr._csr_read_data_T_8\[18\] _06038_ csr.io_mret_vector\[18\] _06463_ VGND
+ VGND VPWR VPWR _07634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_219_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29815_ clknet_leaf_296_clock _02828_ VGND VGND VPWR VPWR decode.regfile.registers_17\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_327_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_327_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_218_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14972_ _10996_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__clkbuf_1
X_29746_ clknet_leaf_285_clock _02759_ VGND VGND VPWR VPWR decode.regfile.registers_15\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_17760_ decode.regfile.registers_10\[24\] _12790_ _12792_ VGND VGND VPWR VPWR _03163_
+ sky130_fd_sc_hd__o21a_1
X_26958_ _10068_ _09849_ VGND VGND VPWR VPWR _09861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13923_ _10031_ _10210_ VGND VGND VPWR VPWR _10214_ sky130_fd_sc_hd__nand2_1
X_16711_ _12576_ decode.regfile.registers_16\[0\] _12580_ _12675_ VGND VGND VPWR VPWR
+ _12676_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17691_ decode.regfile.registers_19\[22\] _12678_ _03075_ _03095_ _12544_ VGND VGND
+ VPWR VPWR _03096_ sky130_fd_sc_hd__o221a_1
X_25909_ net1536 _09242_ _09244_ _09235_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_1002 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29677_ clknet_leaf_282_clock _02690_ VGND VGND VPWR VPWR decode.regfile.registers_13\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_26889_ net1997 _09809_ _09821_ _09812_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16642_ _12606_ VGND VGND VPWR VPWR _12607_ sky130_fd_sc_hd__buf_4
X_19430_ _04153_ _04154_ _04166_ _04164_ _04684_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__a221o_1
X_28628_ clknet_leaf_119_clock _01641_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_13854_ net506 _10167_ _10172_ _10162_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19361_ _04245_ _03705_ _04503_ _04345_ _04362_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__a311o_1
X_16573_ _12537_ VGND VGND VPWR VPWR _12538_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28559_ clknet_leaf_220_clock _01572_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13785_ _10122_ _10075_ VGND VGND VPWR VPWR _10123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15524_ _11127_ decode.regfile.registers_17\[5\] _11105_ _11515_ VGND VGND VPWR VPWR
+ _11516_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18312_ _03621_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19292_ _04050_ _04051_ _04516_ _04529_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_155_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18243_ _03575_ _03576_ _03577_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__nor3_1
X_15455_ _11347_ VGND VGND VPWR VPWR _11448_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14406_ _10097_ _10487_ VGND VGND VPWR VPWR _10493_ sky130_fd_sc_hd__nand2_1
X_18174_ _03463_ _03464_ _03465_ decode.control.io_funct7\[6\] VGND VGND VPWR VPWR
+ _03515_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_108_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15386_ _10655_ _10636_ _11314_ _10660_ VGND VGND VPWR VPWR _11381_ sky130_fd_sc_hd__or4b_4
XFILLER_0_26_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17125_ _13081_ _10937_ decode.regfile.registers_23\[8\] _13041_ VGND VGND VPWR VPWR
+ _13082_ sky130_fd_sc_hd__or4_1
XFILLER_0_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14337_ net935 _10447_ _10452_ _10453_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap204 _03784_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_4
Xhold507 csr.io_ecause\[2\] VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap215 _12635_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold518 decode.regfile.registers_15\[15\] VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ _12530_ _12616_ _12557_ decode.regfile.registers_0\[7\] VGND VGND VPWR VPWR
+ _13014_ sky130_fd_sc_hd__a31o_1
Xhold529 decode.regfile.registers_26\[15\] VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14268_ _10128_ _10375_ VGND VGND VPWR VPWR _10413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16007_ decode.regfile.registers_14\[18\] _11207_ _11273_ decode.regfile.registers_15\[18\]
+ _11361_ VGND VGND VPWR VPWR _11986_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_206_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_206_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14199_ net456 _10333_ _10372_ _10369_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_198_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 decode.regfile.registers_2\[2\] VGND VGND VPWR VPWR net1434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1218 fetch.bht.bhtTable_tag\[4\]\[18\] VGND VGND VPWR VPWR net1445 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_198_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ decode.regfile.registers_13\[29\] _12775_ _03354_ _03355_ _12663_ VGND VGND
+ VPWR VPWR _03356_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1229 execute.csr_write_address_out_reg\[4\] VGND VGND VPWR VPWR net1456 sky130_fd_sc_hd__dlygate4sd3_1
X_16909_ _12765_ _12768_ _12493_ decode.regfile.registers_29\[3\] _12870_ VGND VGND
+ VPWR VPWR _12871_ sky130_fd_sc_hd__o221a_1
XFILLER_0_164_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17889_ _12822_ decode.regfile.registers_21\[27\] _13164_ _03288_ VGND VGND VPWR
+ VPWR _03289_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19628_ _04204_ _04206_ _03638_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19559_ _04211_ _04840_ _04841_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_220_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22570_ csr._minstret_T_3\[40\] _07153_ _07154_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21521_ _06278_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24240_ _08068_ net1725 _08289_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21452_ _06143_ net2012 _06241_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20403_ _05562_ _05522_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_116_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24171_ _08259_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__clkbuf_1
X_21383_ _06204_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_116_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23122_ fetch.bht.bhtTable_target_pc\[0\]\[13\] fetch.bht.bhtTable_target_pc\[1\]\[13\]
+ _07067_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20334_ _10790_ decode.id_ex_pc_reg\[26\] _10854_ _05494_ VGND VGND VPWR VPWR _05502_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27930_ clknet_leaf_161_clock _00009_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_23053_ _06718_ _07472_ VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__nand2_1
X_20265_ _05448_ _05449_ _05420_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_129_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_79_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22004_ csr.mscratch\[24\] _06601_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__or2_1
X_27861_ clknet_leaf_316_clock _00890_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_20196_ _05393_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__nor2_1
Xhold2420 decode.regfile.registers_12\[22\] VGND VGND VPWR VPWR net2647 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2431 csr._mcycle_T_2\[18\] VGND VGND VPWR VPWR net2658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29600_ clknet_leaf_271_clock _02613_ VGND VGND VPWR VPWR decode.regfile.registers_11\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_26812_ net1416 _09766_ _09777_ _09771_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__o211a_1
Xhold2442 fetch.btb.btbTable\[3\]\[1\] VGND VGND VPWR VPWR net2669 sky130_fd_sc_hd__dlygate4sd3_1
X_27792_ clknet_leaf_335_clock _00821_ VGND VGND VPWR VPWR memory.io_wb_readdata\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2453 decode.regfile.registers_0\[19\] VGND VGND VPWR VPWR net2680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2464 decode.id_ex_rs1_data_reg\[16\] VGND VGND VPWR VPWR net2691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1730 csr._mcycle_T_2\[27\] VGND VGND VPWR VPWR net1957 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2475 csr._csr_read_data_T_8\[6\] VGND VGND VPWR VPWR net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2486 decode.immGen._imm_T_10\[0\] VGND VGND VPWR VPWR net2713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1741 decode.regfile.registers_16\[16\] VGND VGND VPWR VPWR net1968 sky130_fd_sc_hd__dlygate4sd3_1
X_26743_ _09422_ _09733_ VGND VGND VPWR VPWR _09738_ sky130_fd_sc_hd__nand2_1
X_29531_ clknet_leaf_313_clock _02544_ VGND VGND VPWR VPWR decode.regfile.registers_9\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1752 fetch.bht.bhtTable_target_pc\[14\]\[6\] VGND VGND VPWR VPWR net1979 sky130_fd_sc_hd__dlygate4sd3_1
X_23955_ net839 _08113_ _06156_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2497 execute.io_reg_pc\[27\] VGND VGND VPWR VPWR net2724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1763 decode.regfile.registers_26\[10\] VGND VGND VPWR VPWR net1990 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1774 fetch.bht.bhtTable_tag\[13\]\[7\] VGND VGND VPWR VPWR net2001 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1785 fetch.bht.bhtTable_tag\[6\]\[20\] VGND VGND VPWR VPWR net2012 sky130_fd_sc_hd__dlygate4sd3_1
X_22906_ _06656_ _06795_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__nand2_1
X_29462_ clknet_leaf_261_clock _02475_ VGND VGND VPWR VPWR decode.regfile.registers_6\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26674_ net2465 _09692_ _09697_ _09688_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__o211a_1
Xhold1796 decode.regfile.registers_9\[29\] VGND VGND VPWR VPWR net2023 sky130_fd_sc_hd__dlygate4sd3_1
X_23886_ _08111_ net2141 _07940_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28413_ clknet_leaf_52_clock _01426_ VGND VGND VPWR VPWR decode.control.io_opcode\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_88_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25625_ net625 _09068_ _09080_ _09074_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__o211a_1
X_22837_ _07314_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29393_ clknet_leaf_259_clock _02406_ VGND VGND VPWR VPWR decode.regfile.registers_4\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28344_ clknet_leaf_203_clock _01357_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25556_ _08931_ _09036_ VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13570_ _09934_ VGND VGND VPWR VPWR _09935_ sky130_fd_sc_hd__buf_4
X_22768_ _07277_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24507_ _08434_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21719_ csr._mcycle_T_2\[30\] _06321_ _06417_ csr.minstret\[30\] VGND VGND VPWR VPWR
+ _06418_ sky130_fd_sc_hd__a211oi_1
X_28275_ clknet_leaf_60_clock _01297_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25487_ net2522 _08995_ _09000_ _08991_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__o211a_1
X_22699_ csr._csr_read_data_T_8\[23\] _07235_ _07238_ _07234_ VGND VGND VPWR VPWR
+ _01307_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15240_ _10657_ _11049_ _11217_ _10662_ VGND VGND VPWR VPWR _11237_ sky130_fd_sc_hd__or4b_2
X_27226_ clknet_leaf_4_clock _00255_ VGND VGND VPWR VPWR decode.regfile.registers_29\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24438_ _08066_ net1335 _08389_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_251_clock clknet_5_18__leaf_clock VGND VGND VPWR VPWR clknet_leaf_251_clock
+ sky130_fd_sc_hd__clkbuf_8
X_27157_ clknet_leaf_355_clock _00186_ VGND VGND VPWR VPWR decode.regfile.registers_27\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_15171_ _10627_ _11091_ _11041_ _11137_ VGND VGND VPWR VPWR _11168_ sky130_fd_sc_hd__and4_1
X_24369_ _08361_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26108_ _09263_ VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__clkbuf_4
X_14122_ net2208 _10288_ _10327_ _10328_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27088_ clknet_leaf_328_clock _00117_ VGND VGND VPWR VPWR decode.regfile.registers_25\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14053_ _10130_ VGND VGND VPWR VPWR _10290_ sky130_fd_sc_hd__clkbuf_4
X_26039_ _08960_ _09310_ VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__nand2_1
X_18930_ _03977_ _03979_ _03982_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__nand3_1
XFILLER_0_162_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_266_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_266_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18861_ decode.id_ex_rs1_data_reg\[10\] _03908_ _04156_ _03700_ _04159_ VGND VGND
+ VPWR VPWR _04160_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_207_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_201_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17812_ decode.regfile.registers_22\[25\] _13100_ _03213_ _13289_ VGND VGND VPWR
+ VPWR _03214_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18792_ decode.id_ex_rs1_data_reg\[15\] _03908_ _04087_ _03914_ _04090_ VGND VGND
+ VPWR VPWR _04091_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_206_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14955_ _10974_ _10982_ VGND VGND VPWR VPWR _10983_ sky130_fd_sc_hd__and2_1
X_29729_ clknet_leaf_289_clock _02742_ VGND VGND VPWR VPWR decode.regfile.registers_15\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_17743_ _12708_ net485 _03110_ _03146_ _03073_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_193_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13906_ _09975_ _10200_ VGND VGND VPWR VPWR _10204_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_193_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17674_ _12138_ _12636_ _12531_ _12728_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__a31o_1
X_14886_ _10618_ VGND VGND VPWR VPWR _10923_ sky130_fd_sc_hd__clkbuf_4
X_19413_ _04443_ _04362_ _04696_ _04701_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__or4b_1
XFILLER_0_212_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13837_ _10008_ _10154_ VGND VGND VPWR VPWR _10163_ sky130_fd_sc_hd__nand2_1
X_16625_ _12497_ _10610_ _10617_ _12488_ VGND VGND VPWR VPWR _12590_ sky130_fd_sc_hd__or4_2
XFILLER_0_98_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_10__f_clock clknet_2_1_0_clock VGND VGND VPWR VPWR clknet_5_10__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_204_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_204_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16556_ _11015_ _10937_ decode.regfile.registers_23\[0\] _12520_ VGND VGND VPWR VPWR
+ _12521_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19344_ _04130_ _04131_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13768_ net2352 _10083_ _10108_ _10077_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15507_ _11371_ decode.regfile.registers_0\[5\] _11155_ _11498_ VGND VGND VPWR VPWR
+ _11499_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_14_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19275_ _04305_ _04372_ _04567_ _04291_ _04568_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__o221a_1
X_16487_ _11263_ decode.regfile.registers_22\[31\] _11404_ _11264_ _11265_ VGND VGND
+ VPWR VPWR _12453_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_85_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13699_ _10021_ memory.io_wb_aluresult\[14\] _10012_ VGND VGND VPWR VPWR _10050_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_152_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18226_ csr.mcycle\[10\] csr.mcycle\[9\] _03559_ _03560_ VGND VGND VPWR VPWR _03561_
+ sky130_fd_sc_hd__and4_1
X_15438_ decode.regfile.registers_23\[3\] _11087_ _11405_ _11431_ VGND VGND VPWR VPWR
+ _11432_ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_219_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_219_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18157_ _03463_ _03464_ _03465_ _10657_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__and4bb_1
X_15369_ _11315_ VGND VGND VPWR VPWR _11364_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17108_ decode.regfile.registers_9\[8\] _10594_ _12690_ _12533_ _13064_ VGND VGND
+ VPWR VPWR _13065_ sky130_fd_sc_hd__a41o_1
Xhold304 decode.id_ex_funct3_reg\[2\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ _03469_ _03467_ _03465_ net1153 VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_106_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold315 decode.regfile.registers_27\[4\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold326 decode.regfile.registers_30\[3\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_229_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold337 decode.regfile.registers_11\[3\] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold348 decode.regfile.registers_16\[9\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_229_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1098 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17039_ _12690_ VGND VGND VPWR VPWR _12998_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_111_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold359 _10063_ VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20050_ decode.id_ex_imm_reg\[7\] decode.id_ex_pc_reg\[7\] VGND VGND VPWR VPWR _05270_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_182_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1004 fetch.bht.bhtTable_target_pc\[15\]\[18\] VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 fetch.bht.bhtTable_tag\[7\]\[1\] VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1026 fetch.bht.bhtTable_target_pc\[1\]\[4\] VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 fetch.bht.bhtTable_tag\[2\]\[16\] VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1048 fetch.bht.bhtTable_tag\[7\]\[16\] VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 fetch.bht.bhtTable_target_pc\[11\]\[11\] VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23740_ _08021_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20952_ _05957_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23671_ _07984_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20883_ _05858_ _09956_ net59 VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25410_ net2385 _08928_ _08949_ _08950_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_81_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22622_ net2530 _07190_ _07191_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__o21a_1
XFILLER_0_192_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26390_ _09533_ VGND VGND VPWR VPWR _09534_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_187_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25341_ _08901_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22553_ csr._minstret_T_3\[35\] csr._minstret_T_3\[34\] _07139_ VGND VGND VPWR VPWR
+ _07143_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_290 _12504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28060_ clknet_leaf_200_clock _01082_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_21504_ _06269_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25272_ _08111_ net2107 _09906_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22484_ fetch.bht.bhtTable_target_pc\[0\]\[0\] fetch.bht.bhtTable_target_pc\[1\]\[0\]
+ fetch.bht.bhtTable_target_pc\[2\]\[0\] fetch.bht.bhtTable_target_pc\[3\]\[0\] _07069_
+ _07072_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__mux4_1
XFILLER_0_185_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27011_ clknet_leaf_341_clock _00040_ VGND VGND VPWR VPWR decode.regfile.registers_22\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24223_ _08051_ net1907 _06241_ VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21435_ _06126_ net1393 _06230_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24154_ _08250_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__clkbuf_1
X_21366_ _06195_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_1056 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23105_ _07545_ _07111_ _07081_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__a21o_1
X_20317_ _05489_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__clkbuf_1
X_28962_ clknet_leaf_134_clock _01975_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_24085_ net1770 execute.io_target_pc\[30\] _07991_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__mux2_1
X_21297_ _06158_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__clkbuf_1
Xhold860 csr._mcycle_T_3\[41\] VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 fetch.bht.bhtTable_tag\[2\]\[14\] VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 csr._mcycle_T_3\[51\] VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__dlygate4sd3_1
X_23036_ fetch.bht.bhtTable_target_pc\[0\]\[8\] fetch.bht.bhtTable_target_pc\[1\]\[8\]
+ fetch.bht.bhtTable_target_pc\[2\]\[8\] fetch.bht.bhtTable_target_pc\[3\]\[8\] _07123_
+ _07101_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__mux4_1
Xhold893 fetch.bht.bhtTable_tag\[10\]\[4\] VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__dlygate4sd3_1
X_27913_ clknet_leaf_66_clock _00942_ VGND VGND VPWR VPWR csr.io_csr_write_address\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20248_ _10704_ _10678_ _05427_ _10730_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__a31o_1
XFILLER_0_229_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28893_ clknet_leaf_177_clock _01906_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20179_ _05369_ _05379_ _05375_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__nand3_1
X_27844_ clknet_leaf_35_clock _00873_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2250 decode.regfile.registers_17\[22\] VGND VGND VPWR VPWR net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2261 decode.regfile.registers_9\[20\] VGND VGND VPWR VPWR net2488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2272 decode.regfile.registers_25\[27\] VGND VGND VPWR VPWR net2499 sky130_fd_sc_hd__dlygate4sd3_1
X_24987_ _08703_ VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__clkbuf_4
Xhold2283 decode.regfile.registers_26\[26\] VGND VGND VPWR VPWR net2510 sky130_fd_sc_hd__dlygate4sd3_1
X_27775_ clknet_leaf_326_clock _00804_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2294 decode.regfile.registers_7\[26\] VGND VGND VPWR VPWR net2521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1560 csr.mcycle\[24\] VGND VGND VPWR VPWR net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1571 fetch.bht.bhtTable_target_pc\[13\]\[11\] VGND VGND VPWR VPWR net1798 sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ _10781_ _10782_ decode.id_ex_pc_reg\[28\] VGND VGND VPWR VPWR _10783_ sky130_fd_sc_hd__o21a_1
X_29514_ clknet_leaf_267_clock _02527_ VGND VGND VPWR VPWR decode.regfile.registers_8\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_23938_ _08139_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__clkbuf_1
X_26726_ _09404_ _09720_ VGND VGND VPWR VPWR _09728_ sky130_fd_sc_hd__nand2_1
Xhold1582 csr.mscratch\[31\] VGND VGND VPWR VPWR net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1593 fetch.bht.bhtTable_target_pc\[14\]\[4\] VGND VGND VPWR VPWR net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14671_ _10687_ decode.id_ex_pc_reg\[27\] execute.io_target_pc\[18\] _10713_ VGND
+ VGND VPWR VPWR _10714_ sky130_fd_sc_hd__o2bb2a_1
X_26657_ _09566_ VGND VGND VPWR VPWR _09688_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_47_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29445_ clknet_leaf_263_clock _02458_ VGND VGND VPWR VPWR decode.regfile.registers_6\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_23869_ _08100_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16410_ _11446_ decode.regfile.registers_28\[28\] _11871_ _11037_ _11448_ VGND VGND
+ VPWR VPWR _12379_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_103_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ memory.csr_read_data_out_reg\[4\] _09942_ _09979_ _09982_ VGND VGND VPWR
+ VPWR _09983_ sky130_fd_sc_hd__a2bb2o_4
X_25608_ _08982_ _09069_ VGND VGND VPWR VPWR _09071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17390_ decode.regfile.registers_15\[15\] _10612_ _10619_ _12589_ _13031_ VGND VGND
+ VPWR VPWR _13340_ sky130_fd_sc_hd__a41o_1
X_29376_ clknet_leaf_256_clock _02389_ VGND VGND VPWR VPWR decode.regfile.registers_4\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26588_ net1837 _09636_ _09647_ _09648_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16341_ _11435_ decode.regfile.registers_24\[27\] _11244_ _11080_ _10991_ VGND VGND
+ VPWR VPWR _12311_ sky130_fd_sc_hd__o2111a_1
X_28327_ clknet_leaf_186_clock _01340_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25539_ _08914_ _09026_ VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__nand2_1
X_13553_ execute.io_mem_rd\[4\] VGND VGND VPWR VPWR _09920_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19060_ _03863_ _04251_ _04252_ _04307_ _04272_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a311o_2
XFILLER_0_109_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_190_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_190_clock
+ sky130_fd_sc_hd__clkbuf_8
X_28258_ clknet_leaf_92_clock _01280_ VGND VGND VPWR VPWR csr._minstret_T_3\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16272_ decode.regfile.registers_2\[25\] _11156_ net348 _11120_ VGND VGND VPWR VPWR
+ _12244_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_81_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27209_ clknet_leaf_363_clock _00238_ VGND VGND VPWR VPWR decode.regfile.registers_28\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15223_ decode.regfile.registers_19\[0\] _11049_ _11215_ _11217_ _11219_ VGND VGND
+ VPWR VPWR _11220_ sky130_fd_sc_hd__o41a_1
X_18011_ net634 _12491_ _12706_ _10940_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28189_ clknet_leaf_85_clock _01211_ VGND VGND VPWR VPWR csr.io_mret_vector\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15154_ _10659_ _10654_ _11150_ VGND VGND VPWR VPWR _11151_ sky130_fd_sc_hd__or3_4
XFILLER_0_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14105_ net2546 _10315_ _10319_ _10317_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19962_ net1214 _03599_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__nor2_1
X_15085_ decode.immGen._imm_T_24\[3\] _10654_ VGND VGND VPWR VPWR _11082_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_201_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14036_ _10117_ _10268_ VGND VGND VPWR VPWR _10279_ sky130_fd_sc_hd__nand2_1
X_18913_ _04197_ _04198_ _04202_ _04207_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_226_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19893_ _03802_ _05128_ _03789_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18844_ _03890_ _04139_ _04140_ _04137_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__o211a_2
XFILLER_0_101_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_220_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18775_ _04070_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_220_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _11199_ _11965_ _11966_ VGND VGND VPWR VPWR _11967_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17726_ decode.regfile.registers_12\[23\] _12542_ _12772_ _12658_ _03129_ VGND VGND
+ VPWR VPWR _03130_ sky130_fd_sc_hd__o311a_1
X_14938_ decode.control.io_opcode\[2\] decode.control.io_opcode\[1\] decode.control.io_opcode\[0\]
+ _10583_ VGND VGND VPWR VPWR _10967_ sky130_fd_sc_hd__and4_1
XFILLER_0_171_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_143_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_143_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17657_ _13250_ decode.regfile.registers_24\[21\] _13170_ _13083_ _13367_ VGND VGND
+ VPWR VPWR _03063_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_77_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14869_ _10577_ _10587_ _10673_ _10911_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__nor4_1
XFILLER_0_148_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16608_ decode.regfile.registers_17\[0\] _12525_ _12569_ _12535_ _12572_ VGND VGND
+ VPWR VPWR _12573_ sky130_fd_sc_hd__a41o_1
XFILLER_0_174_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17588_ net443 _12872_ _13493_ _02995_ _13219_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__o221a_1
XFILLER_0_175_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19327_ _04065_ _04618_ _04445_ _04227_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16539_ _12503_ VGND VGND VPWR VPWR _12504_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_158_clock clknet_5_24__leaf_clock VGND VGND VPWR VPWR clknet_leaf_158_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19258_ _04049_ _04044_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__and2b_1
XFILLER_0_169_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18209_ _10672_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_113_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19189_ _04482_ _04484_ _04268_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21220_ net1498 _06105_ _09912_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_184_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_184_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21151_ _06062_ _06058_ net2531 VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__and3_1
XFILLER_0_229_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold156 io_fetch_data[12] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold167 fetch.bht.bhtTable_valid\[3\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_180_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20102_ decode.id_ex_imm_reg\[15\] _10681_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__nand2_1
Xhold178 execute.csr_write_address_out_reg\[5\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 fetch.btb.btbTable\[8\]\[0\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21082_ execute.csr_read_data_out_reg\[29\] _06025_ _03583_ VGND VGND VPWR VPWR _06028_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_229_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20033_ decode.id_ex_imm_reg\[5\] decode.id_ex_pc_reg\[5\] VGND VGND VPWR VPWR _05255_
+ sky130_fd_sc_hd__nand2_1
X_24910_ csr._mcycle_T_3\[37\] csr._mcycle_T_3\[36\] csr._mcycle_T_3\[35\] _08649_
+ VGND VGND VPWR VPWR _08654_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25890_ net2756 _09226_ _09232_ _09222_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24841_ _08608_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_13 _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27560_ clknet_leaf_55_clock _00589_ VGND VGND VPWR VPWR csr.io_mem_pc\[1\] sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_24 _03369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24772_ _08066_ net1816 _08563_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__mux2_1
XINSDIODE1_35 _08929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21984_ csr._mcycle_T_2\[15\] _06587_ _06595_ _06592_ VGND VGND VPWR VPWR _01235_
+ sky130_fd_sc_hd__o211a_1
XINSDIODE1_46 _09956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26511_ _09415_ _09602_ VGND VGND VPWR VPWR _09604_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_57 _10091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23723_ _08012_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_68 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_205_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20935_ _05948_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__clkbuf_1
XINSDIODE1_79 _10587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27491_ clknet_leaf_31_clock _00520_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29230_ clknet_leaf_123_clock _02243_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26442_ _09424_ _09558_ VGND VGND VPWR VPWR _09564_ sky130_fd_sc_hd__nand2_1
X_23654_ _07975_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20866_ _05910_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29161_ clknet_leaf_205_clock _02174_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_22605_ net2146 _07178_ _07180_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__o21a_1
XFILLER_0_193_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26373_ _09430_ _09515_ VGND VGND VPWR VPWR _09524_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_42_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23585_ _07937_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20797_ net2028 _05867_ _05868_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__and3_1
XFILLER_0_221_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28112_ clknet_leaf_81_clock _01134_ VGND VGND VPWR VPWR csr.minstret\[17\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25324_ _08891_ net2688 VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__and2_1
X_22536_ _07087_ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__buf_8
XFILLER_0_147_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29092_ clknet_leaf_70_clock _02105_ VGND VGND VPWR VPWR csr._mcycle_T_3\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28043_ clknet_leaf_214_clock _01065_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25255_ _08857_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22467_ _06891_ _06893_ _06898_ _07061_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__or4_4
XFILLER_0_63_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24206_ _08277_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__clkbuf_1
X_21418_ _06109_ net1342 _06219_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25186_ _09883_ _10569_ _09881_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__or3b_2
X_22398_ fetch.bht.bhtTable_tag\[12\]\[21\] fetch.bht.bhtTable_tag\[13\]\[21\] _06809_
+ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24137_ net1097 execute.io_target_pc\[23\] _08232_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__mux2_1
X_21349_ _06185_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28945_ clknet_leaf_105_clock _01958_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_24068_ _08206_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__clkbuf_1
Xhold690 fetch.bht.bhtTable_target_pc\[2\]\[0\] VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__dlygate4sd3_1
X_23019_ net227 _07427_ net96 VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__a21oi_1
X_15910_ _11889_ _11890_ _11891_ VGND VGND VPWR VPWR _11892_ sky130_fd_sc_hd__a21o_1
X_28876_ clknet_leaf_87_clock _01889_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16890_ _11019_ _10606_ _10935_ _12649_ VGND VGND VPWR VPWR _12852_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15841_ _10992_ _11066_ _11261_ _11824_ VGND VGND VPWR VPWR _11825_ sky130_fd_sc_hd__a31o_1
X_27827_ clknet_leaf_317_clock _00856_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2080 decode.regfile.registers_13\[20\] VGND VGND VPWR VPWR net2307 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_60_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_60_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold2091 decode.regfile.registers_24\[25\] VGND VGND VPWR VPWR net2318 sky130_fd_sc_hd__dlygate4sd3_1
X_18560_ _03715_ _03725_ _03856_ _03728_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__o31a_1
X_15772_ _11403_ _11754_ _11755_ _11757_ VGND VGND VPWR VPWR _11758_ sky130_fd_sc_hd__a31o_1
X_27758_ clknet_leaf_317_clock _00787_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1390 csr.mcycle\[1\] VGND VGND VPWR VPWR net1617 sky130_fd_sc_hd__dlygate4sd3_1
X_17511_ decode.regfile.registers_3\[18\] _12628_ _12732_ VGND VGND VPWR VPWR _13458_
+ sky130_fd_sc_hd__o21ai_1
X_14723_ csr.io_mem_pc\[19\] csr.io_mem_pc\[20\] csr.io_mem_pc\[21\] _10765_ VGND
+ VGND VPWR VPWR _10766_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26709_ net782 _09709_ _09718_ _09717_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18491_ _03781_ _03788_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__and2_2
X_27689_ clknet_leaf_28_clock _00718_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14654_ decode.id_ex_pc_reg\[29\] VGND VGND VPWR VPWR _10697_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17442_ decode.regfile.registers_10\[16\] _12653_ _13380_ _13390_ VGND VGND VPWR
+ VPWR _13391_ sky130_fd_sc_hd__o22ai_2
X_29428_ clknet_leaf_260_clock _02441_ VGND VGND VPWR VPWR decode.regfile.registers_5\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_75_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_75_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13605_ _09960_ _09961_ memory.io_wb_reg_pc\[2\] VGND VGND VPWR VPWR _09968_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_205_Right_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29359_ clknet_leaf_227_clock _02372_ VGND VGND VPWR VPWR decode.regfile.registers_3\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17373_ decode.regfile.registers_14\[14\] _12669_ _13308_ _13323_ VGND VGND VPWR
+ VPWR _13324_ sky130_fd_sc_hd__o22a_1
X_14585_ _10627_ VGND VGND VPWR VPWR _10628_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_188_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19112_ _04243_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13536_ _09911_ VGND VGND VPWR VPWR _09912_ sky130_fd_sc_hd__buf_4
X_16324_ _11059_ _11149_ _12275_ _12294_ VGND VGND VPWR VPWR _12295_ sky130_fd_sc_hd__o22a_1
XFILLER_0_153_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16255_ decode.regfile.registers_21\[24\] _11267_ _11098_ _11227_ _12227_ VGND VGND
+ VPWR VPWR _12228_ sky130_fd_sc_hd__o311a_1
XFILLER_0_36_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19043_ _04338_ _04339_ _04341_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_42_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15206_ _11202_ VGND VGND VPWR VPWR _11203_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16186_ decode.regfile.registers_20\[22\] _11103_ _11222_ _12160_ VGND VGND VPWR
+ VPWR _12161_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_226_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15137_ _11133_ VGND VGND VPWR VPWR _11134_ sky130_fd_sc_hd__buf_4
XFILLER_0_11_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_13_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_13_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19945_ _05206_ _03627_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__and2_1
X_15068_ _10625_ VGND VGND VPWR VPWR _11065_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14019_ net2169 _10258_ _10269_ _10262_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__o211a_1
X_19876_ _03789_ _03790_ _05120_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_65_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18827_ _03688_ decode.id_ex_rs1_data_reg\[8\] _03700_ _04122_ _04125_ VGND VGND
+ VPWR VPWR _04126_ sky130_fd_sc_hd__o221a_4
Xclkbuf_leaf_28_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_28_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18758_ _04051_ _04054_ _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__or3_1
XFILLER_0_136_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17709_ decode.regfile.registers_17\[23\] _11022_ _12567_ _12586_ VGND VGND VPWR
+ VPWR _03113_ sky130_fd_sc_hd__and4_1
XFILLER_0_172_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18689_ _03984_ _03985_ _03986_ _03987_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20720_ _05804_ _03596_ _05829_ net182 decode.id_ex_rs1_data_reg\[18\] VGND VGND
+ VPWR VPWR _00737_ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20651_ csr.mscratch\[30\] _05591_ _05554_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23370_ fetch.bht.bhtTable_target_pc\[14\]\[28\] fetch.bht.bhtTable_target_pc\[15\]\[28\]
+ _07107_ VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20582_ csr._csr_read_data_T_8\[19\] _05622_ _05718_ _05720_ _05722_ VGND VGND VPWR
+ VPWR _05723_ sky130_fd_sc_hd__a221o_2
XFILLER_0_162_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22321_ _06914_ _06915_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25040_ _03556_ _03561_ net341 VGND VGND VPWR VPWR _08740_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_132_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22252_ _06846_ _06730_ _06686_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21203_ _05867_ _05868_ net2269 VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22183_ fetch.bht.bhtTable_tag\[8\]\[25\] fetch.bht.bhtTable_tag\[9\]\[25\] fetch.bht.bhtTable_tag\[10\]\[25\]
+ fetch.bht.bhtTable_tag\[11\]\[25\] _06619_ _06624_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21134_ _06050_ _06058_ net2358 VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__and3_1
X_26991_ clknet_leaf_334_clock _00020_ VGND VGND VPWR VPWR decode.regfile.registers_22\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28730_ clknet_leaf_178_clock _01743_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25942_ _10130_ VGND VGND VPWR VPWR _09263_ sky130_fd_sc_hd__clkbuf_4
X_21065_ execute.csr_read_data_out_reg\[21\] _06014_ _06010_ VGND VGND VPWR VPWR _06019_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_100_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20016_ decode.id_ex_imm_reg\[3\] _10747_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__or2_1
XFILLER_0_214_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28661_ clknet_leaf_141_clock _01674_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25873_ _09198_ VGND VGND VPWR VPWR _09223_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24824_ _08599_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__clkbuf_1
X_27612_ clknet_leaf_151_clock _00641_ VGND VGND VPWR VPWR execute.io_target_pc\[21\]
+ sky130_fd_sc_hd__dfxtp_4
X_28592_ clknet_leaf_105_clock _01605_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24755_ _08562_ VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__buf_6
X_27543_ clknet_leaf_45_clock _00572_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfxtp_2
X_21967_ net1733 _06572_ _06585_ _06579_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23706_ net1559 _10868_ _08003_ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27474_ clknet_leaf_52_clock _00503_ VGND VGND VPWR VPWR csr.io_csr_address\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20918_ _05939_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_100_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24686_ _08526_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_139_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21898_ _06537_ _06519_ _06520_ _06538_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29213_ clknet_leaf_139_clock _02226_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_23637_ _07966_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__clkbuf_1
X_26425_ net2697 _09548_ _09554_ _09553_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_202_Left_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20849_ _05901_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29144_ clknet_leaf_90_clock _02157_ VGND VGND VPWR VPWR csr.mcycle\[28\] sky130_fd_sc_hd__dfxtp_2
X_26356_ net2033 _09505_ _09514_ _09512_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ net642 _10463_ _10472_ _10468_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__o211a_1
X_23568_ net1871 _07917_ _07928_ _05805_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25307_ _08880_ net2726 VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__and2_1
X_22519_ _06661_ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__buf_4
XFILLER_0_162_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29075_ clknet_leaf_200_clock _02088_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_26287_ _09446_ VGND VGND VPWR VPWR _09475_ sky130_fd_sc_hd__clkbuf_4
X_23499_ _03546_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_190_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _11036_ _11058_ _10632_ VGND VGND VPWR VPWR _12018_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25238_ _08076_ net1684 _08848_ VGND VGND VPWR VPWR _08849_ sky130_fd_sc_hd__mux2_1
X_28026_ clknet_leaf_204_clock _01048_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25169_ _10556_ _10557_ _10568_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__or3b_1
XFILLER_0_62_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_211_Left_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17991_ _12888_ _03386_ _03387_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__o21ai_1
X_19730_ _03888_ _03872_ _04274_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__mux2_1
X_28928_ clknet_leaf_170_clock _01941_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_16942_ _12674_ _12899_ _12902_ VGND VGND VPWR VPWR _12903_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19661_ _04938_ _04939_ _04496_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__and3_1
X_28859_ clknet_leaf_172_clock _01872_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_16873_ _12834_ VGND VGND VPWR VPWR _12835_ sky130_fd_sc_hd__buf_4
XFILLER_0_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18612_ decode.id_ex_rs1_data_reg\[17\] _03908_ _03909_ _03700_ _03910_ VGND VGND
+ VPWR VPWR _03911_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_95_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15824_ _11042_ decode.regfile.registers_4\[13\] _11129_ _10628_ _11082_ VGND VGND
+ VPWR VPWR _11808_ sky130_fd_sc_hd__a2111o_1
X_19592_ _04873_ _04492_ _04508_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18543_ memory.csr_read_data_out_reg\[24\] _09987_ _10104_ _10105_ VGND VGND VPWR
+ VPWR _03842_ sky130_fd_sc_hd__o22a_1
XFILLER_0_158_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15755_ _11046_ decode.regfile.registers_12\[11\] _10649_ _11052_ _10631_ VGND VGND
+ VPWR VPWR _11741_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14706_ execute.io_target_pc\[24\] _10693_ execute.io_target_pc\[3\] _10748_ VGND
+ VGND VPWR VPWR _10749_ sky130_fd_sc_hd__o22a_1
X_18474_ decode.id_ex_islui_reg VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_220_Left_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15686_ _11079_ _11244_ _11261_ _11647_ _11673_ VGND VGND VPWR VPWR _11674_ sky130_fd_sc_hd__a41o_1
XFILLER_0_47_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _13221_ _13372_ _13373_ _13374_ VGND VGND VPWR VPWR _13375_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_215_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14637_ decode.id_ex_pc_reg\[8\] VGND VGND VPWR VPWR _10680_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17356_ _11021_ _12559_ _12534_ _13031_ decode.regfile.registers_16\[14\] VGND VGND
+ VPWR VPWR _13307_ sky130_fd_sc_hd__a32o_1
X_14568_ _10610_ VGND VGND VPWR VPWR _10611_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16307_ decode.regfile.registers_7\[26\] _11378_ _11170_ decode.regfile.registers_6\[26\]
+ _11281_ VGND VGND VPWR VPWR _12278_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_83_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13519_ _09897_ VGND VGND VPWR VPWR _09898_ sky130_fd_sc_hd__buf_4
XFILLER_0_166_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17287_ decode.regfile.registers_15\[12\] _12666_ _12723_ _12575_ VGND VGND VPWR
+ VPWR _13240_ sky130_fd_sc_hd__o31a_1
XFILLER_0_43_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14499_ _10426_ VGND VGND VPWR VPWR _10546_ sky130_fd_sc_hd__buf_4
XFILLER_0_113_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19026_ _04324_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__clkbuf_4
X_16238_ _11156_ _12209_ _12210_ VGND VGND VPWR VPWR _12211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16169_ decode.regfile.registers_5\[22\] _10637_ _11139_ _12142_ _12143_ VGND VGND
+ VPWR VPWR _12144_ sky130_fd_sc_hd__a32o_1
XFILLER_0_140_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19928_ _04443_ _04620_ _05195_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_208_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19859_ _05128_ net212 _05129_ _04444_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__a31o_1
XFILLER_0_223_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22870_ _07331_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21821_ _06481_ csr.io_ecause\[0\] _06316_ _06470_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24540_ _08451_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21752_ _06438_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_121_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20703_ _05804_ _03596_ _05819_ net183 net2725 VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__a32o_1
X_24471_ _08415_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21683_ net843 _06387_ _06388_ _06352_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26210_ _09426_ _09413_ VGND VGND VPWR VPWR _09427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23422_ csr._csr_read_data_T_8\[31\] _07416_ csr.io_mret_vector\[31\] _07417_ _07843_
+ VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__o221a_1
X_20634_ csr.minstret\[27\] _05573_ _05585_ csr.mcycle\[27\] VGND VGND VPWR VPWR _05767_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27190_ clknet_leaf_353_clock _00219_ VGND VGND VPWR VPWR decode.regfile.registers_28\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26141_ net2257 _09373_ _09378_ _09370_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__o211a_1
X_23353_ fetch.bht.bhtTable_target_pc\[0\]\[27\] fetch.bht.bhtTable_target_pc\[1\]\[27\]
+ fetch.bht.bhtTable_target_pc\[2\]\[27\] fetch.bht.bhtTable_target_pc\[3\]\[27\]
+ _07708_ _07710_ VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20565_ csr.minstret\[17\] _05594_ _05595_ csr._minstret_T_3\[49\] VGND VGND VPWR
+ VPWR _05708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22304_ fetch.bht.bhtTable_tag\[4\]\[0\] fetch.bht.bhtTable_tag\[5\]\[0\] _06878_
+ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26072_ _08918_ _09330_ VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__nand2_1
X_23284_ execute.io_target_pc\[22\] _07090_ _06041_ _06038_ VGND VGND VPWR VPWR _07715_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20496_ csr.minstret\[8\] _05572_ _05582_ csr.mcycle\[8\] VGND VGND VPWR VPWR _05648_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25023_ csr._mcycle_T_2\[12\] _08704_ csr.mcycle\[12\] VGND VGND VPWR VPWR _08729_
+ sky130_fd_sc_hd__a21oi_1
X_29900_ clknet_leaf_301_clock _02913_ VGND VGND VPWR VPWR decode.regfile.registers_20\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_22235_ _06623_ _06827_ _06673_ _06829_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29831_ clknet_leaf_298_clock _02844_ VGND VGND VPWR VPWR decode.regfile.registers_18\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_22166_ fetch.bht.bhtTable_tag\[12\]\[13\] fetch.bht.bhtTable_tag\[13\]\[13\] _06680_
+ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21117_ _06050_ _06046_ net648 VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__and3_1
X_29762_ clknet_leaf_291_clock _02775_ VGND VGND VPWR VPWR decode.regfile.registers_16\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22097_ fetch.bht.bhtTable_tag\[12\]\[7\] fetch.bht.bhtTable_tag\[13\]\[7\] _06691_
+ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__mux2_1
X_26974_ net2457 _09866_ _09870_ _09865_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28713_ clknet_leaf_88_clock _01726_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21048_ _06009_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__clkbuf_1
X_25925_ _09241_ VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__clkbuf_4
X_29693_ clknet_leaf_290_clock _02706_ VGND VGND VPWR VPWR decode.regfile.registers_14\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28644_ clknet_leaf_132_clock _01657_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13870_ _10092_ _10177_ VGND VGND VPWR VPWR _10182_ sky130_fd_sc_hd__nand2_1
X_25856_ _08929_ _09210_ VGND VGND VPWR VPWR _09214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24807_ _08590_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__clkbuf_1
X_28575_ clknet_leaf_189_clock _01588_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_22999_ _07097_ _07438_ _07443_ _07445_ VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__a2bb2o_2
X_25787_ _08935_ _09166_ VGND VGND VPWR VPWR _09174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_213_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27526_ clknet_leaf_44_clock _00555_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfxtp_2
XINSDIODE1_108 _10935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15540_ decode.regfile.registers_14\[6\] _11207_ _11273_ decode.regfile.registers_15\[6\]
+ _11201_ VGND VGND VPWR VPWR _11531_ sky130_fd_sc_hd__a221o_1
X_24738_ _08553_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_119 _11058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15471_ decode.regfile.registers_5\[4\] _10637_ _11139_ _11461_ _11463_ VGND VGND
+ VPWR VPWR _11464_ sky130_fd_sc_hd__a32o_1
X_24669_ net1618 execute.io_target_pc\[23\] _08508_ VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__mux2_1
X_27457_ clknet_leaf_137_clock _00486_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17210_ decode.regfile.registers_21\[10\] _12681_ VGND VGND VPWR VPWR _13165_ sky130_fd_sc_hd__or2_1
X_14422_ net476 _10490_ _10501_ _10494_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__o211a_1
X_26408_ net655 _09534_ _09544_ _09540_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18190_ decode.control.io_funct3\[2\] decode.control.io_funct3\[0\] VGND VGND VPWR
+ VPWR _03528_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27388_ clknet_leaf_10_clock _00417_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_29127_ clknet_leaf_76_clock _02140_ VGND VGND VPWR VPWR csr.mcycle\[11\] sky130_fd_sc_hd__dfxtp_2
X_14353_ _10461_ VGND VGND VPWR VPWR _10462_ sky130_fd_sc_hd__clkbuf_4
X_17141_ _12486_ VGND VGND VPWR VPWR _13097_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26339_ _09490_ VGND VGND VPWR VPWR _09505_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17072_ _12666_ _12723_ _12984_ decode.regfile.registers_14\[7\] _13029_ VGND VGND
+ VPWR VPWR _13030_ sky130_fd_sc_hd__o221ai_1
X_29058_ clknet_leaf_213_clock _02071_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14284_ _09970_ _10420_ VGND VGND VPWR VPWR _10423_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28009_ clknet_leaf_191_clock _01031_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_16023_ decode.regfile.registers_16\[18\] _11359_ _11986_ _12001_ _11126_ VGND VGND
+ VPWR VPWR _12002_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_208_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17974_ _12967_ _03369_ _03370_ _03371_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19713_ _04599_ _04600_ _04728_ _04805_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__o211a_1
X_16925_ _10610_ _12615_ _12629_ decode.regfile.registers_3\[4\] _12885_ VGND VGND
+ VPWR VPWR _12886_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_204_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_108_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19644_ _04299_ _04424_ _04056_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__or3_2
X_16856_ _12496_ _12816_ _12817_ _12818_ VGND VGND VPWR VPWR _12819_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_196_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15807_ _11075_ _11790_ _11791_ _11486_ VGND VGND VPWR VPWR _11792_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_217_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19575_ _04844_ _04845_ _04854_ _04857_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_217_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16787_ decode.regfile.registers_16\[1\] _12575_ _12720_ _12750_ VGND VGND VPWR VPWR
+ _12751_ sky130_fd_sc_hd__o22a_1
X_13999_ _10242_ VGND VGND VPWR VPWR _10258_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18526_ _03709_ decode.id_ex_imm_reg\[27\] _03824_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15738_ _10994_ VGND VGND VPWR VPWR _11724_ sky130_fd_sc_hd__buf_2
XFILLER_0_220_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18457_ execute.io_mem_rd\[3\] _03755_ execute.io_mem_rd\[0\] _03721_ VGND VGND VPWR
+ VPWR _03756_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15669_ _11313_ decode.regfile.registers_4\[9\] VGND VGND VPWR VPWR _11657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17408_ decode.regfile.registers_16\[15\] _13011_ _13340_ _13357_ VGND VGND VPWR
+ VPWR _13358_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_146_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18388_ _03686_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__buf_6
XFILLER_0_117_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17339_ _13081_ _13168_ decode.regfile.registers_23\[13\] _13041_ VGND VGND VPWR
+ VPWR _13291_ sky130_fd_sc_hd__or4_1
XFILLER_0_154_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20350_ decode.id_ex_pc_reg\[28\] _10697_ decode.id_ex_pc_reg\[30\] _05502_ VGND
+ VGND VPWR VPWR _05514_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19009_ _03637_ _03633_ _03635_ _03634_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__or4b_2
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20281_ _10694_ _10710_ decode.id_ex_pc_reg\[14\] _05452_ VGND VGND VPWR VPWR _05462_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22020_ _00000_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__buf_8
XFILLER_0_109_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Left_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1901 decode.regfile.registers_2\[4\] VGND VGND VPWR VPWR net2128 sky130_fd_sc_hd__dlygate4sd3_1
X_23971_ _08156_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_127_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1912 fetch.bht.bhtTable_target_pc\[10\]\[12\] VGND VGND VPWR VPWR net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1923 fetch.bht.bhtTable_tag\[8\]\[5\] VGND VGND VPWR VPWR net2150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 fetch.bht.bhtTable_target_pc\[7\]\[28\] VGND VGND VPWR VPWR net2161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22922_ fetch.bht.bhtTable_target_pc\[12\]\[2\] fetch.bht.bhtTable_target_pc\[13\]\[2\]
+ _07068_ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__mux2_1
Xhold1945 decode.regfile.registers_10\[19\] VGND VGND VPWR VPWR net2172 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25710_ _08933_ _09122_ VGND VGND VPWR VPWR _09130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1956 decode.regfile.registers_15\[18\] VGND VGND VPWR VPWR net2183 sky130_fd_sc_hd__dlygate4sd3_1
X_26690_ net2600 _09666_ _09706_ _09702_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_123_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1967 decode.regfile.registers_10\[5\] VGND VGND VPWR VPWR net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1978 fetch.bht.bhtTable_tag\[7\]\[2\] VGND VGND VPWR VPWR net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1989 fetch.bht.bhtTable_tag\[7\]\[13\] VGND VGND VPWR VPWR net2216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22853_ _07322_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25641_ net1874 _09082_ _09089_ _09087_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21804_ csr.io_csr_write_address\[6\] _06469_ _06458_ VGND VGND VPWR VPWR _06472_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_17_1321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28360_ clknet_leaf_236_clock _01373_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25572_ _08945_ _09049_ VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__nand2_1
X_22784_ net1185 _10820_ _07286_ VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24523_ _08083_ net1210 _08439_ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__mux2_1
X_27311_ clknet_leaf_239_clock _00340_ VGND VGND VPWR VPWR fetch.btb.btbTable\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21735_ net1067 _10821_ _06428_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28291_ clknet_leaf_85_clock _01313_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_135_Left_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24454_ _08406_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__clkbuf_1
X_27242_ clknet_leaf_0_clock _00271_ VGND VGND VPWR VPWR decode.regfile.registers_29\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21666_ csr._mcycle_T_2\[19\] _06321_ _06375_ csr.minstret\[19\] VGND VGND VPWR VPWR
+ _06376_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_97_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23405_ csr._csr_read_data_T_8\[30\] _07416_ csr.io_mret_vector\[30\] _07417_ _07827_
+ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__o221a_1
XFILLER_0_35_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20617_ csr.mscratch\[24\] _05593_ _05625_ _05751_ _05752_ VGND VGND VPWR VPWR _05753_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27173_ clknet_leaf_362_clock _00202_ VGND VGND VPWR VPWR decode.regfile.registers_27\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_24385_ net938 execute.io_target_pc\[15\] _08367_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__mux2_1
X_21597_ _06320_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_10_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26124_ _08970_ _09328_ VGND VGND VPWR VPWR _09367_ sky130_fd_sc_hd__nand2_1
X_23336_ fetch.bht.bhtTable_target_pc\[12\]\[26\] fetch.bht.bhtTable_target_pc\[13\]\[26\]
+ fetch.bht.bhtTable_target_pc\[14\]\[26\] fetch.bht.bhtTable_target_pc\[15\]\[26\]
+ _07669_ _07656_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__mux4_1
XFILLER_0_163_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20548_ _05591_ csr.io_mret_vector\[15\] _05565_ _05692_ VGND VGND VPWR VPWR _05693_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26055_ _09930_ _10194_ _09932_ _08902_ VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__and4b_1
X_23267_ fetch.bht.bhtTable_target_pc\[8\]\[21\] fetch.bht.bhtTable_target_pc\[9\]\[21\]
+ fetch.bht.bhtTable_target_pc\[10\]\[21\] fetch.bht.bhtTable_target_pc\[11\]\[21\]
+ _07098_ _07113_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20479_ csr.minstret\[6\] _05574_ _05586_ csr.mcycle\[6\] VGND VGND VPWR VPWR _05633_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25006_ _08716_ _08717_ _08704_ VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__a21o_1
X_22218_ _06691_ fetch.bht.bhtTable_tag\[10\]\[20\] VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23198_ _06887_ _07536_ _07537_ _07633_ _07535_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_144_Left_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29814_ clknet_leaf_296_clock _02827_ VGND VGND VPWR VPWR decode.regfile.registers_17\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22149_ fetch.bht.bhtTable_tag\[4\]\[23\] fetch.bht.bhtTable_tag\[5\]\[23\] _06618_
+ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29745_ clknet_leaf_294_clock _02758_ VGND VGND VPWR VPWR decode.regfile.registers_15\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14971_ _10974_ _10995_ VGND VGND VPWR VPWR _10996_ sky130_fd_sc_hd__and2_1
X_26957_ net802 _09853_ _09860_ _09852_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__o211a_1
X_16710_ decode.regfile.registers_15\[0\] _12585_ _12665_ _12671_ _12674_ VGND VGND
+ VPWR VPWR _12675_ sky130_fd_sc_hd__a221o_1
X_13922_ _10198_ VGND VGND VPWR VPWR _10213_ sky130_fd_sc_hd__buf_2
X_25908_ _09025_ _09243_ VGND VGND VPWR VPWR _09244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17690_ _03076_ _03094_ _12565_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__o21a_1
X_29676_ clknet_leaf_282_clock _02689_ VGND VGND VPWR VPWR decode.regfile.registers_13\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26888_ _09415_ _09819_ VGND VGND VPWR VPWR _09821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28627_ clknet_leaf_140_clock _01640_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16641_ _12605_ VGND VGND VPWR VPWR _12606_ sky130_fd_sc_hd__clkbuf_4
X_13853_ _10053_ _10164_ VGND VGND VPWR VPWR _10172_ sky130_fd_sc_hd__nand2_1
X_25839_ _08912_ _09200_ VGND VGND VPWR VPWR _09204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19360_ _04465_ _04645_ _04428_ _04650_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__a2bb2o_1
X_28558_ clknet_leaf_165_clock _01571_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16572_ _12536_ VGND VGND VPWR VPWR _12537_ sky130_fd_sc_hd__buf_2
XFILLER_0_201_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13784_ net195 VGND VGND VPWR VPWR _10122_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_153_Left_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18311_ decode.id_ex_rs2_data_reg\[21\] _03616_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_191_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _10651_ _11111_ _11118_ _11514_ VGND VGND VPWR VPWR _11515_ sky130_fd_sc_hd__a31o_1
X_27509_ clknet_leaf_9_clock _00538_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_191_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19291_ _04552_ _04580_ _04561_ _04454_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__o31a_1
X_28489_ clknet_leaf_194_clock _01502_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18242_ csr._mcycle_T_3\[41\] csr._mcycle_T_3\[40\] csr._mcycle_T_3\[39\] csr._mcycle_T_3\[38\]
+ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__or4_1
XFILLER_0_155_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15454_ _11349_ VGND VGND VPWR VPWR _11447_ sky130_fd_sc_hd__buf_2
XFILLER_0_155_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14405_ net668 _10490_ _10492_ _10481_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18173_ _03514_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15385_ _11136_ _11377_ _11379_ VGND VGND VPWR VPWR _11380_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17124_ _11013_ VGND VGND VPWR VPWR _13081_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14336_ _10426_ VGND VGND VPWR VPWR _10453_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap205 _03698_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_6
Xmax_cap216 net352 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__buf_1
Xhold508 _06489_ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold519 csr.minstret\[25\] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17055_ decode.regfile.registers_2\[7\] _10608_ net215 net209 VGND VGND VPWR VPWR
+ _13013_ sky130_fd_sc_hd__a31o_1
X_14267_ net874 _10403_ _10412_ _10411_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Left_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16006_ _11493_ decode.regfile.registers_22\[18\] _11450_ _10979_ _10991_ VGND VGND
+ VPWR VPWR _11985_ sky130_fd_sc_hd__o2111a_1
X_14198_ _10147_ _10331_ VGND VGND VPWR VPWR _10372_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_206_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_198_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 fetch.bht.bhtTable_tag\[11\]\[1\] VGND VGND VPWR VPWR net1435 sky130_fd_sc_hd__dlygate4sd3_1
X_17957_ _11019_ _12489_ _12511_ decode.regfile.registers_12\[29\] _12745_ VGND VGND
+ VPWR VPWR _03355_ sky130_fd_sc_hd__o32a_1
Xhold1219 csr.mscratch\[5\] VGND VGND VPWR VPWR net1446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16908_ _12496_ _12867_ _12868_ _12869_ VGND VGND VPWR VPWR _12870_ sky130_fd_sc_hd__a31o_1
X_17888_ decode.regfile.registers_20\[27\] _12770_ _03287_ _12537_ VGND VGND VPWR
+ VPWR _03288_ sky130_fd_sc_hd__a211o_1
XFILLER_0_206_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19627_ _04503_ _04203_ _04445_ _03902_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__and4_1
XFILLER_0_219_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16839_ _12580_ _12800_ _12801_ VGND VGND VPWR VPWR _12802_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19558_ _04840_ _04211_ _04452_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_220_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_215_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18509_ decode.id_ex_rs2_data_reg\[26\] _03747_ _03805_ _03759_ _03727_ VGND VGND
+ VPWR VPWR _03808_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19489_ _04304_ _03704_ _04537_ _04573_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__o2bb2a_1
X_21520_ _06149_ net1750 _06274_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21451_ _06217_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_185_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20402_ _03718_ _05516_ net358 _03737_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__or4_2
X_24170_ _08064_ net1740 _08255_ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21382_ _06130_ net1878 _06199_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23121_ fetch.bht.bhtTable_target_pc\[2\]\[13\] fetch.bht.bhtTable_target_pc\[3\]\[13\]
+ _07119_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20333_ _05420_ _05384_ _05501_ _05454_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23052_ _07085_ _07491_ _07495_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_222_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20264_ _10706_ decode.id_ex_pc_reg\[10\] _05440_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_129_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22003_ net723 _06600_ _06606_ _06605_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__o211a_1
X_27860_ clknet_leaf_318_clock _00889_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_20195_ decode.id_ex_imm_reg\[28\] decode.id_ex_pc_reg\[28\] VGND VGND VPWR VPWR
+ _05394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2410 decode.regfile.registers_24\[30\] VGND VGND VPWR VPWR net2637 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2421 csr.minstret\[17\] VGND VGND VPWR VPWR net2648 sky130_fd_sc_hd__dlygate4sd3_1
X_26811_ _09412_ _09776_ VGND VGND VPWR VPWR _09777_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2432 decode.regfile.registers_9\[5\] VGND VGND VPWR VPWR net2659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2443 execute.io_mem_isbranch VGND VGND VPWR VPWR net2670 sky130_fd_sc_hd__dlygate4sd3_1
X_27791_ clknet_leaf_305_clock _00820_ VGND VGND VPWR VPWR memory.io_wb_readdata\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2454 decode.regfile.registers_16\[26\] VGND VGND VPWR VPWR net2681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1720 csr.mcycle\[27\] VGND VGND VPWR VPWR net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2465 csr._csr_read_data_T_8\[20\] VGND VGND VPWR VPWR net2692 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29530_ clknet_leaf_313_clock _02543_ VGND VGND VPWR VPWR decode.regfile.registers_9\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1731 _01247_ VGND VGND VPWR VPWR net1958 sky130_fd_sc_hd__dlygate4sd3_1
X_26742_ net2109 _09736_ _09737_ _09730_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__o211a_1
Xhold2476 decode.regfile.registers_10\[22\] VGND VGND VPWR VPWR net2703 sky130_fd_sc_hd__dlygate4sd3_1
X_23954_ _08147_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__clkbuf_1
Xhold1742 fetch.bht.bhtTable_tag\[0\]\[2\] VGND VGND VPWR VPWR net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2487 decode.regfile.registers_9\[31\] VGND VGND VPWR VPWR net2714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1753 fetch.bht.bhtTable_target_pc\[7\]\[8\] VGND VGND VPWR VPWR net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2498 decode.id_ex_rs1_data_reg\[11\] VGND VGND VPWR VPWR net2725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1764 decode.regfile.registers_19\[23\] VGND VGND VPWR VPWR net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1775 fetch.bht.bhtTable_tag\[13\]\[3\] VGND VGND VPWR VPWR net2002 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22905_ net90 _06806_ _06670_ net221 _07355_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_4_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29461_ clknet_leaf_264_clock _02474_ VGND VGND VPWR VPWR decode.regfile.registers_6\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1786 fetch.bht.bhtTable_tag\[15\]\[18\] VGND VGND VPWR VPWR net2013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23885_ execute.io_target_pc\[30\] VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__buf_2
X_26673_ _09428_ _09689_ VGND VGND VPWR VPWR _09697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1797 decode.io_id_pc\[6\] VGND VGND VPWR VPWR net2024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28412_ clknet_leaf_143_clock _01425_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_168_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22836_ net1636 csr.io_mem_pc\[31\] _07308_ VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__mux2_1
X_25624_ _08922_ _09079_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29392_ clknet_leaf_259_clock _02405_ VGND VGND VPWR VPWR decode.regfile.registers_4\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28343_ clknet_leaf_210_clock _01356_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22767_ _06140_ net1273 _07276_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_870 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25555_ net618 _09039_ _09040_ _09033_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24506_ _08066_ net1682 _08428_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__mux2_1
X_21718_ csr.minstret\[28\] csr.minstret\[29\] _06413_ VGND VGND VPWR VPWR _06417_
+ sky130_fd_sc_hd__and3_2
X_28274_ clknet_leaf_60_clock _01296_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_25486_ _08937_ _08992_ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22698_ net723 _07236_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27225_ clknet_leaf_4_clock _00254_ VGND VGND VPWR VPWR decode.regfile.registers_29\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24437_ _08397_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__clkbuf_1
X_21649_ csr._mcycle_T_2\[14\] _06325_ _06358_ csr.minstret\[13\] csr.minstret\[14\]
+ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_192_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15170_ _11142_ VGND VGND VPWR VPWR _11167_ sky130_fd_sc_hd__buf_4
X_24368_ net1353 execute.io_target_pc\[7\] _08356_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__mux2_1
X_27156_ clknet_leaf_353_clock _00185_ VGND VGND VPWR VPWR decode.regfile.registers_27\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_90 decode.id_ex_rs2_data_reg\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14121_ _10290_ VGND VGND VPWR VPWR _10328_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23319_ net220 _07740_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26107_ _08954_ _09353_ VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27087_ clknet_leaf_329_clock _00116_ VGND VGND VPWR VPWR decode.regfile.registers_25\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24299_ _08325_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14052_ _09950_ _10288_ VGND VGND VPWR VPWR _10289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26038_ net2586 _09313_ _09317_ _09318_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18860_ _03816_ _04158_ net353 VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17811_ decode.regfile.registers_21\[25\] _12716_ _03186_ _03212_ _13164_ VGND VGND
+ VPWR VPWR _03213_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_201_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18791_ _03816_ _04089_ _03774_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_201_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27989_ clknet_leaf_217_clock _01011_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17742_ _02997_ _13262_ _12965_ decode.regfile.registers_29\[23\] _03145_ VGND VGND
+ VPWR VPWR _03146_ sky130_fd_sc_hd__o221a_1
X_29728_ clknet_leaf_311_clock _02741_ VGND VGND VPWR VPWR decode.regfile.registers_15\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14954_ decode.immGen._imm_T_10\[1\] _10948_ _10975_ _10981_ VGND VGND VPWR VPWR
+ _10982_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13905_ net1374 _10199_ _10203_ _10188_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_193_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17673_ _12636_ _13145_ decode.regfile.registers_0\[22\] VGND VGND VPWR VPWR _03078_
+ sky130_fd_sc_hd__a21oi_1
X_29659_ clknet_leaf_271_clock _02672_ VGND VGND VPWR VPWR decode.regfile.registers_13\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_193_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14885_ _10922_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__clkbuf_1
X_19412_ _04371_ _04421_ _04633_ _04700_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__a211o_1
X_16624_ _12588_ VGND VGND VPWR VPWR _12589_ sky130_fd_sc_hd__clkbuf_4
X_13836_ net1030 _10153_ _10161_ _10162_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19343_ _04515_ _04610_ _04632_ _04634_ _03595_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16555_ _12519_ VGND VGND VPWR VPWR _12520_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13767_ _10107_ _10075_ VGND VGND VPWR VPWR _10108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15506_ decode.regfile.registers_1\[5\] _11115_ _11056_ _11108_ VGND VGND VPWR VPWR
+ _11498_ sky130_fd_sc_hd__and4_1
X_19274_ _04243_ _04541_ _04378_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__or3b_1
XFILLER_0_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16486_ _11435_ decode.regfile.registers_24\[31\] _11065_ _11080_ _10991_ VGND VGND
+ VPWR VPWR _12452_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_57_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13698_ net838 _10027_ _10049_ _10020_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18225_ csr.mcycle\[12\] csr.mcycle\[11\] csr.mcycle\[13\] VGND VGND VPWR VPWR _03560_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_150_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15437_ decode.regfile.registers_21\[3\] _11267_ _11099_ _11228_ _11430_ VGND VGND
+ VPWR VPWR _11431_ sky130_fd_sc_hd__o311a_1
XFILLER_0_84_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18156_ _11067_ _10577_ _10673_ _10911_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__nor4_1
XFILLER_0_5_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15368_ decode.regfile.registers_11\[2\] _11071_ _11204_ _11187_ VGND VGND VPWR VPWR
+ _11363_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_170_Left_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17107_ decode.regfile.registers_8\[8\] _12726_ _13057_ _13063_ _12602_ VGND VGND
+ VPWR VPWR _13064_ sky130_fd_sc_hd__o221a_1
XFILLER_0_80_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14319_ _10069_ _10431_ VGND VGND VPWR VPWR _10443_ sky130_fd_sc_hd__nand2_1
Xhold305 decode.regfile.registers_29\[0\] VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ _10575_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold316 decode.regfile.registers_30\[24\] VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15299_ _10627_ _11107_ _11041_ _11055_ VGND VGND VPWR VPWR _11295_ sky130_fd_sc_hd__nand4_4
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold327 decode.regfile.registers_29\[11\] VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold338 decode.regfile.registers_23\[15\] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold349 fetch.bht.bhtTable_valid\[8\] VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ _10604_ VGND VGND VPWR VPWR _12997_ sky130_fd_sc_hd__buf_2
XFILLER_0_150_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_182_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _04281_ _04283_ _04249_ _04284_ _04287_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1005 fetch.bht.bhtTable_tag\[9\]\[16\] VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 fetch.bht.bhtTable_target_pc\[13\]\[22\] VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 fetch.bht.bhtTable_target_pc\[12\]\[2\] VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1038 decode.regfile.registers_14\[10\] VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 fetch.bht.bhtTable_target_pc\[2\]\[18\] VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_219_Right_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20951_ execute.io_reg_pc\[2\] _05915_ _05911_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_85_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23670_ net2125 _10760_ _07983_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_311_clock clknet_5_18__leaf_clock VGND VGND VPWR VPWR clknet_leaf_311_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20882_ _05919_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22621_ csr._minstret_T_3\[55\] _07190_ _07179_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_81_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25340_ _08891_ net2755 VGND VGND VPWR VPWR _08901_ sky130_fd_sc_hd__and2_1
X_22552_ csr._minstret_T_3\[34\] _07139_ net2323 VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_118_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_280 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21503_ _06132_ net1085 _06263_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_291 _12504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25271_ _08865_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_326_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_326_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22483_ fetch.bht.bhtTable_target_pc\[4\]\[0\] fetch.bht.bhtTable_target_pc\[5\]\[0\]
+ fetch.bht.bhtTable_target_pc\[6\]\[0\] fetch.bht.bhtTable_target_pc\[7\]\[0\] _07069_
+ _07072_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__mux4_1
XFILLER_0_174_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24222_ _08285_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27010_ clknet_leaf_341_clock _00039_ VGND VGND VPWR VPWR decode.regfile.registers_22\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21434_ _06232_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24153_ net990 execute.io_target_pc\[31\] _06427_ VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21365_ _06113_ net1831 _06188_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23104_ fetch.bht.bhtTable_target_pc\[14\]\[12\] fetch.bht.bhtTable_target_pc\[15\]\[12\]
+ _07119_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20316_ _05439_ _05488_ _05425_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__and3b_1
XFILLER_0_82_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24084_ _08214_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__clkbuf_1
X_28961_ clknet_leaf_175_clock _01974_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold850 fetch.bht.bhtTable_tag\[7\]\[0\] VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__dlygate4sd3_1
X_21296_ net1661 _06101_ _06157_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__mux2_1
Xhold861 decode.regfile.registers_27\[19\] VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23035_ fetch.bht.bhtTable_target_pc\[4\]\[8\] fetch.bht.bhtTable_target_pc\[5\]\[8\]
+ fetch.bht.bhtTable_target_pc\[6\]\[8\] fetch.bht.bhtTable_target_pc\[7\]\[8\] _07123_
+ _07101_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__mux4_1
X_27912_ clknet_leaf_23_clock _00941_ VGND VGND VPWR VPWR csr.io_csr_write_address\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold872 decode.regfile.registers_6\[31\] VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 fetch.bht.bhtTable_tag\[14\]\[21\] VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__dlygate4sd3_1
X_20247_ _05412_ _05266_ _05435_ _03517_ _03551_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__a2111oi_1
X_28892_ clknet_leaf_182_clock _01905_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold894 decode.control.io_funct7\[5\] VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__dlygate4sd3_1
X_27843_ clknet_leaf_35_clock _00872_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20178_ decode.id_ex_imm_reg\[23\] _10786_ _05371_ _05365_ _05370_ VGND VGND VPWR
+ VPWR _05379_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_216_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2240 decode.regfile.registers_26\[23\] VGND VGND VPWR VPWR net2467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2251 decode.regfile.registers_27\[16\] VGND VGND VPWR VPWR net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2262 decode.regfile.registers_31\[0\] VGND VGND VPWR VPWR net2489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2273 decode.regfile.registers_18\[1\] VGND VGND VPWR VPWR net2500 sky130_fd_sc_hd__dlygate4sd3_1
X_27774_ clknet_leaf_326_clock _00803_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24986_ csr.io_csr_write_address\[11\] net216 _06314_ _06459_ VGND VGND VPWR VPWR
+ _08703_ sky130_fd_sc_hd__and4_2
Xhold2284 decode.regfile.registers_11\[13\] VGND VGND VPWR VPWR net2511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1550 fetch.bht.bhtTable_target_pc\[0\]\[3\] VGND VGND VPWR VPWR net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2295 decode.regfile.registers_2\[14\] VGND VGND VPWR VPWR net2522 sky130_fd_sc_hd__dlygate4sd3_1
X_29513_ clknet_leaf_265_clock _02526_ VGND VGND VPWR VPWR decode.regfile.registers_8\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1561 fetch.bht.bhtTable_target_pc\[5\]\[25\] VGND VGND VPWR VPWR net1788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26725_ net639 _09723_ _09727_ _09717_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23937_ net1072 _08095_ _08130_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__mux2_1
Xhold1572 fetch.bht.bhtTable_target_pc\[10\]\[28\] VGND VGND VPWR VPWR net1799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1583 decode.io_mret_out VGND VGND VPWR VPWR net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1594 fetch.bht.bhtTable_tag\[4\]\[5\] VGND VGND VPWR VPWR net1821 sky130_fd_sc_hd__dlygate4sd3_1
X_29444_ clknet_leaf_262_clock _02457_ VGND VGND VPWR VPWR decode.regfile.registers_6\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14670_ decode.id_ex_pc_reg\[18\] VGND VGND VPWR VPWR _10713_ sky130_fd_sc_hd__inv_2
X_26656_ _09410_ _09676_ VGND VGND VPWR VPWR _09687_ sky130_fd_sc_hd__nand2_1
X_23868_ _08099_ net1537 _07940_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13621_ _09943_ memory.io_wb_aluresult\[4\] _09981_ memory.io_wb_readdata\[4\] _09977_
+ VGND VGND VPWR VPWR _09982_ sky130_fd_sc_hd__a221oi_2
X_25607_ net707 _09068_ _09070_ _09059_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__o211a_1
X_22819_ net692 csr.io_mem_pc\[23\] _07297_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29375_ clknet_leaf_255_clock _02388_ VGND VGND VPWR VPWR decode.regfile.registers_4\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26587_ _09566_ VGND VGND VPWR VPWR _09648_ sky130_fd_sc_hd__buf_2
X_23799_ execute.io_target_pc\[2\] VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__buf_2
XFILLER_0_196_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28326_ clknet_leaf_191_clock _01339_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_16340_ _11346_ decode.regfile.registers_30\[27\] _12095_ _12096_ _12097_ VGND VGND
+ VPWR VPWR _12310_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_82_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25538_ net2468 _09024_ _09030_ _09017_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13552_ execute.io_mem_rd\[2\] execute.io_mem_rd\[3\] VGND VGND VPWR VPWR _09919_
+ sky130_fd_sc_hd__nor2_1
X_28257_ clknet_leaf_92_clock _01279_ VGND VGND VPWR VPWR csr._minstret_T_3\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16271_ decode.regfile.registers_0\[25\] _11539_ _12242_ VGND VGND VPWR VPWR _12243_
+ sky130_fd_sc_hd__o21bai_1
X_25469_ _10130_ VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__buf_2
XFILLER_0_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18010_ _12493_ decode.regfile.registers_29\[30\] _03375_ _03406_ _12702_ VGND VGND
+ VPWR VPWR _03407_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27208_ clknet_leaf_363_clock _00237_ VGND VGND VPWR VPWR decode.regfile.registers_28\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15222_ _11218_ VGND VGND VPWR VPWR _11219_ sky130_fd_sc_hd__clkbuf_4
X_28188_ clknet_leaf_112_clock _01210_ VGND VGND VPWR VPWR csr.io_mret_vector\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15153_ _10645_ decode.immGen._imm_T_24\[1\] decode.immGen._imm_T_24\[11\] VGND VGND
+ VPWR VPWR _11150_ sky130_fd_sc_hd__nand3b_4
X_27139_ clknet_leaf_358_clock _00168_ VGND VGND VPWR VPWR decode.regfile.registers_26\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14104_ _10097_ _10312_ VGND VGND VPWR VPWR _10319_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19961_ _10731_ _03599_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__nor2_1
X_15084_ _11079_ _10979_ _11080_ VGND VGND VPWR VPWR _11081_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14035_ net1730 _10271_ _10278_ _10275_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__o211a_1
X_18912_ _04208_ _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__nor2b_2
X_19892_ _05159_ _05158_ _03864_ _03862_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_224_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18843_ _04137_ _04141_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_8_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_220_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18774_ _03890_ decode.id_ex_imm_reg\[6\] _04072_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_220_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ decode.regfile.registers_14\[17\] _11360_ _11274_ decode.regfile.registers_15\[17\]
+ _11202_ VGND VGND VPWR VPWR _11966_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17725_ _03116_ _03127_ _12591_ _03128_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14937_ _10964_ _10665_ decode.immGen._imm_T_10\[0\] _10965_ VGND VGND VPWR VPWR
+ _10966_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_19_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17656_ _13081_ _13168_ decode.regfile.registers_23\[21\] _12995_ VGND VGND VPWR
+ VPWR _03062_ sky130_fd_sc_hd__or4_1
X_14868_ _10910_ VGND VGND VPWR VPWR _10911_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16607_ _12571_ VGND VGND VPWR VPWR _12572_ sky130_fd_sc_hd__clkbuf_4
X_13819_ _10151_ VGND VGND VPWR VPWR _10152_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17587_ _13099_ _13262_ _13182_ decode.regfile.registers_29\[19\] _02994_ VGND VGND
+ VPWR VPWR _02995_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14799_ _10730_ _10816_ _10822_ _10823_ _10841_ VGND VGND VPWR VPWR _10842_ sky130_fd_sc_hd__o311a_1
XFILLER_0_57_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19326_ _04442_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16538_ _12502_ VGND VGND VPWR VPWR _12503_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19257_ _04532_ _04545_ _04551_ _10576_ _10910_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_70_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16469_ _10652_ _11112_ _11118_ _12435_ VGND VGND VPWR VPWR _12436_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18208_ net214 _03527_ _03545_ _10999_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19188_ _04247_ _04355_ _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_147_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18139_ _03498_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21150_ _06068_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold146 io_fetch_data[4] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold157 io_fetch_data[14] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold168 fetch.bht.bhtTable_valid\[13\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
X_20101_ _00562_ _05228_ _05313_ _05231_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold179 fetch.btb.btbTable\[13\]\[0\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
X_21081_ _06027_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20032_ decode.id_ex_imm_reg\[5\] _10704_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24840_ _06117_ net1629 _08607_ VGND VGND VPWR VPWR _08608_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_14 _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24771_ _08571_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__clkbuf_1
X_21983_ net1834 _06588_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__or2_1
XINSDIODE1_25 _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_36 _08937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_250_clock clknet_5_19__leaf_clock VGND VGND VPWR VPWR clknet_leaf_250_clock
+ sky130_fd_sc_hd__clkbuf_8
XINSDIODE1_47 _09956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_58 _10091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26510_ net2183 _09592_ _09603_ _09595_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__o211a_1
X_23722_ net958 _10772_ _08003_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__mux2_1
X_20934_ _05937_ _05945_ net52 VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__and3_1
XINSDIODE1_69 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27490_ clknet_leaf_33_clock _00519_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26441_ net2285 _09561_ _09563_ _09553_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__o211a_1
X_23653_ net1753 csr.io_mem_pc\[18\] _07972_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__mux2_1
X_20865_ net119 _05903_ _05899_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29160_ clknet_leaf_213_clock _02173_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_22604_ csr._minstret_T_3\[49\] _07178_ _07179_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23584_ _06115_ net2030 _07930_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__mux2_1
X_26372_ net2596 _09518_ _09523_ _09512_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_265_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_265_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20796_ _05872_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28111_ clknet_leaf_80_clock _01133_ VGND VGND VPWR VPWR csr.minstret\[16\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_147_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22535_ _07097_ _07105_ _07118_ _07128_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__o2bb2a_1
X_25323_ _08892_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29091_ clknet_leaf_71_clock _02104_ VGND VGND VPWR VPWR csr._mcycle_T_3\[39\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_137_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28042_ clknet_leaf_53_clock _01064_ VGND VGND VPWR VPWR decode.control.io_opcode\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_49_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25254_ _08093_ net1635 _08848_ VGND VGND VPWR VPWR _08857_ sky130_fd_sc_hd__mux2_1
X_22466_ _06916_ _06977_ _07007_ _07060_ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__or4b_4
XFILLER_0_84_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24205_ _08099_ net1290 _06251_ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__mux2_1
X_21417_ _06223_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25185_ _08821_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__clkbuf_1
X_22397_ fetch.bht.bhtTable_tag\[8\]\[21\] fetch.bht.bhtTable_tag\[9\]\[21\] fetch.bht.bhtTable_tag\[10\]\[21\]
+ fetch.bht.bhtTable_tag\[11\]\[21\] _06707_ _06730_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24136_ _08241_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__clkbuf_1
X_21348_ net1055 csr.io_mem_pc\[31\] _06179_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28944_ clknet_leaf_106_clock _01957_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_24067_ net1031 execute.io_target_pc\[21\] _08198_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__mux2_1
Xhold680 fetch.bht.bhtTable_target_pc\[1\]\[24\] VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_203_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_203_clock
+ sky130_fd_sc_hd__clkbuf_8
X_21279_ net1302 _06145_ _06141_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold691 decode.regfile.registers_31\[3\] VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd3_1
X_23018_ net96 net227 _07427_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__and3_1
X_28875_ clknet_leaf_89_clock _01888_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15840_ decode.regfile.registers_23\[13\] _11087_ _11797_ _11823_ VGND VGND VPWR
+ VPWR _11824_ sky130_fd_sc_hd__o22a_1
X_27826_ clknet_leaf_317_clock _00855_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_9_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2070 decode.regfile.registers_9\[12\] VGND VGND VPWR VPWR net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2081 decode.regfile.registers_22\[30\] VGND VGND VPWR VPWR net2308 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_218_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_218_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold2092 decode.regfile.registers_23\[25\] VGND VGND VPWR VPWR net2319 sky130_fd_sc_hd__dlygate4sd3_1
X_15771_ _11756_ decode.regfile.registers_28\[11\] _11067_ _11681_ _11440_ VGND VGND
+ VPWR VPWR _11757_ sky130_fd_sc_hd__o2111a_1
X_27757_ clknet_leaf_325_clock _00786_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_24969_ _08692_ VGND VGND VPWR VPWR _08693_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_188_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17510_ decode.regfile.registers_2\[18\] _10616_ _12729_ VGND VGND VPWR VPWR _13457_
+ sky130_fd_sc_hd__o21ai_1
Xhold1380 decode.regfile.registers_10\[9\] VGND VGND VPWR VPWR net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1391 fetch.bht.bhtTable_target_pc\[12\]\[23\] VGND VGND VPWR VPWR net1618 sky130_fd_sc_hd__dlygate4sd3_1
X_14722_ csr.io_mem_pc\[16\] csr.io_mem_pc\[17\] csr.io_mem_pc\[18\] _10764_ VGND
+ VGND VPWR VPWR _10765_ sky130_fd_sc_hd__and4_1
X_26708_ _09385_ _09710_ VGND VGND VPWR VPWR _09718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18490_ _03781_ _03788_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__nor2_2
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27688_ clknet_leaf_21_clock _00717_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17441_ _13388_ _12726_ _13389_ VGND VGND VPWR VPWR _13390_ sky130_fd_sc_hd__a21oi_1
X_29427_ clknet_leaf_260_clock _02440_ VGND VGND VPWR VPWR decode.regfile.registers_5\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_14653_ _10694_ execute.io_target_pc\[12\] VGND VGND VPWR VPWR _10696_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26639_ _09392_ _09676_ VGND VGND VPWR VPWR _09678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13604_ _09939_ memory.io_wb_readdata\[2\] _09966_ VGND VGND VPWR VPWR _09967_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_200_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29358_ clknet_leaf_227_clock _02371_ VGND VGND VPWR VPWR decode.regfile.registers_3\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_17372_ decode.regfile.registers_12\[14\] _12745_ _13309_ _13322_ _12658_ VGND VGND
+ VPWR VPWR _13323_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14584_ decode.immGen._imm_T_24\[1\] VGND VGND VPWR VPWR _10627_ sky130_fd_sc_hd__buf_4
XFILLER_0_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19111_ _04225_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_188_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28309_ clknet_leaf_219_clock _01322_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16323_ decode.regfile.registers_16\[26\] _11124_ _12276_ _12293_ _11127_ VGND VGND
+ VPWR VPWR _12294_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13535_ _09910_ VGND VGND VPWR VPWR _09911_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_188_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29289_ clknet_leaf_242_clock _02302_ VGND VGND VPWR VPWR decode.regfile.registers_1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19042_ _04297_ _04261_ _04263_ _04340_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16254_ decode.regfile.registers_20\[24\] _11102_ _11327_ _12226_ VGND VGND VPWR
+ VPWR _12227_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15205_ _11201_ VGND VGND VPWR VPWR _11202_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16185_ decode.regfile.registers_19\[22\] _11453_ _11219_ _12159_ VGND VGND VPWR
+ VPWR _12160_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15136_ net320 _10624_ _11058_ VGND VGND VPWR VPWR _11133_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_226_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19944_ decode.id_ex_memread_reg VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__clkbuf_2
X_15067_ _11063_ VGND VGND VPWR VPWR _11064_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_222_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14018_ _10074_ _10268_ VGND VGND VPWR VPWR _10269_ sky130_fd_sc_hd__nand2_1
X_19875_ _03803_ _05123_ _05144_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18826_ _03817_ _04124_ _03774_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_223_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18757_ _04055_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__buf_2
XFILLER_0_175_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15969_ decode.regfile.registers_9\[17\] _11280_ _11134_ _11183_ VGND VGND VPWR VPWR
+ _11949_ sky130_fd_sc_hd__a31o_1
XFILLER_0_222_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17708_ decode.regfile.registers_18\[23\] _10925_ _12569_ _11023_ _11008_ VGND VGND
+ VPWR VPWR _03112_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_37_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18688_ decode.id_ex_imm_reg\[0\] _03726_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_177_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17639_ decode.regfile.registers_8\[21\] _12892_ _12603_ VGND VGND VPWR VPWR _03045_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20650_ _05780_ _05671_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19309_ _04417_ _04431_ _04272_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20581_ csr._minstret_T_3\[51\] _05577_ _05578_ _05721_ VGND VGND VPWR VPWR _05722_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22320_ _06907_ _06913_ net227 VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22251_ fetch.bht.bhtTable_tag\[14\]\[19\] fetch.bht.bhtTable_tag\[15\]\[19\] _06809_
+ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21202_ _06096_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22182_ _06774_ _06661_ _06633_ _06776_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_83_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21133_ _06059_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26990_ net905 _09840_ _09878_ _06396_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25941_ _08939_ _09253_ VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__nand2_1
X_21064_ _06018_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20015_ _05238_ _05239_ _00550_ _05227_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__o22a_1
X_28660_ clknet_leaf_119_clock _01673_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25872_ net2237 _09213_ _09221_ _09222_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_213_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27611_ clknet_leaf_158_clock _00640_ VGND VGND VPWR VPWR execute.io_target_pc\[20\]
+ sky130_fd_sc_hd__dfxtp_4
X_24823_ _06101_ net1267 _08422_ VGND VGND VPWR VPWR _08599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28591_ clknet_leaf_107_clock _01604_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27542_ clknet_leaf_45_clock _00571_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24754_ _08561_ VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__buf_6
X_21966_ csr.mscratch\[8\] _06574_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23705_ _07991_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__buf_4
X_27473_ clknet_leaf_53_clock _00502_ VGND VGND VPWR VPWR csr.io_csr_address\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20917_ _05937_ _05933_ net43 VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__and3_1
X_24685_ net1441 execute.io_target_pc\[31\] _07285_ VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__mux2_1
X_21897_ net2798 _06521_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29212_ clknet_leaf_128_clock _02225_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26424_ _09404_ _09545_ VGND VGND VPWR VPWR _09554_ sky130_fd_sc_hd__nand2_1
X_23636_ net765 _10878_ _07961_ VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__mux2_1
X_20848_ net110 _05891_ _05899_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29143_ clknet_leaf_92_clock _02156_ VGND VGND VPWR VPWR csr.mcycle\[27\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_182_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26355_ _09410_ _09502_ VGND VGND VPWR VPWR _09514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23567_ net2772 _07918_ decode.id_ex_memread_reg VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__or3b_1
XFILLER_0_119_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20779_ net133 execute.io_mem_zero net134 VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_25_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25306_ _03580_ net442 VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22518_ _07111_ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__buf_4
X_29074_ clknet_leaf_197_clock _02087_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_23498_ net2777 _07875_ _07888_ _07879_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__o211a_1
X_26286_ net1608 _09462_ _09474_ _09471_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28025_ clknet_leaf_200_clock _01047_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25237_ _09905_ VGND VGND VPWR VPWR _08848_ sky130_fd_sc_hd__clkbuf_8
X_22449_ _07042_ _07043_ _06635_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25168_ _08812_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_142_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_142_clock
+ sky130_fd_sc_hd__clkbuf_8
X_24119_ net1379 execute.io_target_pc\[14\] _08232_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25099_ _08777_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17990_ decode.regfile.registers_8\[30\] _12843_ _12605_ VGND VGND VPWR VPWR _03387_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28927_ clknet_leaf_180_clock _01940_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16941_ decode.regfile.registers_16\[4\] _12674_ _12901_ VGND VGND VPWR VPWR _12902_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_208_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19660_ _04935_ _04912_ _04936_ _04192_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__o211ai_1
X_28858_ clknet_leaf_128_clock _01871_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_157_clock clknet_5_24__leaf_clock VGND VGND VPWR VPWR clknet_leaf_157_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16872_ _12833_ VGND VGND VPWR VPWR _12834_ sky130_fd_sc_hd__buf_2
XFILLER_0_216_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18611_ _03817_ _03905_ _03774_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__a21oi_2
X_15823_ decode.regfile.registers_2\[13\] _11295_ _11151_ _11806_ VGND VGND VPWR VPWR
+ _11807_ sky130_fd_sc_hd__o211a_1
X_27809_ clknet_leaf_326_clock _00838_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_19591_ _04349_ _04358_ _04370_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28789_ clknet_leaf_116_clock _01802_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18542_ execute.io_reg_pc\[24\] _03777_ _03666_ net116 _03840_ VGND VGND VPWR VPWR
+ _03841_ sky130_fd_sc_hd__o221a_1
X_15754_ _11382_ decode.regfile.registers_10\[11\] _11315_ _11739_ VGND VGND VPWR
+ VPWR _11740_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14705_ _10747_ VGND VGND VPWR VPWR _10748_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18473_ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__clkbuf_8
X_15685_ decode.regfile.registers_23\[9\] _11262_ _11089_ _11493_ _11672_ VGND VGND
+ VPWR VPWR _11673_ sky130_fd_sc_hd__o221a_1
XFILLER_0_158_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17424_ _13215_ decode.regfile.registers_28\[15\] _13093_ VGND VGND VPWR VPWR _13374_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14636_ execute.io_target_pc\[6\] _10678_ VGND VGND VPWR VPWR _10679_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_215_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_215_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17355_ decode.regfile.registers_18\[14\] _12570_ _12560_ VGND VGND VPWR VPWR _13306_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14567_ _10609_ VGND VGND VPWR VPWR _10610_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16306_ decode.regfile.registers_10\[26\] _11184_ _11181_ VGND VGND VPWR VPWR _12277_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13518_ _09896_ VGND VGND VPWR VPWR _09897_ sky130_fd_sc_hd__clkbuf_8
X_17286_ decode.regfile.registers_13\[12\] _12659_ _13224_ _13238_ _12984_ VGND VGND
+ VPWR VPWR _13239_ sky130_fd_sc_hd__o221a_1
X_14498_ _10142_ _10505_ VGND VGND VPWR VPWR _10545_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19025_ _04264_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16237_ _10660_ _10655_ net346 decode.regfile.registers_2\[24\] _11296_ VGND VGND
+ VPWR VPWR _12210_ sky130_fd_sc_hd__o32a_1
XFILLER_0_113_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16168_ _11313_ decode.regfile.registers_4\[22\] _10647_ _10629_ _11462_ VGND VGND
+ VPWR VPWR _12143_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_3_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15119_ _11115_ VGND VGND VPWR VPWR _11116_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16099_ _12018_ _12056_ _12073_ _12075_ VGND VGND VPWR VPWR _12076_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19927_ _04225_ _03766_ _04424_ _03705_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__or4b_1
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19858_ _03801_ _03802_ _05126_ _03830_ _04219_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18809_ _10039_ _10040_ memory.csr_read_data_out_reg\[12\] _09942_ VGND VGND VPWR
+ VPWR _04108_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_69_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19789_ _04325_ _05006_ _04317_ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_69_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21820_ _06479_ net1158 _06396_ _06483_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21751_ net985 _10807_ _06428_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20702_ _05818_ decode.id_ex_rs1_data_reg\[11\] _05670_ VGND VGND VPWR VPWR _05819_
+ sky130_fd_sc_hd__a21oi_1
X_24470_ _08097_ net1967 _08411_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__mux2_1
X_21682_ csr._mcycle_T_2\[23\] _06321_ _06387_ csr.minstret\[23\] VGND VGND VPWR VPWR
+ _06388_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_176_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20633_ csr._minstret_T_3\[59\] _05616_ _05618_ csr._csr_read_data_T_8\[27\] _05765_
+ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23421_ execute.io_target_pc\[31\] _07091_ _07831_ _07842_ _06032_ VGND VGND VPWR
+ VPWR _07843_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_134_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23352_ fetch.bht.bhtTable_target_pc\[4\]\[27\] fetch.bht.bhtTable_target_pc\[5\]\[27\]
+ fetch.bht.bhtTable_target_pc\[6\]\[27\] fetch.bht.bhtTable_target_pc\[7\]\[27\]
+ _07555_ _07710_ VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_199_Left_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26140_ _09377_ _09374_ VGND VGND VPWR VPWR _09378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20564_ csr.minstret\[17\] _05574_ _05586_ csr.mcycle\[17\] _05706_ VGND VGND VPWR
+ VPWR _05707_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_24_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22303_ _06894_ _06895_ _06896_ _06897_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23283_ _07709_ _07711_ _07712_ _07713_ _07122_ _07084_ VGND VGND VPWR VPWR _07714_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26071_ net2194 _09329_ _09337_ _09333_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__o211a_1
X_20495_ csr._csr_read_data_T_8\[8\] _05591_ _05516_ _05528_ _05646_ VGND VGND VPWR
+ VPWR _05647_ sky130_fd_sc_hd__a41o_1
XFILLER_0_132_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22234_ _06828_ _06678_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__or2b_1
X_25022_ _08728_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29830_ clknet_leaf_297_clock _02843_ VGND VGND VPWR VPWR decode.regfile.registers_18\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_22165_ _06673_ _06755_ _06757_ _06759_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_74_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_74_clock
+ sky130_fd_sc_hd__clkbuf_8
X_21116_ _05857_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__clkbuf_2
X_29761_ clknet_leaf_310_clock _02774_ VGND VGND VPWR VPWR decode.regfile.registers_16\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_22096_ net302 VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__clkbuf_8
X_26973_ _10101_ _09862_ VGND VGND VPWR VPWR _09870_ sky130_fd_sc_hd__nand2_1
Xfanout220 net84 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_4
XFILLER_0_227_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28712_ clknet_leaf_99_clock _01725_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25924_ net1690 _09242_ _09252_ _09250_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__o211a_1
X_21047_ execute.csr_read_data_out_reg\[13\] _06002_ _05998_ VGND VGND VPWR VPWR _06009_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_121_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29692_ clknet_leaf_290_clock _02705_ VGND VGND VPWR VPWR decode.regfile.registers_14\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28643_ clknet_leaf_132_clock _01656_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25855_ _09198_ VGND VGND VPWR VPWR _09213_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_213_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_89_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_89_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24806_ _08099_ net1354 _08585_ VGND VGND VPWR VPWR _08590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28574_ clknet_leaf_186_clock _01587_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25786_ net2209 _09170_ _09173_ _09169_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__o211a_1
X_22998_ _07444_ _07406_ _07085_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__a21oi_1
X_27525_ clknet_leaf_44_clock _00554_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfxtp_2
X_24737_ _08099_ net1217 _06283_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21949_ net559 _06572_ _06575_ _10546_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__o211a_1
XINSDIODE1_109 _10935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_12_clock
+ sky130_fd_sc_hd__clkbuf_8
X_27456_ clknet_leaf_137_clock _00485_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15470_ _11313_ decode.regfile.registers_4\[4\] _11191_ _10630_ _11462_ VGND VGND
+ VPWR VPWR _11463_ sky130_fd_sc_hd__a2111o_1
X_24668_ _08517_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26407_ _09387_ _09535_ VGND VGND VPWR VPWR _09544_ sky130_fd_sc_hd__nand2_1
X_14421_ _10136_ _10462_ VGND VGND VPWR VPWR _10501_ sky130_fd_sc_hd__nand2_1
X_23619_ _06149_ net1700 _07952_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27387_ clknet_leaf_15_clock _00416_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24599_ net1089 execute.io_target_pc\[21\] _08473_ VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29126_ clknet_leaf_76_clock _02139_ VGND VGND VPWR VPWR csr.mcycle\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17140_ _12708_ net435 _13056_ _13096_ _12705_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__o221a_1
X_26338_ net712 _09491_ _09504_ _09499_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__o211a_1
X_14352_ _10373_ _10195_ _09932_ _10149_ VGND VGND VPWR VPWR _10461_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_210_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_27_clock
+ sky130_fd_sc_hd__clkbuf_8
X_29057_ clknet_leaf_170_clock _02070_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_17071_ _13012_ _13027_ _13028_ VGND VGND VPWR VPWR _13029_ sky130_fd_sc_hd__o21ai_1
X_26269_ _09400_ _09459_ VGND VGND VPWR VPWR _09465_ sky130_fd_sc_hd__nand2_1
X_14283_ net2187 _10419_ _10422_ _10411_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28008_ clknet_leaf_190_clock _01030_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_16022_ decode.regfile.registers_12\[18\] _10639_ _11690_ _11198_ _12000_ VGND VGND
+ VPWR VPWR _12001_ sky130_fd_sc_hd__o311a_1
XFILLER_0_126_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_208_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_208_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17973_ _10929_ decode.regfile.registers_28\[29\] _12697_ VGND VGND VPWR VPWR _03371_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_209_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16924_ decode.regfile.registers_2\[4\] _12835_ _12836_ _12884_ VGND VGND VPWR VPWR
+ _12885_ sky130_fd_sc_hd__a211o_1
X_19712_ _04546_ _04428_ _04792_ _04988_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_204_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19643_ net309 _04290_ _04301_ _04707_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__or4b_1
X_16855_ _12701_ decode.regfile.registers_28\[2\] _12698_ VGND VGND VPWR VPWR _12818_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_205_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15806_ decode.regfile.registers_25\[12\] _11483_ _11484_ decode.regfile.registers_24\[12\]
+ VGND VGND VPWR VPWR _11791_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19574_ _04295_ _04293_ _04779_ _04856_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__o31a_2
XFILLER_0_220_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_196_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16786_ _12650_ _12723_ _12669_ decode.regfile.registers_14\[1\] _12749_ VGND VGND
+ VPWR VPWR _12750_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_217_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13998_ net452 _10243_ _10257_ _10249_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18525_ decode.id_ex_rs2_data_reg\[27\] _03747_ _03822_ _03823_ VGND VGND VPWR VPWR
+ _03824_ sky130_fd_sc_hd__o211a_1
X_15737_ _10981_ VGND VGND VPWR VPWR _11723_ sky130_fd_sc_hd__buf_2
XFILLER_0_133_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18456_ _03719_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__buf_6
XFILLER_0_213_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15668_ _10659_ _10654_ _11150_ decode.regfile.registers_3\[9\] VGND VGND VPWR VPWR
+ _11656_ sky130_fd_sc_hd__or4b_1
XFILLER_0_146_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17407_ _12666_ _12773_ _12984_ decode.regfile.registers_14\[15\] _13356_ VGND VGND
+ VPWR VPWR _13357_ sky130_fd_sc_hd__o221a_1
X_14619_ _10660_ VGND VGND VPWR VPWR _10662_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_173_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18387_ _03675_ _03685_ _03655_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__o21ai_4
X_15599_ decode.regfile.registers_11\[7\] _11070_ _11470_ _11278_ VGND VGND VPWR VPWR
+ _11589_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17338_ decode.regfile.registers_22\[13\] _12528_ _13288_ _13289_ VGND VGND VPWR
+ VPWR _13290_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17269_ decode.regfile.registers_20\[12\] _11024_ _12553_ _12823_ _12824_ VGND VGND
+ VPWR VPWR _13222_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_12_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19008_ _04274_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_168_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20280_ decode.id_ex_pc_reg\[14\] _05458_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_1__f_clock clknet_2_0_0_clock VGND VGND VPWR VPWR clknet_5_1__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_90_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23970_ net1282 execute.io_target_pc\[6\] _08153_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__mux2_1
Xhold1902 decode.io_id_pc\[14\] VGND VGND VPWR VPWR net2129 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1913 csr._minstret_T_3\[58\] VGND VGND VPWR VPWR net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1924 fetch.bht.bhtTable_target_pc\[10\]\[14\] VGND VGND VPWR VPWR net2151 sky130_fd_sc_hd__dlygate4sd3_1
X_22921_ _07369_ _07370_ _07371_ VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__mux2_1
Xhold1935 decode.regfile.registers_2\[0\] VGND VGND VPWR VPWR net2162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1946 decode.regfile.registers_4\[17\] VGND VGND VPWR VPWR net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1957 decode.io_id_pc\[15\] VGND VGND VPWR VPWR net2184 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_123_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1968 decode.io_id_pc\[5\] VGND VGND VPWR VPWR net2195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1979 decode.regfile.registers_8\[2\] VGND VGND VPWR VPWR net2206 sky130_fd_sc_hd__dlygate4sd3_1
X_25640_ _08939_ _09079_ VGND VGND VPWR VPWR _09089_ sky130_fd_sc_hd__nand2_1
X_22852_ net1019 _10871_ _09898_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21803_ _06457_ _06466_ _06470_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__and3b_1
X_25571_ _09023_ VGND VGND VPWR VPWR _09049_ sky130_fd_sc_hd__buf_2
XFILLER_0_195_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22783_ _07285_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27310_ clknet_leaf_9_clock _00339_ VGND VGND VPWR VPWR decode.regfile.registers_31\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24522_ _08442_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__clkbuf_1
X_28290_ clknet_leaf_85_clock _01312_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_21734_ _06429_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27241_ clknet_leaf_0_clock _00270_ VGND VGND VPWR VPWR decode.regfile.registers_29\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24453_ _08081_ net2265 _08400_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__mux2_1
X_21665_ _06374_ _06372_ _06327_ _06375_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_35_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1090 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23404_ _07064_ _07819_ _07820_ _07826_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20616_ _05627_ csr.io_mret_vector\[24\] _05603_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__o21a_1
X_27172_ clknet_leaf_362_clock _00201_ VGND VGND VPWR VPWR decode.regfile.registers_27\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_24384_ _08369_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21596_ csr.minstret\[0\] net578 csr.io_inst_retired _06318_ _06324_ VGND VGND VPWR
+ VPWR _01117_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_46_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26123_ net2346 _09356_ _09366_ _09359_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__o211a_1
X_23335_ fetch.bht.bhtTable_target_pc\[8\]\[26\] fetch.bht.bhtTable_target_pc\[9\]\[26\]
+ fetch.bht.bhtTable_target_pc\[10\]\[26\] fetch.bht.bhtTable_target_pc\[11\]\[26\]
+ _07068_ _07656_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__mux4_1
X_20547_ _05691_ _05572_ _05561_ csr.mcycle\[15\] VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26054_ net2714 _09287_ _09326_ _09318_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__o211a_1
X_23266_ fetch.bht.bhtTable_target_pc\[12\]\[21\] fetch.bht.bhtTable_target_pc\[13\]\[21\]
+ fetch.bht.bhtTable_target_pc\[14\]\[21\] fetch.bht.bhtTable_target_pc\[15\]\[21\]
+ _07098_ _07113_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__mux4_1
X_20478_ csr._minstret_T_3\[38\] _05616_ _05622_ csr._csr_read_data_T_8\[6\] _05631_
+ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25005_ csr.mcycle\[4\] csr.mcycle\[3\] csr.mcycle\[5\] _03557_ csr.mcycle\[6\] VGND
+ VGND VPWR VPWR _08717_ sky130_fd_sc_hd__a41o_1
XFILLER_0_30_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22217_ _06707_ fetch.bht.bhtTable_tag\[11\]\[20\] _06649_ VGND VGND VPWR VPWR _06812_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23197_ _07619_ _07573_ _07620_ _07632_ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_56_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22148_ fetch.bht.bhtTable_tag\[6\]\[23\] fetch.bht.bhtTable_tag\[7\]\[23\] _06646_
+ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__mux2_1
X_29813_ clknet_leaf_296_clock _02826_ VGND VGND VPWR VPWR decode.regfile.registers_17\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22079_ _06643_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__buf_6
X_14970_ decode.immGen._imm_T_10\[4\] _10667_ _10975_ _10994_ VGND VGND VPWR VPWR
+ _10995_ sky130_fd_sc_hd__a22o_1
X_29744_ clknet_leaf_284_clock _02757_ VGND VGND VPWR VPWR decode.regfile.registers_15\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_26956_ net586 _09849_ VGND VGND VPWR VPWR _09860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13921_ net491 _10199_ _10212_ _10206_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__o211a_1
X_25907_ _09241_ VGND VGND VPWR VPWR _09243_ sky130_fd_sc_hd__buf_2
X_29675_ clknet_leaf_278_clock _02688_ VGND VGND VPWR VPWR decode.regfile.registers_13\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26887_ net1514 _09809_ _09820_ _09812_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__o211a_1
X_28626_ clknet_leaf_107_clock _01639_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16640_ _12592_ _12531_ _10592_ VGND VGND VPWR VPWR _12605_ sky130_fd_sc_hd__and3_2
X_13852_ net1970 _10167_ _10171_ _10162_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__o211a_1
X_25838_ net2422 _09199_ _09203_ _09194_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28557_ clknet_leaf_235_clock _01570_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16571_ _12524_ _12523_ _12535_ VGND VGND VPWR VPWR _12536_ sky130_fd_sc_hd__and3_1
X_13783_ memory.csr_read_data_out_reg\[27\] _09987_ _10120_ VGND VGND VPWR VPWR _10121_
+ sky130_fd_sc_hd__o21ai_4
X_25769_ net2650 _09156_ _09163_ _09153_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18310_ _03620_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15522_ decode.regfile.registers_16\[5\] _11122_ _11496_ _11513_ VGND VGND VPWR VPWR
+ _11514_ sky130_fd_sc_hd__o22a_1
X_27508_ clknet_leaf_15_clock _00537_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19290_ _04226_ _04582_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_191_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28488_ clknet_leaf_206_clock _01501_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18241_ csr._mcycle_T_3\[37\] csr._mcycle_T_3\[36\] csr._mcycle_T_3\[35\] csr._mcycle_T_3\[34\]
+ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__or4_1
XFILLER_0_155_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27439_ clknet_leaf_146_clock _00468_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_15453_ _10959_ VGND VGND VPWR VPWR _11446_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_194_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14404_ _10092_ _10487_ VGND VGND VPWR VPWR _10492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18172_ _03463_ _03464_ _03465_ decode.control.io_funct7\[5\] VGND VGND VPWR VPWR
+ _03514_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_26_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15384_ decode.regfile.registers_7\[2\] _11378_ _11170_ decode.regfile.registers_6\[2\]
+ _11281_ VGND VGND VPWR VPWR _11379_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17123_ decode.regfile.registers_22\[8\] _12527_ _13078_ _13079_ _12686_ VGND VGND
+ VPWR VPWR _13080_ sky130_fd_sc_hd__a221o_1
X_29109_ clknet_leaf_16_clock _02122_ VGND VGND VPWR VPWR csr._mcycle_T_3\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14335_ _10107_ _10444_ VGND VGND VPWR VPWR _10452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap206 _03724_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_8
Xhold509 _01186_ VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap217 _06313_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
X_17054_ decode.regfile.registers_12\[7\] _12745_ _12587_ _12533_ VGND VGND VPWR VPWR
+ _13012_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_64_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14266_ _10122_ _10400_ VGND VGND VPWR VPWR _10412_ sky130_fd_sc_hd__nand2_1
X_16005_ _11446_ decode.regfile.registers_26\[18\] _11447_ _11348_ _10993_ VGND VGND
+ VPWR VPWR _11984_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_21_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14197_ net487 _10333_ _10371_ _10369_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_206_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17956_ _03340_ _03352_ _12591_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__o211ai_1
Xhold1209 fetch.bht.bhtTable_target_pc\[4\]\[17\] VGND VGND VPWR VPWR net1436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16907_ _12701_ decode.regfile.registers_28\[3\] _12698_ VGND VGND VPWR VPWR _12869_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17887_ decode.regfile.registers_19\[27\] _12678_ _03264_ _03286_ _12544_ VGND VGND
+ VPWR VPWR _03287_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_1202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19626_ _04512_ _04905_ _04883_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_206_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16838_ decode.regfile.registers_17\[2\] _12580_ _12566_ VGND VGND VPWR VPWR _12801_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16769_ decode.regfile.registers_2\[1\] _12633_ _12627_ decode.regfile.registers_3\[1\]
+ _12732_ VGND VGND VPWR VPWR _12733_ sky130_fd_sc_hd__o221a_1
X_19557_ _04637_ _04170_ _04835_ _04839_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_88_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18508_ net239 _03797_ net196 VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_157_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19488_ _04570_ _04567_ _04371_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18439_ _03737_ decode.io_wb_rd\[1\] VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21450_ _06240_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20401_ csr.io_csr_address\[11\] net218 _05520_ _05524_ VGND VGND VPWR VPWR _05561_
+ sky130_fd_sc_hd__and4_2
X_21381_ _06203_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23120_ fetch.bht.bhtTable_target_pc\[4\]\[13\] fetch.bht.bhtTable_target_pc\[5\]\[13\]
+ fetch.bht.bhtTable_target_pc\[6\]\[13\] fetch.bht.bhtTable_target_pc\[7\]\[13\]
+ _07099_ _07101_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__mux4_1
XFILLER_0_189_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20332_ _05499_ _05500_ _05416_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23051_ _07406_ _07492_ _07494_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_187_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20263_ _10706_ _05440_ decode.id_ex_pc_reg\[10\] VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__a21oi_1
X_22002_ csr.mscratch\[23\] _06601_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20194_ decode.id_ex_imm_reg\[28\] decode.id_ex_pc_reg\[28\] VGND VGND VPWR VPWR
+ _05393_ sky130_fd_sc_hd__and2_1
Xhold2400 decode.regfile.registers_9\[24\] VGND VGND VPWR VPWR net2627 sky130_fd_sc_hd__dlygate4sd3_1
X_26810_ _09751_ VGND VGND VPWR VPWR _09776_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_51_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2411 csr._mcycle_T_3\[53\] VGND VGND VPWR VPWR net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2422 _01135_ VGND VGND VPWR VPWR net2649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27790_ clknet_leaf_322_clock _00819_ VGND VGND VPWR VPWR memory.io_wb_readdata\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2433 decode.regfile.registers_22\[20\] VGND VGND VPWR VPWR net2660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2444 decode.regfile.registers_11\[20\] VGND VGND VPWR VPWR net2671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1710 _01231_ VGND VGND VPWR VPWR net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2455 decode.regfile.registers_18\[29\] VGND VGND VPWR VPWR net2682 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2466 decode.regfile.registers_0\[26\] VGND VGND VPWR VPWR net2693 sky130_fd_sc_hd__dlygate4sd3_1
X_26741_ _09420_ _09733_ VGND VGND VPWR VPWR _09737_ sky130_fd_sc_hd__nand2_1
Xhold1721 decode.regfile.registers_5\[21\] VGND VGND VPWR VPWR net1948 sky130_fd_sc_hd__dlygate4sd3_1
X_23953_ net1201 _08111_ _06156_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__mux2_1
Xhold1732 fetch.bht.bhtTable_tag\[15\]\[9\] VGND VGND VPWR VPWR net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2477 csr.minstret\[3\] VGND VGND VPWR VPWR net2704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1743 decode.regfile.registers_23\[13\] VGND VGND VPWR VPWR net1970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2488 execute.io_mem_rd\[2\] VGND VGND VPWR VPWR net2715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2499 decode.regfile.registers_0\[15\] VGND VGND VPWR VPWR net2726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1754 decode.regfile.registers_3\[14\] VGND VGND VPWR VPWR net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1765 fetch.bht.bhtTable_target_pc\[7\]\[22\] VGND VGND VPWR VPWR net1992 sky130_fd_sc_hd__dlygate4sd3_1
X_22904_ net69 _06794_ _06806_ net90 VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_4_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29460_ clknet_leaf_261_clock _02473_ VGND VGND VPWR VPWR decode.regfile.registers_6\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26672_ net1915 _09692_ _09696_ _09688_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__o211a_1
Xhold1776 decode.regfile.registers_5\[24\] VGND VGND VPWR VPWR net2003 sky130_fd_sc_hd__dlygate4sd3_1
X_23884_ _08110_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__clkbuf_1
Xhold1787 csr.mscratch\[26\] VGND VGND VPWR VPWR net2014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1798 fetch.bht.bhtTable_tag\[6\]\[14\] VGND VGND VPWR VPWR net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28411_ clknet_leaf_142_clock _01424_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_4
X_25623_ _09067_ VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22835_ _07313_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__clkbuf_1
X_29391_ clknet_leaf_259_clock _02404_ VGND VGND VPWR VPWR decode.regfile.registers_4\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28342_ clknet_leaf_210_clock _01355_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25554_ _08929_ _09036_ VGND VGND VPWR VPWR _09040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22766_ _09901_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24505_ _08433_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21717_ net2679 _06415_ _06416_ _06352_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__a211oi_1
X_28273_ clknet_leaf_61_clock _01295_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_25485_ net2072 _08995_ _08999_ _08991_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22697_ csr._csr_read_data_T_8\[22\] _07235_ _07237_ _07234_ VGND VGND VPWR VPWR
+ _01306_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27224_ clknet_leaf_6_clock _00253_ VGND VGND VPWR VPWR decode.regfile.registers_29\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_24436_ _08064_ net2005 _08389_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21648_ _06317_ _06361_ _06362_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27155_ clknet_leaf_354_clock _00184_ VGND VGND VPWR VPWR decode.regfile.registers_27\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_24367_ _08360_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__clkbuf_1
X_21579_ _06310_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_80 _11892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 decode.regfile.registers_11\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26106_ net1154 _09356_ _09357_ _09346_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__o211a_1
X_14120_ _10142_ _10286_ VGND VGND VPWR VPWR _10327_ sky130_fd_sc_hd__nand2_1
X_23318_ csr._csr_read_data_T_8\[25\] _06480_ csr.io_mret_vector\[25\] _07621_ VGND
+ VGND VPWR VPWR _07746_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27086_ clknet_leaf_330_clock _00115_ VGND VGND VPWR VPWR decode.regfile.registers_24\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_24298_ _08060_ net1662 _08323_ VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14051_ _10286_ VGND VGND VPWR VPWR _10288_ sky130_fd_sc_hd__buf_2
X_26037_ _09263_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__buf_4
X_23249_ _07678_ _07679_ _07680_ _07681_ _07081_ _06740_ VGND VGND VPWR VPWR _07682_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17810_ _03187_ _03211_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18790_ net106 _03664_ _04088_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_201_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27988_ clknet_leaf_166_clock _01010_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _12967_ _03142_ _03143_ _03144_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__a31o_1
X_14953_ _10980_ VGND VGND VPWR VPWR _10981_ sky130_fd_sc_hd__clkbuf_8
X_26939_ net1543 _09839_ _09850_ _09836_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__o211a_1
X_29727_ clknet_leaf_311_clock _02740_ VGND VGND VPWR VPWR decode.regfile.registers_15\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13904_ _09970_ _10200_ VGND VGND VPWR VPWR _10203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17672_ decode.regfile.registers_15\[22\] _10611_ _10923_ _12876_ _12672_ VGND VGND
+ VPWR VPWR _03077_ sky130_fd_sc_hd__a41o_1
X_14884_ _10912_ _10913_ _10921_ decode.immGen._imm_T_10\[4\] VGND VGND VPWR VPWR
+ _10922_ sky130_fd_sc_hd__and4bb_1
X_29658_ clknet_leaf_288_clock _02671_ VGND VGND VPWR VPWR decode.regfile.registers_13\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_193_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19411_ _04273_ _04410_ _04290_ _04412_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__o211a_1
X_16623_ _12587_ VGND VGND VPWR VPWR _12588_ sky130_fd_sc_hd__clkbuf_4
X_28609_ clknet_leaf_174_clock _01622_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13835_ _10131_ VGND VGND VPWR VPWR _10162_ sky130_fd_sc_hd__clkbuf_4
X_29589_ clknet_leaf_274_clock _02602_ VGND VGND VPWR VPWR decode.regfile.registers_10\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19342_ _04443_ _04362_ _04633_ _04628_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__or4_1
X_16554_ _12518_ VGND VGND VPWR VPWR _12519_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13766_ _10106_ VGND VGND VPWR VPWR _10107_ sky130_fd_sc_hd__buf_6
XFILLER_0_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15505_ decode.regfile.registers_7\[5\] _11465_ _11466_ decode.regfile.registers_6\[5\]
+ _11281_ VGND VGND VPWR VPWR _11497_ sky130_fd_sc_hd__a221o_1
XFILLER_0_210_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19273_ _04356_ _04382_ _04541_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16485_ _11346_ net2331 _11038_ _10981_ _10994_ VGND VGND VPWR VPWR _12451_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_85_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13697_ _10048_ _10016_ VGND VGND VPWR VPWR _10049_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_152_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18224_ csr.mcycle\[6\] csr.mcycle\[8\] csr.mcycle\[7\] _03558_ VGND VGND VPWR VPWR
+ _03559_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15436_ decode.regfile.registers_20\[3\] _11103_ _11222_ _11429_ VGND VGND VPWR VPWR
+ _11430_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_152_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18155_ _11251_ _10577_ _10673_ _10911_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__nor4_1
XFILLER_0_182_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15367_ decode.regfile.registers_14\[2\] _11360_ _11274_ decode.regfile.registers_15\[2\]
+ _11361_ VGND VGND VPWR VPWR _11362_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17106_ _13060_ _13061_ _13062_ VGND VGND VPWR VPWR _13063_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14318_ net517 _10434_ _10442_ _10440_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18086_ _03468_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__clkbuf_1
X_15298_ decode.regfile.registers_3\[1\] _11292_ _11293_ _10635_ VGND VGND VPWR VPWR
+ _11294_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold306 decode.regfile.registers_14\[9\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold317 decode.regfile.registers_20\[9\] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold328 decode.regfile.registers_14\[2\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ _11014_ _10936_ decode.regfile.registers_23\[6\] _12995_ VGND VGND VPWR VPWR
+ _12996_ sky130_fd_sc_hd__or4_1
Xhold339 decode.regfile.registers_29\[3\] VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_229_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14249_ net1528 _10390_ _10402_ _10398_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_229_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_182_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18988_ _04251_ _04252_ _04285_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1006 decode.regfile.registers_28\[13\] VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 fetch.bht.bhtTable_target_pc\[12\]\[3\] VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1028 fetch.bht.bhtTable_target_pc\[9\]\[28\] VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_183_Right_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17939_ _10926_ decode.regfile.registers_22\[29\] _12554_ _11009_ _12546_ VGND VGND
+ VPWR VPWR _03337_ sky130_fd_sc_hd__o2111a_1
Xhold1039 _10690_ VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20950_ _05956_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19609_ _04888_ _04452_ _04889_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__or3b_1
XFILLER_0_89_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20881_ _05858_ _09956_ net56 VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__and3_1
XFILLER_0_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22620_ _06377_ _07188_ _07190_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_81_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22551_ csr._minstret_T_3\[34\] _07139_ _07141_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_118_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_270 _08937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_281 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21502_ _06268_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__clkbuf_1
X_25270_ _08109_ net1522 _09906_ VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__mux2_1
XINSDIODE1_292 _12504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22482_ _07073_ _07074_ _07076_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24221_ _08049_ net1278 _06241_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21433_ _06124_ net2202 _06230_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24152_ _08249_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__clkbuf_1
X_21364_ _06194_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23103_ _07101_ _07543_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__and2b_1
X_20315_ _05358_ _05362_ decode.id_ex_rdsel_reg _05486_ _05487_ VGND VGND VPWR VPWR
+ _05488_ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24083_ net1078 execute.io_target_pc\[29\] _07991_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__mux2_1
X_21295_ _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__buf_4
X_28960_ clknet_leaf_161_clock _01973_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold840 fetch.bht.bhtTable_tag\[4\]\[1\] VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold851 fetch.bht.bhtTable_target_pc\[3\]\[29\] VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold862 fetch.bht.bhtTable_target_pc\[11\]\[21\] VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23034_ _07476_ _07477_ _07112_ _07478_ _07082_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__o221a_1
Xhold873 fetch.bht.bhtTable_target_pc\[12\]\[17\] VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__dlygate4sd3_1
X_20246_ _05433_ _05434_ _05415_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__o21a_1
X_27911_ clknet_leaf_23_clock _00940_ VGND VGND VPWR VPWR csr.io_csr_write_address\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold884 fetch.bht.bhtTable_target_pc\[15\]\[1\] VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__dlygate4sd3_1
X_28891_ clknet_leaf_173_clock _01904_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold895 fetch.bht.bhtTable_target_pc\[1\]\[2\] VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27842_ clknet_leaf_326_clock _00871_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_20177_ _05068_ _05247_ _05378_ _05267_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_228_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2230 decode.regfile.registers_21\[23\] VGND VGND VPWR VPWR net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2241 decode.regfile.registers_3\[3\] VGND VGND VPWR VPWR net2468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2252 decode.regfile.registers_30\[1\] VGND VGND VPWR VPWR net2479 sky130_fd_sc_hd__dlygate4sd3_1
X_27773_ clknet_leaf_326_clock _00802_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24985_ net559 net569 _08701_ _08702_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__o31a_1
Xhold2263 decode.regfile.registers_22\[2\] VGND VGND VPWR VPWR net2490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2274 csr._minstret_T_3\[43\] VGND VGND VPWR VPWR net2501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1540 decode.regfile.registers_18\[17\] VGND VGND VPWR VPWR net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2285 decode.regfile.registers_6\[28\] VGND VGND VPWR VPWR net2512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 csr.mscratch\[12\] VGND VGND VPWR VPWR net1778 sky130_fd_sc_hd__dlygate4sd3_1
X_26724_ _09402_ _09720_ VGND VGND VPWR VPWR _09727_ sky130_fd_sc_hd__nand2_1
Xhold2296 decode.regfile.registers_24\[19\] VGND VGND VPWR VPWR net2523 sky130_fd_sc_hd__dlygate4sd3_1
X_29512_ clknet_leaf_267_clock _02525_ VGND VGND VPWR VPWR decode.regfile.registers_8\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1562 fetch.bht.bhtTable_target_pc\[14\]\[15\] VGND VGND VPWR VPWR net1789 sky130_fd_sc_hd__dlygate4sd3_1
X_23936_ _08138_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1573 csr._mcycle_T_3\[32\] VGND VGND VPWR VPWR net1800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1584 execute.csr_write_address_out_reg\[0\] VGND VGND VPWR VPWR net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1595 fetch.bht.bhtTable_target_pc\[15\]\[3\] VGND VGND VPWR VPWR net1822 sky130_fd_sc_hd__dlygate4sd3_1
X_29443_ clknet_leaf_253_clock _02456_ VGND VGND VPWR VPWR decode.regfile.registers_6\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_26655_ net1724 _09679_ _09686_ _09675_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__o211a_1
X_23867_ execute.io_target_pc\[24\] VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__buf_2
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13620_ _09980_ VGND VGND VPWR VPWR _09981_ sky130_fd_sc_hd__buf_4
X_25606_ _09025_ _09069_ VGND VGND VPWR VPWR _09070_ sky130_fd_sc_hd__nand2_1
X_22818_ _07304_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__clkbuf_1
X_29374_ clknet_leaf_255_clock _02387_ VGND VGND VPWR VPWR decode.regfile.registers_4\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_26586_ _09415_ _09645_ VGND VGND VPWR VPWR _09647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23798_ _08052_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28325_ clknet_leaf_192_clock _01338_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25537_ _08912_ _09026_ VGND VGND VPWR VPWR _09030_ sky130_fd_sc_hd__nand2_1
X_13551_ execute.io_mem_rd\[0\] execute.io_mem_rd\[1\] VGND VGND VPWR VPWR _09918_
+ sky130_fd_sc_hd__nor2_1
X_22749_ _07267_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28256_ clknet_leaf_92_clock _01278_ VGND VGND VPWR VPWR csr._minstret_T_3\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_16270_ decode.regfile.registers_1\[25\] _11300_ VGND VGND VPWR VPWR _12242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25468_ _08920_ _08980_ VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27207_ clknet_leaf_363_clock _00236_ VGND VGND VPWR VPWR decode.regfile.registers_28\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15221_ _11058_ _10633_ _10642_ _11085_ VGND VGND VPWR VPWR _11218_ sky130_fd_sc_hd__or4_4
X_24419_ _10556_ _10557_ _09900_ _09917_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__or4b_4
X_28187_ clknet_leaf_85_clock _01209_ VGND VGND VPWR VPWR csr.io_mret_vector\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25399_ net2664 _08928_ _08942_ _08927_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15152_ _11148_ VGND VGND VPWR VPWR _11149_ sky130_fd_sc_hd__buf_6
X_27138_ clknet_leaf_358_clock _00167_ VGND VGND VPWR VPWR decode.regfile.registers_26\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14103_ net2316 _10315_ _10318_ _10317_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19960_ _05212_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27069_ clknet_leaf_346_clock _00098_ VGND VGND VPWR VPWR decode.regfile.registers_24\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_15083_ _11072_ VGND VGND VPWR VPWR _11080_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14034_ _10112_ _10268_ VGND VGND VPWR VPWR _10278_ sky130_fd_sc_hd__nand2_1
X_18911_ _03708_ decode.id_ex_imm_reg\[16\] _04209_ _03932_ VGND VGND VPWR VPWR _04210_
+ sky130_fd_sc_hd__a211o_1
X_19891_ _05158_ _05159_ _03865_ _04526_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_120_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18842_ _03707_ _04139_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_224_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15985_ decode.regfile.registers_13\[17\] _11276_ _11407_ decode.regfile.registers_12\[17\]
+ _11964_ VGND VGND VPWR VPWR _11965_ sky130_fd_sc_hd__a221o_1
X_18773_ decode.id_ex_rs2_data_reg\[6\] _03746_ _03764_ _04068_ _04071_ VGND VGND
+ VPWR VPWR _04072_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_220_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_220_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14936_ decode.control.io_opcode\[5\] VGND VGND VPWR VPWR _10965_ sky130_fd_sc_hd__buf_2
X_17724_ _12498_ _12504_ _12649_ decode.regfile.registers_11\[23\] VGND VGND VPWR
+ VPWR _03128_ sky130_fd_sc_hd__or4b_1
XFILLER_0_76_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14867_ _10909_ VGND VGND VPWR VPWR _10910_ sky130_fd_sc_hd__buf_4
X_17655_ decode.regfile.registers_22\[21\] _12527_ _03059_ _03060_ _12686_ VGND VGND
+ VPWR VPWR _03061_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_19_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16606_ _12570_ VGND VGND VPWR VPWR _12571_ sky130_fd_sc_hd__clkbuf_4
X_13818_ _09930_ _10149_ _10150_ _09935_ VGND VGND VPWR VPWR _10151_ sky130_fd_sc_hd__and4_1
XFILLER_0_203_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17586_ _13221_ _02989_ _02991_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14798_ _10824_ _10825_ _10827_ _10839_ _10840_ VGND VGND VPWR VPWR _10841_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_202_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16537_ _12501_ VGND VGND VPWR VPWR _12502_ sky130_fd_sc_hd__clkbuf_4
X_19325_ _04454_ _04612_ _04613_ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__a31oi_1
X_13749_ _10092_ _10075_ VGND VGND VPWR VPWR _10093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19256_ _04295_ _04546_ _04301_ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__or4b_2
X_16468_ decode.regfile.registers_16\[30\] _11123_ _12418_ _12434_ VGND VGND VPWR
+ VPWR _12435_ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18207_ _10944_ _03528_ _03533_ _03534_ _03544_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__o41a_1
X_15419_ decode.regfile.registers_2\[3\] _10646_ _11298_ VGND VGND VPWR VPWR _11413_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_72_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19187_ _04381_ _03998_ _03997_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_113_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16399_ decode.regfile.registers_18\[28\] _11269_ _12366_ _12367_ _11456_ VGND VGND
+ VPWR VPWR _12368_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18138_ _03495_ _03493_ _03487_ net2138 VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_147_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18069_ _10579_ _10964_ _10580_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__and3b_2
XFILLER_0_145_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold147 io_fetch_data[31] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20100_ _05310_ _05312_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__xnor2_1
Xhold158 io_fetch_data[29] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold169 fetch.bht.bhtTable_valid\[7\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21080_ execute.csr_read_data_out_reg\[28\] _06025_ _03583_ VGND VGND VPWR VPWR _06027_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_106_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20031_ _05231_ _00552_ _05247_ _05253_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_6_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24770_ _08064_ net1986 _08563_ VGND VGND VPWR VPWR _08571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_15 _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21982_ net806 _06587_ _06594_ _06592_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__o211a_1
XINSDIODE1_26 _04589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_37 _08943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23721_ _08011_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__clkbuf_1
XINSDIODE1_48 _09956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_59 _10091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20933_ _05947_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26440_ _09422_ _09558_ VGND VGND VPWR VPWR _09563_ sky130_fd_sc_hd__nand2_1
X_23652_ _07974_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ _05909_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22603_ _10576_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26371_ _09428_ _09515_ VGND VGND VPWR VPWR _09523_ sky130_fd_sc_hd__nand2_1
X_23583_ _07936_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20795_ execute.io_mem_rd\[3\] _05867_ _05868_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__and3_1
X_28110_ clknet_leaf_80_clock _01132_ VGND VGND VPWR VPWR csr.minstret\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25322_ _08891_ decode.regfile.registers_0\[22\] VGND VGND VPWR VPWR _08892_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22534_ _07121_ _07122_ _07126_ _07127_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__a31o_1
XFILLER_0_174_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29090_ clknet_leaf_71_clock _02103_ VGND VGND VPWR VPWR csr._mcycle_T_3\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28041_ clknet_leaf_52_clock _01063_ VGND VGND VPWR VPWR decode.control.io_opcode\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25253_ _08856_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22465_ _07018_ _07035_ _07059_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__and3b_1
XFILLER_0_91_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24204_ _08276_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21416_ _06107_ net1401 _06219_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25184_ _10573_ net2623 _08820_ VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22396_ net73 _06990_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24135_ net1307 execute.io_target_pc\[22\] _08232_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21347_ _06184_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24066_ net1346 VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28943_ clknet_leaf_107_clock _01956_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21278_ _10759_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__buf_2
Xhold670 decode.regfile.registers_26\[0\] VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 execute.csr_write_data_out_reg\[2\] VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 fetch.bht.bhtTable_target_pc\[4\]\[16\] VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlygate4sd3_1
X_23017_ _07097_ _07456_ _07460_ _07462_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_120_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20229_ _05417_ _05238_ _05421_ _05414_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28874_ clknet_leaf_100_clock _01887_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27825_ clknet_leaf_318_clock _00854_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2060 fetch.bht.bhtTable_tag\[7\]\[3\] VGND VGND VPWR VPWR net2287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2071 decode.io_id_pc\[25\] VGND VGND VPWR VPWR net2298 sky130_fd_sc_hd__dlygate4sd3_1
X_15770_ _10959_ VGND VGND VPWR VPWR _11756_ sky130_fd_sc_hd__clkbuf_4
Xhold2082 decode.regfile.registers_21\[24\] VGND VGND VPWR VPWR net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2093 fetch.bht.bhtTable_tag\[12\]\[14\] VGND VGND VPWR VPWR net2320 sky130_fd_sc_hd__dlygate4sd3_1
X_27756_ clknet_leaf_321_clock _00785_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_24968_ csr._mcycle_T_3\[58\] csr._mcycle_T_3\[57\] _08689_ VGND VGND VPWR VPWR _08692_
+ sky130_fd_sc_hd__and3_1
Xhold1370 decode.regfile.registers_6\[29\] VGND VGND VPWR VPWR net1597 sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ csr.io_mem_pc\[13\] csr.io_mem_pc\[14\] csr.io_mem_pc\[15\] _10763_ VGND
+ VGND VPWR VPWR _10764_ sky130_fd_sc_hd__and4_1
Xhold1381 decode.regfile.registers_12\[19\] VGND VGND VPWR VPWR net1608 sky130_fd_sc_hd__dlygate4sd3_1
X_23919_ _08129_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__clkbuf_1
X_26707_ net733 _09709_ _09716_ _09717_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__o211a_1
Xhold1392 fetch.bht.bhtTable_target_pc\[2\]\[20\] VGND VGND VPWR VPWR net1619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27687_ clknet_leaf_27_clock _00716_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_24899_ _07199_ net621 _08647_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__nor3_1
XFILLER_0_58_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17440_ decode.regfile.registers_8\[16\] _12726_ _12601_ VGND VGND VPWR VPWR _13389_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_197_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14652_ _10694_ execute.io_target_pc\[12\] VGND VGND VPWR VPWR _10695_ sky130_fd_sc_hd__and2_1
X_26638_ net1086 _09665_ _09677_ _09675_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__o211a_1
X_29426_ clknet_leaf_260_clock _02439_ VGND VGND VPWR VPWR decode.regfile.registers_5\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13603_ _09939_ memory.io_wb_aluresult\[2\] _09940_ VGND VGND VPWR VPWR _09966_ sky130_fd_sc_hd__a21o_1
X_17371_ _12599_ _13320_ _13321_ VGND VGND VPWR VPWR _13322_ sky130_fd_sc_hd__o21a_1
Xclkbuf_5_29__f_clock clknet_2_3_0_clock VGND VGND VPWR VPWR clknet_5_29__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_29357_ clknet_leaf_226_clock _02370_ VGND VGND VPWR VPWR decode.regfile.registers_3\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_26569_ _09398_ _09632_ VGND VGND VPWR VPWR _09638_ sky130_fd_sc_hd__nand2_1
X_14583_ _10625_ _10613_ VGND VGND VPWR VPWR _10626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19110_ _04407_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__dlymetal6s2s_1
X_16322_ _11048_ _11054_ _11318_ _12292_ VGND VGND VPWR VPWR _12293_ sky130_fd_sc_hd__o31a_1
XFILLER_0_94_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13534_ _09909_ VGND VGND VPWR VPWR _09910_ sky130_fd_sc_hd__buf_4
X_28308_ clknet_leaf_236_clock _01321_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_188_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29288_ clknet_leaf_242_clock _02301_ VGND VGND VPWR VPWR decode.regfile.registers_1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19041_ _04117_ _04100_ _03989_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__mux2_1
X_28239_ clknet_leaf_73_clock _01261_ VGND VGND VPWR VPWR csr._minstret_T_3\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_16253_ decode.regfile.registers_19\[24\] _11406_ _11325_ _12225_ VGND VGND VPWR
+ VPWR _12226_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15204_ _10624_ _11111_ _11045_ _10648_ VGND VGND VPWR VPWR _11201_ sky130_fd_sc_hd__and4_4
XFILLER_0_51_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16184_ _12137_ _12157_ _12158_ VGND VGND VPWR VPWR _12159_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone81 net206 net207 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__nor2_2
XFILLER_0_180_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_226_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15135_ _11131_ VGND VGND VPWR VPWR _11132_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_226_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_310_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_310_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_147_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19943_ _05205_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_1
X_15066_ _10979_ _11050_ _11054_ _11062_ VGND VGND VPWR VPWR _11063_ sky130_fd_sc_hd__or4_4
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_222_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_222_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14017_ _10242_ VGND VGND VPWR VPWR _10268_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19874_ _03789_ _03790_ _05120_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__or3b_1
X_18825_ net130 _03666_ _04123_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_325_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_325_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18756_ _03706_ decode.id_ex_imm_reg\[4\] _04036_ _04037_ VGND VGND VPWR VPWR _04055_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_106_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ decode.regfile.registers_19\[17\] _11406_ VGND VGND VPWR VPWR _11948_ sky130_fd_sc_hd__nor2_1
X_17707_ decode.regfile.registers_20\[23\] _12525_ _12552_ _12823_ _12824_ VGND VGND
+ VPWR VPWR _03111_ sky130_fd_sc_hd__a41o_1
X_14919_ _10667_ VGND VGND VPWR VPWR _10948_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_177_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15899_ decode.regfile.registers_3\[15\] _11110_ _11141_ _11146_ VGND VGND VPWR VPWR
+ _11881_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18687_ _03715_ _03725_ net273 _03978_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_203_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_177_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17638_ decode.regfile.registers_7\[21\] _12612_ _12889_ VGND VGND VPWR VPWR _03044_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17569_ _12566_ _02974_ _02975_ _02976_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19308_ _04503_ _04599_ _04600_ _04346_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20580_ _03554_ _05551_ _05559_ csr.minstret\[19\] VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19239_ _04269_ _04289_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22250_ _06684_ _06844_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21201_ _06086_ _05868_ net448 VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__and3_1
X_22181_ _06624_ _06775_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__and2b_1
XFILLER_0_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21132_ _06050_ _06058_ net719 VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_1197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25940_ net2127 _09256_ _09261_ _09250_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__o211a_1
X_21063_ execute.csr_read_data_out_reg\[20\] _06014_ _06010_ VGND VGND VPWR VPWR _06018_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20014_ _05222_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25871_ _09128_ VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__buf_2
XFILLER_0_225_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24822_ _08598_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__clkbuf_1
X_27610_ clknet_leaf_151_clock _00639_ VGND VGND VPWR VPWR execute.io_target_pc\[19\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_226_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28590_ clknet_leaf_110_clock _01603_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27541_ clknet_leaf_45_clock _00570_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_2
X_24753_ _09900_ _06281_ _09887_ VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__or3b_4
XFILLER_0_154_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21965_ csr._mcycle_T_2\[7\] _06572_ _06584_ _06579_ VGND VGND VPWR VPWR _01227_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23704_ _08002_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27472_ clknet_leaf_53_clock _00501_ VGND VGND VPWR VPWR csr.io_csr_address\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20916_ _05938_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__clkbuf_1
X_24684_ _08525_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21896_ csr.io_mret_vector\[18\] csr.io_mem_pc\[18\] _06515_ VGND VGND VPWR VPWR
+ _06537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29211_ clknet_leaf_130_clock _02224_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_26423_ net2071 _09548_ _09552_ _09553_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23635_ _07965_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__clkbuf_1
X_20847_ _05900_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29142_ clknet_leaf_91_clock _02155_ VGND VGND VPWR VPWR csr.mcycle\[26\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_181_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26354_ net2720 _09505_ _09513_ _09512_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__o211a_1
X_23566_ net2792 _07917_ _07927_ _05805_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_61_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20778_ net100 net133 VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__nand2_1
X_25305_ _08883_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22517_ _07110_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__buf_4
XFILLER_0_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29073_ clknet_leaf_193_clock _02086_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26285_ _09415_ _09472_ VGND VGND VPWR VPWR _09474_ sky130_fd_sc_hd__nand2_1
X_23497_ net2280 _07876_ _07887_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28024_ clknet_leaf_204_clock _01046_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_25236_ _08847_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__clkbuf_1
X_22448_ _06674_ fetch.btb.btbTable\[7\]\[1\] fetch.bht.bhtTable_valid\[7\] _06626_
+ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25167_ _10573_ net2514 _08811_ VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__mux2_1
X_22379_ _06970_ _06972_ _06973_ _06790_ _06641_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24118_ _06426_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25098_ _06115_ net1641 _08596_ VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28926_ clknet_leaf_131_clock _01939_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24049_ _08196_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__clkbuf_1
X_16940_ _12900_ VGND VGND VPWR VPWR _12901_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28857_ clknet_leaf_128_clock _01870_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_16871_ _12597_ _10934_ _10605_ _10607_ VGND VGND VPWR VPWR _12833_ sky130_fd_sc_hd__and4_1
XFILLER_0_216_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18610_ _10067_ _10066_ memory.csr_read_data_out_reg\[17\] _09986_ VGND VGND VPWR
+ VPWR _03909_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_217_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15822_ _10645_ _11147_ _11804_ _11805_ VGND VGND VPWR VPWR _11806_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_126_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27808_ clknet_leaf_327_clock _00837_ VGND VGND VPWR VPWR memory.io_wb_readdata\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19590_ _04859_ _04871_ _04465_ _04198_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__o2bb2a_1
X_28788_ clknet_leaf_118_clock _01801_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15753_ decode.regfile.registers_9\[11\] _11547_ _11737_ _11738_ _11509_ VGND VGND
+ VPWR VPWR _11739_ sky130_fd_sc_hd__a221o_1
X_18541_ execute.csr_read_data_out_reg\[24\] _03661_ _03660_ VGND VGND VPWR VPWR _03840_
+ sky130_fd_sc_hd__or3_1
X_27739_ clknet_leaf_37_clock _00768_ VGND VGND VPWR VPWR decode.io_wb_rd\[2\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_172_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14704_ decode.id_ex_pc_reg\[3\] VGND VGND VPWR VPWR _10747_ sky130_fd_sc_hd__clkbuf_4
X_15684_ decode.regfile.registers_22\[9\] _11096_ _11232_ _11671_ VGND VGND VPWR VPWR
+ _11672_ sky130_fd_sc_hd__a211o_1
X_18472_ _03768_ _03769_ _03770_ net232 VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__o31a_4
XFILLER_0_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14635_ decode.id_ex_pc_reg\[6\] VGND VGND VPWR VPWR _10678_ sky130_fd_sc_hd__clkbuf_4
X_17423_ _13091_ _13176_ decode.regfile.registers_27\[15\] _13050_ VGND VGND VPWR
+ VPWR _13373_ sky130_fd_sc_hd__or4_1
X_29409_ clknet_leaf_247_clock _02422_ VGND VGND VPWR VPWR decode.regfile.registers_5\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_215_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17354_ _10926_ decode.regfile.registers_22\[14\] _12554_ _11009_ _12546_ VGND VGND
+ VPWR VPWR _13305_ sky130_fd_sc_hd__o2111a_1
X_14566_ _10608_ VGND VGND VPWR VPWR _10609_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13517_ _09895_ VGND VGND VPWR VPWR _09896_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16305_ decode.regfile.registers_15\[26\] _11036_ _11205_ _11203_ VGND VGND VPWR
+ VPWR _12276_ sky130_fd_sc_hd__a31o_1
X_17285_ decode.regfile.registers_11\[12\] _12878_ _12772_ _12541_ _13237_ VGND VGND
+ VPWR VPWR _13238_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14497_ net445 _10533_ _10544_ _10535_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16236_ decode.regfile.registers_1\[24\] decode.regfile.registers_0\[24\] _11371_
+ VGND VGND VPWR VPWR _12209_ sky130_fd_sc_hd__mux2_1
X_19024_ _04027_ _04320_ _04322_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16167_ decode.regfile.registers_3\[22\] _11614_ _12140_ _12141_ _11146_ VGND VGND
+ VPWR VPWR _12142_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15118_ decode.immGen._imm_T_24\[1\] decode.immGen._imm_T_24\[11\] VGND VGND VPWR
+ VPWR _11115_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_11_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16098_ _11194_ decode.regfile.registers_12\[20\] decode.regfile.registers_13\[20\]
+ _11196_ _12074_ VGND VGND VPWR VPWR _12075_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15049_ _11045_ VGND VGND VPWR VPWR _11046_ sky130_fd_sc_hd__clkbuf_4
X_19926_ _04620_ _04408_ _04505_ _05193_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__o22a_1
XFILLER_0_220_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_264_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_264_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19857_ _03803_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_179_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18808_ _04106_ _04104_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__nand2_4
XFILLER_0_208_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19788_ _04297_ _04261_ _04263_ _05061_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_69_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18739_ _03889_ decode.id_ex_imm_reg\[4\] _04036_ _04037_ VGND VGND VPWR VPWR _04038_
+ sky130_fd_sc_hd__o2bb2ai_4
Xclkbuf_leaf_279_clock clknet_5_21__leaf_clock VGND VGND VPWR VPWR clknet_leaf_279_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21750_ _06437_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20701_ _03728_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__buf_2
X_21681_ _06384_ _06386_ _06387_ _06352_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_148_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_202_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_202_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_176_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23420_ _03592_ _07841_ _07064_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__a21o_1
X_20632_ csr.mcycle\[27\] _05587_ _05594_ csr.minstret\[27\] VGND VGND VPWR VPWR _05765_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23351_ fetch.bht.bhtTable_target_pc\[8\]\[27\] fetch.bht.bhtTable_target_pc\[9\]\[27\]
+ fetch.bht.bhtTable_target_pc\[10\]\[27\] fetch.bht.bhtTable_target_pc\[11\]\[27\]
+ _07555_ _07710_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20563_ _05627_ csr.io_mret_vector\[17\] _05603_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22302_ net224 _06767_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_8_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_229_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26070_ _08916_ _09330_ VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__nand2_1
X_23282_ fetch.bht.bhtTable_target_pc\[4\]\[22\] fetch.bht.bhtTable_target_pc\[5\]\[22\]
+ fetch.bht.bhtTable_target_pc\[6\]\[22\] fetch.bht.bhtTable_target_pc\[7\]\[22\]
+ _07708_ _07103_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_217_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_217_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20494_ _05591_ _03741_ _05528_ _05595_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_95_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25021_ _10019_ _08726_ _08727_ VGND VGND VPWR VPWR _08728_ sky130_fd_sc_hd__and3_1
X_22233_ fetch.bht.bhtTable_tag\[14\]\[15\] fetch.bht.bhtTable_tag\[15\]\[15\] _06680_
+ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22164_ _06758_ _06685_ _06687_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21115_ _06049_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__clkbuf_1
X_29760_ clknet_leaf_309_clock _02773_ VGND VGND VPWR VPWR decode.regfile.registers_16\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_22095_ _06621_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__buf_4
XFILLER_0_160_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26972_ net2027 _09866_ _09869_ _09865_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__o211a_1
Xfanout221 net83 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_4
XFILLER_0_227_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28711_ clknet_leaf_118_clock _01724_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25923_ _08920_ _09243_ VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__nand2_1
X_21046_ _06008_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__clkbuf_1
X_29691_ clknet_leaf_289_clock _02704_ VGND VGND VPWR VPWR decode.regfile.registers_14\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28642_ clknet_leaf_133_clock _01655_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25854_ net633 _09199_ _09212_ _09209_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24805_ _08589_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28573_ clknet_leaf_191_clock _01586_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_25785_ _08933_ _09166_ VGND VGND VPWR VPWR _09173_ sky130_fd_sc_hd__nand2_1
X_22997_ fetch.bht.bhtTable_target_pc\[8\]\[6\] fetch.bht.bhtTable_target_pc\[9\]\[6\]
+ fetch.bht.bhtTable_target_pc\[10\]\[6\] fetch.bht.bhtTable_target_pc\[11\]\[6\]
+ _07108_ _07125_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__mux4_1
XFILLER_0_213_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24736_ _08552_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27524_ clknet_leaf_43_clock _00553_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_179_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21948_ net830 _06574_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27455_ clknet_leaf_137_clock _00484_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24667_ net1500 execute.io_target_pc\[22\] _08508_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21879_ csr._mcycle_T_2\[12\] _06521_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26406_ net743 _09534_ _09543_ _09540_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__o211a_1
X_14420_ net635 _10490_ _10500_ _10494_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__o211a_1
X_23618_ _07955_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27386_ clknet_leaf_10_clock _00415_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[27\]
+ sky130_fd_sc_hd__dfxtp_2
X_24598_ net1703 VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__clkbuf_1
X_29125_ clknet_leaf_76_clock _02138_ VGND VGND VPWR VPWR csr.mcycle\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_135_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26337_ _09392_ _09502_ VGND VGND VPWR VPWR _09504_ sky130_fd_sc_hd__nand2_1
X_14351_ net500 _10420_ _10460_ _10453_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_210_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23549_ net2171 _07918_ _07915_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__or3b_1
XFILLER_0_108_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_210_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29056_ clknet_leaf_170_clock _02069_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17070_ decode.regfile.registers_13\[7\] _12775_ _12663_ VGND VGND VPWR VPWR _13028_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26268_ net2421 _09462_ _09464_ _09458_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__o211a_1
X_14282_ _09964_ _10420_ VGND VGND VPWR VPWR _10422_ sky130_fd_sc_hd__nand2_1
X_16021_ decode.regfile.registers_13\[18\] _11046_ _11690_ _11987_ _11999_ VGND VGND
+ VPWR VPWR _12000_ sky130_fd_sc_hd__o32a_1
X_25219_ _08057_ net1599 _08837_ VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__mux2_1
X_28007_ clknet_leaf_195_clock _01029_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26199_ _09372_ VGND VGND VPWR VPWR _09419_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_208_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17972_ _10939_ _03068_ decode.regfile.registers_27\[29\] _12506_ VGND VGND VPWR
+ VPWR _03370_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19711_ _04618_ net219 _04982_ _04949_ _04987_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__a311o_1
X_28909_ clknet_leaf_102_clock _01922_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16923_ decode.regfile.registers_1\[4\] _12778_ _12830_ _12882_ _12883_ VGND VGND
+ VPWR VPWR _12884_ sky130_fd_sc_hd__o221a_1
X_29889_ clknet_leaf_304_clock _02902_ VGND VGND VPWR VPWR decode.regfile.registers_20\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_204_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19642_ _04244_ _04302_ _04921_ _04308_ _04206_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__o32a_1
XFILLER_0_189_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16854_ _10940_ _12706_ decode.regfile.registers_27\[2\] _12507_ VGND VGND VPWR VPWR
+ _12817_ sky130_fd_sc_hd__or4_1
X_15805_ decode.regfile.registers_23\[12\] _11088_ _11764_ _11789_ VGND VGND VPWR
+ VPWR _11790_ sky130_fd_sc_hd__o22a_1
X_19573_ _04618_ _04386_ _04855_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__o21ai_2
X_13997_ _10025_ _10255_ VGND VGND VPWR VPWR _10257_ sky130_fd_sc_hd__nand2_1
X_16785_ _12658_ _12746_ _12747_ _12748_ VGND VGND VPWR VPWR _12749_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_217_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18524_ net239 _03797_ _10121_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__or3b_1
XFILLER_0_88_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15736_ _11038_ VGND VGND VPWR VPWR _11722_ sky130_fd_sc_hd__buf_2
XFILLER_0_150_1320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18455_ execute.io_mem_rd\[4\] csr.io_csr_address\[4\] VGND VGND VPWR VPWR _03754_
+ sky130_fd_sc_hd__or2_1
X_15667_ _11156_ _11653_ _11654_ VGND VGND VPWR VPWR _11655_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17406_ decode.regfile.registers_13\[15\] _12775_ _13354_ _13355_ _12663_ VGND VGND
+ VPWR VPWR _13356_ sky130_fd_sc_hd__a221o_1
X_14618_ _10660_ decode.id_ex_ex_rd_reg\[3\] VGND VGND VPWR VPWR _10661_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15598_ decode.regfile.registers_10\[7\] _10638_ _11132_ _11575_ _11587_ VGND VGND
+ VPWR VPWR _11588_ sky130_fd_sc_hd__o32a_1
X_18386_ _03679_ _03682_ _03683_ _03684_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_172_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14549_ _10591_ VGND VGND VPWR VPWR _10592_ sky130_fd_sc_hd__clkbuf_4
X_17337_ _12686_ VGND VGND VPWR VPWR _13289_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17268_ _12495_ VGND VGND VPWR VPWR _13221_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_168_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19007_ _03635_ _03634_ _03633_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_70_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16219_ decode.regfile.registers_19\[23\] _11453_ _11219_ _12192_ VGND VGND VPWR
+ VPWR _12193_ sky130_fd_sc_hd__o211a_1
X_17199_ _12594_ _13152_ _13153_ _12590_ VGND VGND VPWR VPWR _13154_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_141_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19909_ net339 _05157_ _05177_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_209_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1903 fetch.bht.bhtTable_tag\[0\]\[10\] VGND VGND VPWR VPWR net2130 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1914 fetch.bht.bhtTable_target_pc\[15\]\[30\] VGND VGND VPWR VPWR net2141 sky130_fd_sc_hd__dlygate4sd3_1
X_22920_ _07080_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__buf_6
Xhold1925 decode.io_id_pc\[18\] VGND VGND VPWR VPWR net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1936 decode.regfile.registers_3\[4\] VGND VGND VPWR VPWR net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1947 decode.regfile.registers_7\[30\] VGND VGND VPWR VPWR net2174 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_3_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1958 decode.regfile.registers_2\[31\] VGND VGND VPWR VPWR net2185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1969 decode.regfile.registers_3\[22\] VGND VGND VPWR VPWR net2196 sky130_fd_sc_hd__dlygate4sd3_1
X_22851_ _07321_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21802_ csr.io_csr_write_address\[6\] _06469_ _06458_ VGND VGND VPWR VPWR _06470_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_91_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25570_ net2279 _09039_ _09048_ _09046_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__o211a_1
X_22782_ _07284_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24521_ _08081_ net1667 _08439_ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_141_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_141_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21733_ net1114 _10820_ _06428_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27240_ clknet_leaf_0_clock _00269_ VGND VGND VPWR VPWR decode.regfile.registers_29\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_24452_ _08405_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21664_ csr.minstret\[17\] csr.minstret\[18\] _06370_ VGND VGND VPWR VPWR _06375_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_164_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23403_ execute.io_target_pc\[30\] _10757_ _07088_ _07825_ _10971_ VGND VGND VPWR
+ VPWR _07826_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20615_ csr.minstret\[24\] _05574_ _05586_ csr.mcycle\[24\] VGND VGND VPWR VPWR _05751_
+ sky130_fd_sc_hd__a22o_1
X_27171_ clknet_leaf_362_clock _00200_ VGND VGND VPWR VPWR decode.regfile.registers_27\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_24383_ net1213 execute.io_target_pc\[14\] _08367_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__mux2_1
X_21595_ net559 _06321_ _06323_ csr.minstret\[0\] VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__a211oi_1
Xclkbuf_leaf_156_clock clknet_5_24__leaf_clock VGND VGND VPWR VPWR clknet_leaf_156_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26122_ _08968_ _09328_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__nand2_1
X_23334_ net220 _07706_ _07707_ _07761_ _07705_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_10_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_49_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20546_ csr.minstret\[15\] VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__buf_2
XFILLER_0_149_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26053_ _08975_ _09285_ VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__nand2_1
X_23265_ _07694_ _07075_ _07696_ _06740_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20477_ csr.mcycle\[6\] _05552_ _05575_ csr.minstret\[6\] VGND VGND VPWR VPWR _05631_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25004_ csr.mcycle\[6\] _03558_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_197_Right_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22216_ _06631_ _06810_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23196_ csr._csr_read_data_T_8\[17\] _06480_ csr.io_mret_vector\[17\] _07621_ _07631_
+ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__o221a_1
XFILLER_0_162_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29812_ clknet_leaf_295_clock _02825_ VGND VGND VPWR VPWR decode.regfile.registers_17\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22147_ _06632_ _06741_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1090 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29743_ clknet_leaf_285_clock _02756_ VGND VGND VPWR VPWR decode.regfile.registers_15\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22078_ _06672_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__buf_4
X_26955_ net528 _09853_ _09859_ _09852_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13920_ _10025_ _10210_ VGND VGND VPWR VPWR _10212_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_58_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25906_ _09241_ VGND VGND VPWR VPWR _09242_ sky130_fd_sc_hd__buf_2
X_21029_ _05999_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
X_29674_ clknet_leaf_277_clock _02687_ VGND VGND VPWR VPWR decode.regfile.registers_13\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_26886_ _09412_ _09819_ VGND VGND VPWR VPWR _09820_ sky130_fd_sc_hd__nand2_1
X_28625_ clknet_leaf_104_clock _01638_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_13851_ _10048_ _10164_ VGND VGND VPWR VPWR _10171_ sky130_fd_sc_hd__nand2_1
X_25837_ _08910_ _09200_ VGND VGND VPWR VPWR _09203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28556_ clknet_leaf_219_clock _01569_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16570_ _12534_ VGND VGND VPWR VPWR _12535_ sky130_fd_sc_hd__buf_4
X_13782_ memory.io_wb_reg_pc\[27\] _10001_ _10005_ _10119_ VGND VGND VPWR VPWR _10120_
+ sky130_fd_sc_hd__a211o_1
X_25768_ _08916_ _09157_ VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_109_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_109_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15521_ _11511_ _11512_ VGND VGND VPWR VPWR _11513_ sky130_fd_sc_hd__and2_1
X_27507_ clknet_leaf_20_clock _00536_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dfxtp_1
X_24719_ _08081_ net1807 _08542_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28487_ clknet_leaf_204_clock _01500_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25699_ _08922_ _09122_ VGND VGND VPWR VPWR _09123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18240_ csr._mcycle_T_3\[33\] csr._mcycle_T_3\[32\] csr.mcycle\[31\] VGND VGND VPWR
+ VPWR _03575_ sky130_fd_sc_hd__or3_1
XFILLER_0_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15452_ _11398_ VGND VGND VPWR VPWR _11445_ sky130_fd_sc_hd__clkbuf_4
X_27438_ clknet_leaf_145_clock _00467_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_167_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14403_ net936 _10490_ _10491_ _10481_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18171_ _03513_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_67_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15383_ _11308_ VGND VGND VPWR VPWR _11378_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27369_ clknet_leaf_33_clock _00398_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17122_ decode.regfile.registers_21\[8\] _12682_ _12909_ VGND VGND VPWR VPWR _13079_
+ sky130_fd_sc_hd__o21a_1
X_14334_ net740 _10447_ _10451_ _10440_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__o211a_1
X_29108_ clknet_leaf_16_clock _02121_ VGND VGND VPWR VPWR csr._mcycle_T_3\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17053_ _12575_ VGND VGND VPWR VPWR _13011_ sky130_fd_sc_hd__clkbuf_4
X_29039_ clknet_leaf_107_clock _02052_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14265_ net664 _10403_ _10410_ _10411_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__o211a_1
Xmax_cap207 net208 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_4
Xmax_cap218 _05523_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_1
X_16004_ _11942_ decode.regfile.registers_30\[18\] _11722_ _11723_ _11724_ VGND VGND
+ VPWR VPWR _11983_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_208_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14196_ _10142_ _10331_ VGND VGND VPWR VPWR _10371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_206_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17955_ _12498_ _12977_ _12649_ decode.regfile.registers_11\[29\] VGND VGND VPWR
+ VPWR _03353_ sky130_fd_sc_hd__or4b_1
XFILLER_0_225_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16906_ _10940_ _12706_ decode.regfile.registers_27\[3\] _12507_ VGND VGND VPWR VPWR
+ _12868_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17886_ _03265_ _03285_ _12565_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19625_ _03594_ _04345_ _03636_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__and3_1
XFILLER_0_205_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16837_ decode.regfile.registers_16\[2\] _12576_ _12799_ VGND VGND VPWR VPWR _12800_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_221_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_215_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19556_ _04180_ net254 _04837_ _04838_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_215_1147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16768_ _12731_ VGND VGND VPWR VPWR _12732_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18507_ _03656_ _03805_ decode.id_ex_rs1_data_reg\[26\] _03689_ VGND VGND VPWR VPWR
+ _03806_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_157_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15719_ _11705_ decode.regfile.registers_13\[10\] _11276_ VGND VGND VPWR VPWR _11706_
+ sky130_fd_sc_hd__mux2_1
X_19487_ _04618_ _04294_ _04620_ _04772_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_83_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16699_ _12663_ VGND VGND VPWR VPWR _12664_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_83_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18438_ csr.io_csr_address\[1\] VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_73_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18369_ execute.io_mem_memtoreg\[1\] execute.io_mem_memtoreg\[0\] execute.io_reg_pc\[31\]
+ _03667_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_21_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20400_ csr.io_csr_address\[11\] _05526_ net218 _05520_ _05559_ VGND VGND VPWR VPWR
+ _05560_ sky130_fd_sc_hd__a41o_1
XFILLER_0_16_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21380_ _06128_ net2216 _06199_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20331_ _10790_ decode.id_ex_pc_reg\[26\] _05494_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_88_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_187_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23050_ _07122_ _07493_ _07127_ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20262_ _05417_ _05281_ _05447_ _05414_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22001_ net1093 _06600_ _06604_ _06605_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20193_ _05391_ _05383_ _05386_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_11_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_11_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_179_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2401 decode.regfile.registers_2\[24\] VGND VGND VPWR VPWR net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2412 decode.regfile.registers_9\[22\] VGND VGND VPWR VPWR net2639 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2423 decode.regfile.registers_6\[5\] VGND VGND VPWR VPWR net2650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2434 decode.regfile.registers_15\[25\] VGND VGND VPWR VPWR net2661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2445 decode.regfile.registers_4\[20\] VGND VGND VPWR VPWR net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1700 decode.regfile.registers_23\[17\] VGND VGND VPWR VPWR net1927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1711 fetch.bht.bhtTable_tag\[14\]\[8\] VGND VGND VPWR VPWR net1938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23952_ _08146_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__clkbuf_1
Xhold2456 decode.regfile.registers_13\[25\] VGND VGND VPWR VPWR net2683 sky130_fd_sc_hd__dlygate4sd3_1
X_26740_ _09708_ VGND VGND VPWR VPWR _09736_ sky130_fd_sc_hd__buf_2
Xhold1722 fetch.bht.bhtTable_target_pc\[14\]\[13\] VGND VGND VPWR VPWR net1949 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2467 decode.regfile.registers_0\[16\] VGND VGND VPWR VPWR net2694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2478 _06334_ VGND VGND VPWR VPWR net2705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 decode.regfile.registers_17\[4\] VGND VGND VPWR VPWR net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1744 fetch.bht.bhtTable_target_pc\[6\]\[22\] VGND VGND VPWR VPWR net1971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2489 decode.regfile.registers_11\[24\] VGND VGND VPWR VPWR net2716 sky130_fd_sc_hd__dlygate4sd3_1
X_22903_ _06944_ _06928_ _07018_ _07353_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__nor4_2
Xhold1755 decode.regfile.registers_11\[6\] VGND VGND VPWR VPWR net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1766 decode.regfile.registers_21\[27\] VGND VGND VPWR VPWR net1993 sky130_fd_sc_hd__dlygate4sd3_1
X_26671_ _09426_ _09689_ VGND VGND VPWR VPWR _09696_ sky130_fd_sc_hd__nand2_1
X_23883_ _08109_ net1336 _07940_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_26_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_26_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1777 decode.regfile.registers_25\[2\] VGND VGND VPWR VPWR net2004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1788 _01246_ VGND VGND VPWR VPWR net2015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1799 fetch.bht.bhtTable_target_pc\[15\]\[25\] VGND VGND VPWR VPWR net2026 sky130_fd_sc_hd__dlygate4sd3_1
X_28410_ clknet_leaf_142_clock _01423_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_168_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22834_ net1646 _10777_ _07308_ VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25622_ net1483 _09068_ _09078_ _09074_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__o211a_1
X_29390_ clknet_leaf_258_clock _02403_ VGND VGND VPWR VPWR decode.regfile.registers_4\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28341_ clknet_leaf_203_clock _01354_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_25553_ _09023_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_49_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22765_ _07275_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24504_ _08064_ net1238 _08428_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21716_ csr._mcycle_T_2\[29\] _06325_ _06413_ csr.minstret\[28\] csr.minstret\[29\]
+ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__a221oi_1
X_28272_ clknet_leaf_61_clock _01294_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25484_ _08935_ _08992_ VGND VGND VPWR VPWR _08999_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22696_ net2774 _07236_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24435_ _08396_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27223_ clknet_leaf_5_clock _00252_ VGND VGND VPWR VPWR decode.regfile.registers_29\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_21647_ csr.minstret\[4\] csr.minstret\[5\] csr.minstret\[14\] _06333_ VGND VGND
+ VPWR VPWR _06362_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27154_ clknet_leaf_353_clock _00183_ VGND VGND VPWR VPWR decode.regfile.registers_27\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_24366_ net1704 execute.io_target_pc\[6\] _08356_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__mux2_1
X_21578_ _06149_ net1964 _06306_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__mux2_1
XANTENNA_70 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 _12076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26105_ _08952_ _09353_ VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23317_ net221 _07706_ _07707_ _07745_ _07705_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__o311a_1
XFILLER_0_133_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_92 decode.regfile.registers_11\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20529_ csr._minstret_T_3\[44\] _05556_ csr.minstret\[12\] _05658_ _05537_ VGND VGND
+ VPWR VPWR _05677_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27085_ clknet_leaf_330_clock _00114_ VGND VGND VPWR VPWR decode.regfile.registers_24\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_24297_ _08324_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14050_ _10286_ VGND VGND VPWR VPWR _10287_ sky130_fd_sc_hd__clkbuf_4
X_26036_ _08958_ _09310_ VGND VGND VPWR VPWR _09317_ sky130_fd_sc_hd__nand2_1
X_23248_ fetch.bht.bhtTable_target_pc\[8\]\[20\] fetch.bht.bhtTable_target_pc\[9\]\[20\]
+ fetch.bht.bhtTable_target_pc\[10\]\[20\] fetch.bht.bhtTable_target_pc\[11\]\[20\]
+ _07669_ _07656_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23179_ csr._csr_read_data_T_8\[16\] _06038_ csr.io_mret_vector\[16\] _06462_ VGND
+ VGND VPWR VPWR _07616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27987_ clknet_leaf_183_clock _01009_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_201_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_201_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17740_ _10929_ decode.regfile.registers_28\[23\] _02992_ VGND VGND VPWR VPWR _03144_
+ sky130_fd_sc_hd__o21a_1
X_29726_ clknet_leaf_312_clock _02739_ VGND VGND VPWR VPWR decode.regfile.registers_15\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_197_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14952_ _10979_ VGND VGND VPWR VPWR _10980_ sky130_fd_sc_hd__clkbuf_4
X_26938_ _10014_ _09849_ VGND VGND VPWR VPWR _09850_ sky130_fd_sc_hd__nand2_1
X_13903_ net2360 _10199_ _10202_ _10188_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17671_ decode.regfile.registers_17\[22\] _11021_ _12559_ _12534_ VGND VGND VPWR
+ VPWR _03076_ sky130_fd_sc_hd__and4_1
X_29657_ clknet_leaf_288_clock _02670_ VGND VGND VPWR VPWR decode.regfile.registers_12\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_193_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14883_ _10915_ VGND VGND VPWR VPWR _10921_ sky130_fd_sc_hd__clkbuf_2
X_26869_ net540 _09809_ _09810_ _09799_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_193_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19410_ _04360_ _04689_ _04694_ _04698_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__a31o_1
X_28608_ clknet_leaf_170_clock _01621_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_16622_ _12582_ VGND VGND VPWR VPWR _12587_ sky130_fd_sc_hd__clkbuf_4
X_13834_ _09999_ _10154_ VGND VGND VPWR VPWR _10161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29588_ clknet_leaf_275_clock _02601_ VGND VGND VPWR VPWR decode.regfile.registers_10\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19341_ _03704_ _04537_ _04345_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28539_ clknet_leaf_210_clock _01552_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_16553_ _10594_ _10604_ _10924_ VGND VGND VPWR VPWR _12518_ sky130_fd_sc_hd__or3b_4
X_13765_ memory.csr_read_data_out_reg\[24\] _09988_ _10104_ _10105_ VGND VGND VPWR
+ VPWR _10106_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_167_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15504_ decode.regfile.registers_14\[5\] _11206_ _11272_ decode.regfile.registers_15\[5\]
+ _11201_ VGND VGND VPWR VPWR _11496_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19272_ _04465_ _04553_ _04565_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13696_ _10047_ VGND VGND VPWR VPWR _10048_ sky130_fd_sc_hd__buf_4
X_16484_ _12133_ net634 _12416_ _12450_ _12132_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_14_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18223_ csr.mcycle\[4\] csr.mcycle\[3\] csr.mcycle\[5\] _03557_ VGND VGND VPWR VPWR
+ _03558_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_152_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15435_ decode.regfile.registers_19\[3\] _11406_ _11325_ _11428_ VGND VGND VPWR VPWR
+ _11429_ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18154_ _03506_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15366_ _11201_ VGND VGND VPWR VPWR _11361_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17105_ decode.regfile.registers_4\[8\] _12549_ _12532_ decode.regfile.registers_5\[8\]
+ _12626_ VGND VGND VPWR VPWR _13062_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_29_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14317_ _10064_ _10431_ VGND VGND VPWR VPWR _10442_ sky130_fd_sc_hd__nand2_1
X_18085_ _03463_ _03467_ _03465_ net2280 VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__and4bb_1
X_15297_ _10645_ decode.immGen._imm_T_24\[3\] decode.immGen._imm_T_24\[1\] decode.immGen._imm_T_24\[2\]
+ VGND VGND VPWR VPWR _11293_ sky130_fd_sc_hd__or4b_4
Xhold307 decode.regfile.registers_23\[28\] VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold318 memory.csr_read_data_out_reg\[11\] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_106_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14248_ _10081_ _10400_ VGND VGND VPWR VPWR _10402_ sky130_fd_sc_hd__nand2_1
X_17036_ _12519_ VGND VGND VPWR VPWR _12995_ sky130_fd_sc_hd__clkbuf_2
Xhold329 decode.regfile.registers_10\[10\] VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_229_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14179_ _10097_ _10355_ VGND VGND VPWR VPWR _10362_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_182_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _03986_ _03985_ _03984_ _03987_ _03703_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__a311o_1
Xhold1007 fetch.bht.bhtTable_tag\[8\]\[14\] VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1018 fetch.bht.bhtTable_target_pc\[5\]\[10\] VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17938_ _12765_ net476 _12486_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1029 csr.mcycle\[6\] VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17869_ decode.regfile.registers_3\[27\] _10615_ _12728_ _12837_ VGND VGND VPWR VPWR
+ _03269_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_1_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19608_ _03912_ _04862_ _04863_ _04201_ _03938_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__a311o_1
XFILLER_0_178_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20880_ _05918_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1088 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19539_ _04225_ _04094_ _04444_ _04091_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__and4_1
XFILLER_0_193_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22550_ csr._minstret_T_3\[34\] _06417_ _07140_ _06422_ VGND VGND VPWR VPWR _07141_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_260 net2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_200_Right_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21501_ _06130_ net1781 _06263_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_271 _10096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_282 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22481_ _07075_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__buf_4
XINSDIODE1_293 _12542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24220_ _08284_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21432_ _06231_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24151_ net2018 execute.io_target_pc\[30\] _06427_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21363_ _06111_ net1671 _06188_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23102_ fetch.bht.bhtTable_target_pc\[12\]\[12\] fetch.bht.bhtTable_target_pc\[13\]\[12\]
+ _07068_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20314_ _10864_ _05482_ decode.id_ex_rdsel_reg VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24082_ _08213_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold830 fetch.bht.bhtTable_target_pc\[10\]\[26\] VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__dlygate4sd3_1
X_21294_ _06155_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold841 fetch.bht.bhtTable_tag\[1\]\[18\] VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 fetch.bht.bhtTable_target_pc\[3\]\[27\] VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23033_ fetch.bht.bhtTable_target_pc\[8\]\[8\] fetch.bht.bhtTable_target_pc\[9\]\[8\]
+ _07407_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27910_ clknet_leaf_19_clock _00939_ VGND VGND VPWR VPWR csr._mcycle_T_2\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20245_ _10704_ _05427_ _10678_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__a21oi_1
Xhold863 decode.regfile.registers_7\[16\] VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__dlygate4sd3_1
X_28890_ clknet_leaf_178_clock _01903_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold874 _08512_ VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold885 fetch.bht.bhtTable_tag\[1\]\[4\] VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold896 fetch.bht.bhtTable_target_pc\[2\]\[30\] VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27841_ clknet_leaf_54_clock _00870_ VGND VGND VPWR VPWR csr.io_mret sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_38_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20176_ _05376_ _05377_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__xnor2_1
Xhold2220 decode.regfile.registers_7\[31\] VGND VGND VPWR VPWR net2447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2231 decode.regfile.registers_26\[11\] VGND VGND VPWR VPWR net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2242 decode.regfile.registers_8\[4\] VGND VGND VPWR VPWR net2469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27772_ clknet_leaf_324_clock _00801_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2253 decode.regfile.registers_5\[23\] VGND VGND VPWR VPWR net2480 sky130_fd_sc_hd__dlygate4sd3_1
X_24984_ _08701_ csr.mcycle\[0\] _06318_ VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__a21oi_1
Xhold2264 decode.regfile.registers_26\[24\] VGND VGND VPWR VPWR net2491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1530 decode.regfile.registers_5\[2\] VGND VGND VPWR VPWR net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2275 decode.regfile.registers_15\[29\] VGND VGND VPWR VPWR net2502 sky130_fd_sc_hd__dlygate4sd3_1
X_29511_ clknet_leaf_265_clock _02524_ VGND VGND VPWR VPWR decode.regfile.registers_8\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1541 fetch.bht.bhtTable_target_pc\[9\]\[6\] VGND VGND VPWR VPWR net1768 sky130_fd_sc_hd__dlygate4sd3_1
X_26723_ net728 _09723_ _09726_ _09717_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__o211a_1
Xhold2286 decode.regfile.registers_20\[23\] VGND VGND VPWR VPWR net2513 sky130_fd_sc_hd__dlygate4sd3_1
X_23935_ net845 _08093_ _08130_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__mux2_1
Xhold1552 _01232_ VGND VGND VPWR VPWR net1779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2297 decode.regfile.registers_12\[14\] VGND VGND VPWR VPWR net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1563 fetch.bht.bhtTable_target_pc\[11\]\[12\] VGND VGND VPWR VPWR net1790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1574 _02097_ VGND VGND VPWR VPWR net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1585 decode.regfile.registers_11\[4\] VGND VGND VPWR VPWR net1812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29442_ clknet_leaf_255_clock _02455_ VGND VGND VPWR VPWR decode.regfile.registers_6\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_23866_ _08098_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__clkbuf_1
Xhold1596 fetch.bht.bhtTable_tag\[13\]\[13\] VGND VGND VPWR VPWR net1823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26654_ _09408_ _09676_ VGND VGND VPWR VPWR _09686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22817_ net1026 _10787_ _07297_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__mux2_1
X_25605_ _09067_ VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__buf_2
XFILLER_0_66_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29373_ clknet_leaf_255_clock _02386_ VGND VGND VPWR VPWR decode.regfile.registers_4\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_23797_ _08051_ net1111 _07952_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__mux2_1
X_26585_ net2201 _09636_ _09646_ _09635_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28324_ clknet_leaf_187_clock _01337_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13550_ _09914_ _09892_ _09917_ net390 VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__a31o_1
X_22748_ _06122_ net1998 _07265_ VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25536_ net686 _09024_ _09029_ _09017_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28255_ clknet_leaf_92_clock _01277_ VGND VGND VPWR VPWR csr._minstret_T_3\[55\]
+ sky130_fd_sc_hd__dfxtp_2
X_25467_ net1976 _08979_ _08988_ _08972_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22679_ csr._mcycle_T_2\[15\] _07223_ VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__or2_1
X_15220_ _11216_ VGND VGND VPWR VPWR _11217_ sky130_fd_sc_hd__clkbuf_4
X_24418_ _08386_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27206_ clknet_leaf_364_clock _00235_ VGND VGND VPWR VPWR decode.regfile.registers_28\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_28186_ clknet_leaf_85_clock _01208_ VGND VGND VPWR VPWR csr.io_mret_vector\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_25398_ _08941_ _08923_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15151_ _11147_ VGND VGND VPWR VPWR _11148_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24349_ _08111_ net1673 _06187_ VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27137_ clknet_leaf_359_clock _00166_ VGND VGND VPWR VPWR decode.regfile.registers_26\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14102_ _10092_ _10312_ VGND VGND VPWR VPWR _10318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15082_ _10990_ VGND VGND VPWR VPWR _11079_ sky130_fd_sc_hd__buf_2
X_27068_ clknet_leaf_345_clock _00097_ VGND VGND VPWR VPWR decode.regfile.registers_24\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14033_ net2565 _10271_ _10277_ _10275_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__o211a_1
X_26019_ net2609 _09300_ _09307_ _09305_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__o211a_1
X_18910_ decode.id_ex_rs1_data_reg\[16\] _03688_ _03925_ _03701_ _03928_ VGND VGND
+ VPWR VPWR _04209_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_129_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19890_ _03781_ _05142_ _05146_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18841_ _03889_ decode.id_ex_imm_reg\[9\] VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_224_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1055 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18772_ _03715_ _03725_ _04067_ _03726_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__o31a_1
X_15984_ _11181_ _11962_ _11963_ VGND VGND VPWR VPWR _11964_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_220_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29709_ clknet_leaf_284_clock _02722_ VGND VGND VPWR VPWR decode.regfile.registers_14\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_17723_ decode.regfile.registers_9\[23\] _12607_ _03125_ _03126_ _12600_ VGND VGND
+ VPWR VPWR _03127_ sky130_fd_sc_hd__a221oi_2
X_14935_ decode.control.io_opcode\[4\] VGND VGND VPWR VPWR _10964_ sky130_fd_sc_hd__buf_2
XFILLER_0_188_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17654_ decode.regfile.registers_21\[21\] _12822_ _12909_ VGND VGND VPWR VPWR _03060_
+ sky130_fd_sc_hd__o21a_1
X_14866_ _10908_ _10758_ VGND VGND VPWR VPWR _10909_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_19_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16605_ _10923_ _12559_ _11020_ _12555_ VGND VGND VPWR VPWR _12570_ sky130_fd_sc_hd__and4b_2
XFILLER_0_202_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13817_ decode.io_wb_rd\[0\] decode.io_wb_rd\[1\] VGND VGND VPWR VPWR _10150_ sky130_fd_sc_hd__and2_4
XFILLER_0_187_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17585_ _13215_ decode.regfile.registers_28\[19\] _02992_ VGND VGND VPWR VPWR _02993_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_225_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14797_ _10816_ _10822_ _10730_ VGND VGND VPWR VPWR _10840_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19324_ _04452_ _04615_ _04505_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16536_ _10934_ _10597_ VGND VGND VPWR VPWR _12501_ sky130_fd_sc_hd__nand2_1
X_13748_ _10091_ VGND VGND VPWR VPWR _10092_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_175_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19255_ _04281_ _04283_ _04548_ _04549_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__o31a_1
XFILLER_0_73_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16467_ _10650_ _10625_ _11053_ _12433_ VGND VGND VPWR VPWR _12434_ sky130_fd_sc_hd__o31a_1
XFILLER_0_112_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13679_ _10012_ _10021_ memory.io_wb_readdata\[11\] VGND VGND VPWR VPWR _10033_ sky130_fd_sc_hd__and3b_1
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18206_ _03540_ _03458_ _10965_ _03543_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15418_ _11154_ decode.regfile.registers_0\[3\] _11156_ _11411_ VGND VGND VPWR VPWR
+ _11412_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19186_ _04251_ _04252_ _04375_ _04481_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__a31o_1
XFILLER_0_182_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16398_ _11225_ _11125_ _11216_ decode.regfile.registers_17\[28\] _11128_ VGND VGND
+ VPWR VPWR _12367_ sky130_fd_sc_hd__o32a_1
XFILLER_0_53_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18137_ _03497_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15349_ _11243_ VGND VGND VPWR VPWR _11344_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_184_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18068_ _03457_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold148 io_fetch_data[30] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold159 io_fetch_data[25] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17019_ decode.regfile.registers_9\[6\] _11018_ _12977_ _12510_ _12653_ VGND VGND
+ VPWR VPWR _12978_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_74_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20030_ _05250_ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__xor2_1
XFILLER_0_226_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21981_ csr.mscratch\[14\] _06588_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_16 _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_27 _05155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23720_ net1350 csr.io_mem_pc\[23\] _08003_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__mux2_1
XINSDIODE1_38 _08945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_49 _09956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20932_ _05937_ _05945_ net51 VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23651_ net1689 _10803_ _07972_ VGND VGND VPWR VPWR _07974_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20863_ net118 _05903_ _05899_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22602_ _06377_ _07176_ _07178_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__nor3_1
XFILLER_0_53_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26370_ net2573 _09518_ _09522_ _09512_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_102_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23582_ _06113_ net1922 _07930_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20794_ _05871_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25321_ _10018_ VGND VGND VPWR VPWR _08891_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22533_ _06740_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25252_ _08091_ net1687 _08848_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28040_ clknet_leaf_51_clock _01062_ VGND VGND VPWR VPWR decode.control.io_opcode\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22464_ _07037_ _07048_ _07058_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24203_ _08097_ net1996 _08266_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21415_ _06222_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25183_ net404 _08820_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__xnor2_1
X_22395_ _06699_ _06981_ _06983_ _06989_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__o31a_1
XFILLER_0_115_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24134_ _08240_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21346_ net1252 _10777_ _06179_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_978 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24065_ net1345 execute.io_target_pc\[20\] _08198_ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__mux2_1
X_28942_ clknet_leaf_87_clock _01955_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold660 fetch.bht.bhtTable_tag\[12\]\[12\] VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__dlygate4sd3_1
X_21277_ _06144_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__clkbuf_1
Xhold671 decode.regfile.registers_21\[19\] VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23016_ _07461_ _07406_ _07085_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__a21oi_1
Xhold682 decode.regfile.registers_21\[13\] VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 fetch.bht.bhtTable_target_pc\[12\]\[9\] VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__dlygate4sd3_1
X_20228_ _05420_ _10834_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_229_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28873_ clknet_leaf_87_clock _01886_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_228_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27824_ clknet_leaf_322_clock _00853_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_20159_ _00570_ _05226_ _05363_ _05239_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__o22a_1
Xhold2050 decode.regfile.registers_17\[28\] VGND VGND VPWR VPWR net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2061 fetch.bht.bhtTable_target_pc\[15\]\[15\] VGND VGND VPWR VPWR net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2072 decode.regfile.registers_18\[23\] VGND VGND VPWR VPWR net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2083 decode.regfile.registers_24\[20\] VGND VGND VPWR VPWR net2310 sky130_fd_sc_hd__dlygate4sd3_1
X_27755_ clknet_leaf_323_clock _00784_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2094 decode.regfile.registers_9\[17\] VGND VGND VPWR VPWR net2321 sky130_fd_sc_hd__dlygate4sd3_1
X_24967_ net949 _08689_ net636 VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_225_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1360 decode.regfile.registers_11\[30\] VGND VGND VPWR VPWR net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 fetch.bht.bhtTable_target_pc\[11\]\[8\] VGND VGND VPWR VPWR net1598 sky130_fd_sc_hd__dlygate4sd3_1
X_14720_ csr.io_mem_pc\[10\] csr.io_mem_pc\[11\] csr.io_mem_pc\[12\] _10762_ VGND
+ VGND VPWR VPWR _10763_ sky130_fd_sc_hd__and4_4
X_26706_ _09701_ VGND VGND VPWR VPWR _09717_ sky130_fd_sc_hd__clkbuf_4
X_23918_ net1288 _08076_ _08119_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__mux2_1
Xhold1382 csr.mscratch\[16\] VGND VGND VPWR VPWR net1609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1393 _08171_ VGND VGND VPWR VPWR net1620 sky130_fd_sc_hd__dlygate4sd3_1
X_27686_ clknet_leaf_28_clock _00715_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24898_ csr._mcycle_T_3\[33\] csr._mcycle_T_3\[32\] csr.mcycle\[31\] _08646_ VGND
+ VGND VPWR VPWR _08647_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29425_ clknet_leaf_261_clock _02438_ VGND VGND VPWR VPWR decode.regfile.registers_5\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14651_ decode.id_ex_pc_reg\[12\] VGND VGND VPWR VPWR _10694_ sky130_fd_sc_hd__clkbuf_4
X_26637_ _09389_ _09676_ VGND VGND VPWR VPWR _09677_ sky130_fd_sc_hd__nand2_1
X_23849_ execute.io_target_pc\[18\] VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__buf_2
XFILLER_0_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13602_ net1751 _09938_ _09965_ _09957_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__o211a_1
X_29356_ clknet_leaf_227_clock _02369_ VGND VGND VPWR VPWR decode.regfile.registers_3\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_17370_ _11018_ _12977_ _12649_ decode.regfile.registers_10\[14\] _12652_ VGND VGND
+ VPWR VPWR _13321_ sky130_fd_sc_hd__o32a_1
X_26568_ net2387 _09636_ _09637_ _09635_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14582_ _10624_ VGND VGND VPWR VPWR _10625_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28307_ clknet_leaf_223_clock _01320_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16321_ decode.regfile.registers_14\[26\] _12018_ _12290_ _12291_ VGND VGND VPWR
+ VPWR _12292_ sky130_fd_sc_hd__a22o_1
X_13533_ _09879_ _09882_ fetch.bht.bhtTable_tag_MPORT_en _09892_ VGND VGND VPWR VPWR
+ _09909_ sky130_fd_sc_hd__and4b_1
X_25519_ net2668 _09008_ _09018_ _09017_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29287_ clknet_leaf_230_clock _02300_ VGND VGND VPWR VPWR decode.regfile.registers_1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_188_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26499_ net2188 _09592_ _09597_ _09595_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_188_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19040_ _04081_ _04091_ _03989_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__mux2_1
X_28238_ clknet_leaf_73_clock _01260_ VGND VGND VPWR VPWR csr._minstret_T_3\[38\]
+ sky130_fd_sc_hd__dfxtp_2
X_16252_ _11106_ _12223_ _12224_ VGND VGND VPWR VPWR _12225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15203_ _11194_ decode.regfile.registers_12\[0\] decode.regfile.registers_13\[0\]
+ _11196_ _11199_ VGND VGND VPWR VPWR _11200_ sky130_fd_sc_hd__o221a_1
XFILLER_0_168_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28169_ clknet_leaf_53_clock _01191_ VGND VGND VPWR VPWR csr.io_mret_vector\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16183_ decode.regfile.registers_18\[22\] _11455_ _11456_ VGND VGND VPWR VPWR _12158_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15134_ _11130_ VGND VGND VPWR VPWR _11131_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_226_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1090 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19942_ _03581_ _05201_ net2016 VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__and3b_1
X_15065_ _11061_ VGND VGND VPWR VPWR _11062_ sky130_fd_sc_hd__buf_4
XFILLER_0_26_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_222_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14016_ net2232 _10258_ _10267_ _10262_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19873_ _05142_ _03781_ _04225_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18824_ _03659_ execute.csr_read_data_out_reg\[8\] execute.io_reg_pc\[8\] _03777_
+ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__o22a_1
XFILLER_0_207_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18755_ _04034_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_106_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ decode.regfile.registers_21\[17\] _11222_ VGND VGND VPWR VPWR _11947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17706_ _13451_ net741 _13492_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14918_ _10947_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_1003 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18686_ _03714_ _03724_ decode.id_ex_rs2_data_reg\[0\] _03744_ VGND VGND VPWR VPWR
+ _03985_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_188_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15898_ _11191_ _11097_ decode.regfile.registers_5\[15\] VGND VGND VPWR VPWR _11880_
+ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_177_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17637_ _12649_ _12615_ _12880_ decode.regfile.registers_6\[21\] _03042_ VGND VGND
+ VPWR VPWR _03043_ sky130_fd_sc_hd__o221ai_4
X_14849_ _10678_ net337 _10891_ VGND VGND VPWR VPWR _10892_ sky130_fd_sc_hd__nor3_1
XFILLER_0_114_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17568_ decode.regfile.registers_18\[19\] _10925_ _12569_ _11023_ _11008_ VGND VGND
+ VPWR VPWR _02976_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_50_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19307_ _04410_ _04534_ _04598_ _04290_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16519_ _10961_ _11252_ _11944_ net500 _12484_ VGND VGND VPWR VPWR _12485_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17499_ _13091_ _13176_ decode.regfile.registers_27\[17\] _13050_ VGND VGND VPWR
+ VPWR _13447_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19238_ _04297_ _04261_ _04263_ _04284_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__a211o_1
XFILLER_0_171_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19169_ _04308_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21200_ _06095_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22180_ fetch.bht.bhtTable_tag\[0\]\[25\] fetch.bht.bhtTable_tag\[1\]\[25\] _06646_
+ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21131_ _09955_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_197_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21062_ _06017_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20013_ _05236_ _05237_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__nand2_1
X_25870_ _08943_ _09210_ VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_226_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24821_ _08113_ net2374 _08596_ VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27540_ clknet_5_7__leaf_clock _00569_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_2
X_24752_ _08560_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21964_ net2019 _06574_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23703_ net1240 _10807_ _07992_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__mux2_1
X_20915_ _05937_ _05933_ net42 VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__and3_1
X_24683_ net1868 execute.io_target_pc\[30\] _07285_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__mux2_1
X_27471_ clknet_leaf_52_clock _00500_ VGND VGND VPWR VPWR csr.io_csr_address\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_21895_ _06535_ _06519_ _06520_ _06536_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29210_ clknet_leaf_134_clock _02223_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23634_ net906 _10817_ _07961_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__mux2_1
X_26422_ _09417_ VGND VGND VPWR VPWR _09553_ sky130_fd_sc_hd__clkbuf_4
X_20846_ net109 _05891_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29141_ clknet_leaf_91_clock net1912 VGND VGND VPWR VPWR csr.mcycle\[25\] sky130_fd_sc_hd__dfxtp_2
X_23565_ net2289 _07918_ _07915_ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__or3b_1
XFILLER_0_147_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26353_ _09408_ _09502_ VGND VGND VPWR VPWR _09513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20777_ net100 net133 VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22516_ _07070_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__clkbuf_4
X_25304_ _08880_ decode.regfile.registers_0\[13\] VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29072_ clknet_leaf_208_clock _02085_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_26284_ net2537 _09462_ _09473_ _09471_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23496_ decode.id_ex_memread_reg VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28023_ clknet_leaf_214_clock _01045_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_25235_ _08074_ net1632 _08837_ VGND VGND VPWR VPWR _08847_ sky130_fd_sc_hd__mux2_1
X_22447_ _06674_ fetch.btb.btbTable\[6\]\[1\] fetch.bht.bhtTable_valid\[6\] VGND VGND
+ VPWR VPWR _07042_ sky130_fd_sc_hd__and3b_1
XFILLER_0_17_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25166_ net414 _08811_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22378_ fetch.bht.bhtTable_tag\[8\]\[16\] fetch.bht.bhtTable_tag\[9\]\[16\] fetch.bht.bhtTable_tag\[10\]\[16\]
+ fetch.bht.bhtTable_tag\[11\]\[16\] _06691_ _06677_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24117_ net853 VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21329_ net1162 _10787_ _06168_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__mux2_1
X_25097_ _08776_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28925_ clknet_leaf_178_clock _01938_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24048_ net826 execute.io_target_pc\[12\] _08187_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__mux2_1
Xhold490 decode.regfile.registers_3\[31\] VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28856_ clknet_leaf_124_clock _01869_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_16870_ _12830_ _12831_ VGND VGND VPWR VPWR _12832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15821_ _11153_ decode.regfile.registers_0\[13\] VGND VGND VPWR VPWR _11805_ sky130_fd_sc_hd__nand2_1
X_27807_ clknet_leaf_327_clock _00836_ VGND VGND VPWR VPWR memory.io_wb_readdata\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28787_ clknet_leaf_140_clock _01800_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25999_ _08920_ _09287_ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_216_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18540_ _03835_ _03838_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__or2_1
X_15752_ decode.regfile.registers_8\[11\] _11044_ _11174_ VGND VGND VPWR VPWR _11738_
+ sky130_fd_sc_hd__a21o_1
X_27738_ clknet_leaf_34_clock _00767_ VGND VGND VPWR VPWR decode.io_wb_rd\[1\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_137_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1190 csr.mscratch\[17\] VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__dlygate4sd3_1
X_14703_ _10711_ execute.io_target_pc\[2\] _10743_ execute.io_target_pc\[28\] VGND
+ VGND VPWR VPWR _10746_ sky130_fd_sc_hd__a22o_1
X_18471_ decode.id_ex_ex_rs1_reg\[3\] _03640_ _03650_ _03653_ _03651_ VGND VGND VPWR
+ VPWR _03770_ sky130_fd_sc_hd__o2111ai_4
X_15683_ decode.regfile.registers_21\[9\] _11648_ _11649_ _11670_ _11227_ VGND VGND
+ VPWR VPWR _11671_ sky130_fd_sc_hd__o221a_1
X_27669_ clknet_leaf_27_clock _00698_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17422_ _13183_ _13369_ _13370_ _13371_ VGND VGND VPWR VPWR _13372_ sky130_fd_sc_hd__a31o_1
X_29408_ clknet_leaf_247_clock _02421_ VGND VGND VPWR VPWR decode.regfile.registers_5\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14634_ decode.id_ex_pc_reg\[22\] VGND VGND VPWR VPWR _10677_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_215_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_215_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_215_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29339_ clknet_leaf_256_clock _02352_ VGND VGND VPWR VPWR decode.regfile.registers_3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_17353_ _11025_ _12690_ _12535_ VGND VGND VPWR VPWR _13304_ sky130_fd_sc_hd__and3_1
XFILLER_0_200_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14565_ _10607_ VGND VGND VPWR VPWR _10608_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16304_ decode.regfile.registers_17\[26\] _10988_ _11113_ _11118_ VGND VGND VPWR
+ VPWR _12275_ sky130_fd_sc_hd__and4_1
X_13516_ _09879_ _09882_ fetch.bht.bhtTable_tag_MPORT_en _09894_ VGND VGND VPWR VPWR
+ _09895_ sky130_fd_sc_hd__and4b_1
XFILLER_0_125_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17284_ _13225_ _13235_ _13236_ VGND VGND VPWR VPWR _13237_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14496_ _10136_ _10505_ VGND VGND VPWR VPWR _10544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19023_ _04321_ _04255_ _04248_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16235_ decode.regfile.registers_3\[24\] _11614_ _11367_ _11178_ VGND VGND VPWR VPWR
+ _12208_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_181_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16166_ _10659_ _10654_ net345 decode.regfile.registers_2\[22\] _11296_ VGND VGND
+ VPWR VPWR _12141_ sky130_fd_sc_hd__o32a_1
XFILLER_0_140_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15117_ _11113_ VGND VGND VPWR VPWR _11114_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_71_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16097_ _10649_ _10638_ _11052_ _10625_ VGND VGND VPWR VPWR _12074_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15048_ _11044_ VGND VGND VPWR VPWR _11045_ sky130_fd_sc_hd__buf_4
X_19925_ _04442_ _03766_ _03854_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19856_ _05126_ _03830_ _04219_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18807_ _03890_ decode.id_ex_imm_reg\[13\] _04101_ _04102_ _04105_ VGND VGND VPWR
+ VPWR _04106_ sky130_fd_sc_hd__a221o_2
X_19787_ _03835_ _03844_ _04234_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16999_ _10928_ decode.regfile.registers_26\[5\] _12814_ _11011_ _11027_ VGND VGND
+ VPWR VPWR _12959_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_69_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18738_ _09983_ net290 net273 VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__and3_1
XFILLER_0_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18669_ net330 _03645_ _03641_ _03643_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__and4_1
XFILLER_0_149_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20700_ _05801_ _05808_ decode.id_ex_rs1_data_reg\[10\] _05817_ _00697_ VGND VGND
+ VPWR VPWR _00729_ sky130_fd_sc_hd__a32o_1
X_21680_ csr.minstret\[21\] csr.minstret\[22\] _06381_ VGND VGND VPWR VPWR _06387_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20631_ _05761_ _05764_ _05630_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_28_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23350_ fetch.bht.bhtTable_target_pc\[12\]\[27\] fetch.bht.bhtTable_target_pc\[13\]\[27\]
+ fetch.bht.bhtTable_target_pc\[14\]\[27\] fetch.bht.bhtTable_target_pc\[15\]\[27\]
+ _07708_ _07103_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_178_Right_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20562_ net1417 _05592_ _05625_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__or3_1
XFILLER_0_190_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22301_ net226 _06877_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23281_ fetch.bht.bhtTable_target_pc\[0\]\[22\] fetch.bht.bhtTable_target_pc\[1\]\[22\]
+ fetch.bht.bhtTable_target_pc\[2\]\[22\] fetch.bht.bhtTable_target_pc\[3\]\[22\]
+ _07708_ _07710_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20493_ csr.mcycle\[8\] _05588_ _05575_ csr.minstret\[8\] VGND VGND VPWR VPWR _05645_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_229_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25020_ net2643 _08725_ VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22232_ fetch.bht.bhtTable_tag\[12\]\[15\] fetch.bht.bhtTable_tag\[13\]\[15\] _06700_
+ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22163_ fetch.bht.bhtTable_tag\[6\]\[13\] fetch.bht.bhtTable_tag\[7\]\[13\] _06644_
+ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21114_ _05949_ _06046_ net1058 VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22094_ _06673_ _06676_ _06682_ _06688_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__o22a_1
X_26971_ _10096_ _09862_ VGND VGND VPWR VPWR _09869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28710_ clknet_leaf_95_clock _01723_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout222 net82 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_4
X_25922_ net2384 _09242_ _09251_ _09250_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__o211a_1
X_21045_ execute.csr_read_data_out_reg\[12\] _06002_ _05998_ VGND VGND VPWR VPWR _06008_
+ sky130_fd_sc_hd__and3_1
X_29690_ clknet_leaf_289_clock _02703_ VGND VGND VPWR VPWR decode.regfile.registers_14\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28641_ clknet_leaf_174_clock _01654_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25853_ _08925_ _09210_ VGND VGND VPWR VPWR _09212_ sky130_fd_sc_hd__nand2_1
X_24804_ _08097_ net1735 _08585_ VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__mux2_1
X_28572_ clknet_leaf_191_clock _01585_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_25784_ net751 _09170_ _09172_ _09169_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__o211a_1
X_22996_ _07440_ _07441_ _07112_ _07442_ _07076_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_69_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27523_ clknet_leaf_44_clock _00552_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_4
X_24735_ _08097_ net1523 _08542_ VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21947_ _06573_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_179_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27454_ clknet_leaf_150_clock _00483_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24666_ _08516_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__clkbuf_1
X_21878_ csr.io_mret_vector\[12\] csr.io_mem_pc\[12\] _06515_ VGND VGND VPWR VPWR
+ _06525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26405_ _09385_ _09535_ VGND VGND VPWR VPWR _09543_ sky130_fd_sc_hd__nand2_1
X_23617_ _06147_ net1075 _07952_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__mux2_1
X_20829_ _05890_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27385_ clknet_leaf_10_clock _00414_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24597_ net1702 execute.io_target_pc\[20\] _08473_ VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29124_ clknet_leaf_73_clock _02137_ VGND VGND VPWR VPWR csr.mcycle\[8\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26336_ net1045 _09491_ _09503_ _09499_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__o211a_1
X_14350_ _10147_ _10418_ VGND VGND VPWR VPWR _10460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23548_ _10670_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_210_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_210_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29055_ clknet_leaf_180_clock _02068_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14281_ net532 _10419_ _10421_ _10411_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_324_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_324_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_163_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23479_ decode.control.io_funct7\[0\] _07876_ _07873_ VGND VGND VPWR VPWR _07878_
+ sky130_fd_sc_hd__or3b_1
X_26267_ _09398_ _09459_ VGND VGND VPWR VPWR _09464_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28006_ clknet_leaf_187_clock _01028_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16020_ decode.regfile.registers_9\[18\] _11365_ _11988_ _11997_ _11998_ VGND VGND
+ VPWR VPWR _11999_ sky130_fd_sc_hd__o221a_2
X_25218_ _08838_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26198_ net2665 _09395_ _09416_ _09418_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25149_ net420 _08802_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_339_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_339_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17971_ _12968_ _03366_ _03367_ _03368_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_208_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19710_ _04600_ _04359_ _04439_ _04986_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__a31o_1
X_28908_ clknet_leaf_108_clock _01921_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16922_ _12531_ _10592_ _12558_ decode.regfile.registers_0\[4\] VGND VGND VPWR VPWR
+ _12883_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29888_ clknet_leaf_305_clock _02901_ VGND VGND VPWR VPWR decode.regfile.registers_20\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19641_ _04541_ _04814_ _04920_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__o21a_1
XFILLER_0_217_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28839_ clknet_leaf_113_clock _01852_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16853_ _12695_ _12810_ _12813_ _12815_ VGND VGND VPWR VPWR _12816_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15804_ decode.regfile.registers_21\[12\] _11062_ _11100_ _11229_ _11788_ VGND VGND
+ VPWR VPWR _11789_ sky130_fd_sc_hd__o311a_1
X_19572_ _04442_ _03705_ _04306_ _03636_ _03593_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__o311a_1
XFILLER_0_176_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16784_ decode.regfile.registers_13\[1\] _12533_ _12582_ _12662_ VGND VGND VPWR VPWR
+ _12748_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13996_ net489 _10243_ _10256_ _10249_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_217_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18523_ _03797_ _03819_ _03708_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15735_ _11344_ net514 _11685_ _11721_ _11249_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_1126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18454_ execute.io_mem_rd\[4\] csr.io_csr_address\[4\] VGND VGND VPWR VPWR _03753_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15666_ _10659_ _10654_ net344 decode.regfile.registers_2\[9\] _11296_ VGND VGND
+ VPWR VPWR _11654_ sky130_fd_sc_hd__o32a_1
XFILLER_0_157_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17405_ _12499_ _12489_ _12511_ decode.regfile.registers_12\[15\] _12745_ VGND VGND
+ VPWR VPWR _13355_ sky130_fd_sc_hd__o32a_1
XFILLER_0_96_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14617_ _10659_ VGND VGND VPWR VPWR _10660_ sky130_fd_sc_hd__buf_6
XFILLER_0_28_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18385_ _03652_ decode.io_wb_rd\[4\] VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__nand2_1
Xclkbuf_5_13__f_clock clknet_2_1_0_clock VGND VGND VPWR VPWR clknet_5_13__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_15597_ _11576_ _11585_ _11586_ VGND VGND VPWR VPWR _11587_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17336_ _13263_ _13286_ _13164_ _13287_ VGND VGND VPWR VPWR _13288_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14548_ decode.immGen._imm_T_24\[19\] VGND VGND VPWR VPWR _10591_ sky130_fd_sc_hd__clkinv_4
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17267_ _13055_ decode.regfile.registers_30\[12\] _13097_ VGND VGND VPWR VPWR _13220_
+ sky130_fd_sc_hd__o21a_1
X_14479_ net822 _10533_ _10534_ _10535_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19006_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16218_ _11106_ _12190_ _12191_ VGND VGND VPWR VPWR _12192_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_1181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17198_ _12497_ _12503_ _12637_ decode.regfile.registers_11\[10\] VGND VGND VPWR
+ VPWR _13153_ sky130_fd_sc_hd__or4b_1
XFILLER_0_70_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16149_ decode.regfile.registers_21\[21\] _11061_ _11100_ _11229_ _12124_ VGND VGND
+ VPWR VPWR _12125_ sky130_fd_sc_hd__o311a_1
XFILLER_0_87_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19908_ _05168_ _05175_ _05176_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_127_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1904 decode.regfile.registers_13\[13\] VGND VGND VPWR VPWR net2131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1915 csr._mcycle_T_2\[24\] VGND VGND VPWR VPWR net2142 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19839_ _04509_ _04905_ _04511_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__and3_1
Xhold1926 decode.regfile.registers_19\[4\] VGND VGND VPWR VPWR net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1937 fetch.bht.bhtTable_tag\[13\]\[4\] VGND VGND VPWR VPWR net2164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1948 fetch.bht.bhtTable_target_pc\[6\]\[19\] VGND VGND VPWR VPWR net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1959 decode.regfile.registers_14\[17\] VGND VGND VPWR VPWR net2186 sky130_fd_sc_hd__dlygate4sd3_1
X_22850_ net1171 csr.io_mem_pc\[12\] _09898_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21801_ csr.io_csr_write_address\[5\] csr.io_csr_write_address\[4\] csr.io_csr_write_address\[7\]
+ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__nor3_1
XFILLER_0_79_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_870 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22781_ _09880_ _09882_ _09885_ _09892_ VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__and4_4
XFILLER_0_151_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24520_ _08441_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__clkbuf_1
X_21732_ _06427_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24451_ _08078_ net1840 _08400_ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__mux2_1
X_21663_ csr._mcycle_T_2\[18\] _06329_ csr.minstret\[18\] VGND VGND VPWR VPWR _06374_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23402_ _07821_ _07822_ _07823_ _07824_ _07080_ _06637_ VGND VGND VPWR VPWR _07825_
+ sky130_fd_sc_hd__mux4_2
X_20614_ csr._minstret_T_3\[56\] _05616_ _05618_ csr._csr_read_data_T_8\[24\] _05749_
+ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24382_ net997 VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__clkbuf_1
X_27170_ clknet_leaf_362_clock _00199_ VGND VGND VPWR VPWR decode.regfile.registers_27\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_21594_ _06322_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23333_ _06248_ _10915_ _07746_ _07760_ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26121_ net1502 _09356_ _09365_ _09359_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__o211a_1
X_20545_ _05685_ _05690_ _05630_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__o21a_2
XFILLER_0_7_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_104_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23264_ _07695_ _07114_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26052_ net2729 _09287_ _09325_ _09318_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__o211a_1
X_20476_ _05624_ _05629_ _05630_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22215_ fetch.bht.bhtTable_tag\[12\]\[20\] fetch.bht.bhtTable_tag\[13\]\[20\] fetch.bht.bhtTable_tag\[14\]\[20\]
+ fetch.bht.bhtTable_tag\[15\]\[20\] _06809_ _06649_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__mux4_1
X_25003_ net1370 csr.mcycle\[5\] _08701_ _08715_ _05856_ VGND VGND VPWR VPWR _02134_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_30_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23195_ execute.io_target_pc\[17\] _07091_ _06032_ _07630_ VGND VGND VPWR VPWR _07631_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29811_ clknet_leaf_296_clock _02824_ VGND VGND VPWR VPWR decode.regfile.registers_17\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22146_ fetch.bht.bhtTable_tag\[0\]\[23\] fetch.bht.bhtTable_tag\[1\]\[23\] fetch.bht.bhtTable_tag\[2\]\[23\]
+ fetch.bht.bhtTable_tag\[3\]\[23\] _06618_ _06652_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__mux4_1
XFILLER_0_219_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29742_ clknet_leaf_285_clock _02755_ VGND VGND VPWR VPWR decode.regfile.registers_15\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_22077_ _00002_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__buf_4
X_26954_ _10057_ _09849_ VGND VGND VPWR VPWR _09859_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25905_ _09240_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__clkbuf_4
X_21028_ execute.csr_read_data_out_reg\[4\] _05989_ _05998_ VGND VGND VPWR VPWR _05999_
+ sky130_fd_sc_hd__and3_1
X_29673_ clknet_leaf_277_clock _02686_ VGND VGND VPWR VPWR decode.regfile.registers_13\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_26885_ _09794_ VGND VGND VPWR VPWR _09819_ sky130_fd_sc_hd__buf_2
XFILLER_0_214_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_113_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28624_ clknet_leaf_120_clock _01637_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13850_ net647 _10167_ _10170_ _10162_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__o211a_1
X_25836_ net1169 _09199_ _09202_ _09194_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_214_Right_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28555_ clknet_leaf_234_clock _01568_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13781_ _10060_ memory.io_wb_aluresult\[27\] _10004_ memory.io_wb_readdata\[27\]
+ VGND VGND VPWR VPWR _10119_ sky130_fd_sc_hd__a22o_1
X_25767_ net1126 _09156_ _09162_ _09153_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__o211a_1
X_22979_ net94 net93 _07393_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15520_ _11193_ decode.regfile.registers_12\[5\] decode.regfile.registers_13\[5\]
+ _11195_ _11198_ VGND VGND VPWR VPWR _11512_ sky130_fd_sc_hd__o221a_1
X_27506_ clknet_leaf_14_clock _00535_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dfxtp_1
X_24718_ _08543_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__clkbuf_1
X_28486_ clknet_leaf_211_clock _01499_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25698_ _09110_ VGND VGND VPWR VPWR _09122_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_191_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27437_ clknet_leaf_146_clock _00466_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15451_ _10962_ decode.regfile.registers_30\[4\] _11039_ _11032_ _11033_ VGND VGND
+ VPWR VPWR _11444_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24649_ net1203 VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14402_ _10087_ _10487_ VGND VGND VPWR VPWR _10491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18170_ _03463_ _03464_ _10921_ decode.control.io_funct7\[4\] VGND VGND VPWR VPWR
+ _03513_ sky130_fd_sc_hd__and4bb_1
Xclkbuf_leaf_263_clock clknet_5_22__leaf_clock VGND VGND VPWR VPWR clknet_leaf_263_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_182_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27368_ clknet_leaf_33_clock _00397_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15382_ _11376_ decode.regfile.registers_5\[2\] _11291_ VGND VGND VPWR VPWR _11377_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_122_Left_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17121_ decode.regfile.registers_20\[8\] _12771_ _13076_ _13077_ _12538_ VGND VGND
+ VPWR VPWR _13078_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29107_ clknet_leaf_17_clock _02120_ VGND VGND VPWR VPWR csr._mcycle_T_3\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14333_ _10102_ _10444_ VGND VGND VPWR VPWR _10451_ sky130_fd_sc_hd__nand2_1
X_26319_ _09450_ _09492_ VGND VGND VPWR VPWR _09494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27299_ clknet_leaf_13_clock _00328_ VGND VGND VPWR VPWR decode.regfile.registers_31\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29038_ clknet_leaf_109_clock _02051_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052_ _11023_ _12552_ _12523_ _12561_ decode.regfile.registers_19\[7\] VGND VGND
+ VPWR VPWR _13010_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_150_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14264_ _10290_ VGND VGND VPWR VPWR _10411_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap208 _03714_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_4
XFILLER_0_151_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap219 _04391_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
X_16003_ _11761_ net411 _11943_ _11982_ _11760_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_278_clock clknet_5_21__leaf_clock VGND VGND VPWR VPWR clknet_leaf_278_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_180_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14195_ net2723 _10359_ _10370_ _10369_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_201_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_201_clock
+ sky130_fd_sc_hd__clkbuf_8
X_17954_ decode.regfile.registers_9\[29\] _12607_ _03350_ _03351_ _12600_ VGND VGND
+ VPWR VPWR _03352_ sky130_fd_sc_hd__a221oi_2
XPHY_EDGE_ROW_131_Left_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16905_ _12695_ _12864_ _12865_ _12866_ VGND VGND VPWR VPWR _12867_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17885_ decode.regfile.registers_16\[27\] _12575_ _03266_ _03284_ _12578_ VGND VGND
+ VPWR VPWR _03285_ sky130_fd_sc_hd__o221a_1
XFILLER_0_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19624_ _04893_ _04895_ _04903_ _04904_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__o31a_1
X_16836_ decode.regfile.registers_15\[2\] _12585_ _12674_ _12798_ VGND VGND VPWR VPWR
+ _12799_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_7_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_7_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_122_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_216_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_216_clock
+ sky130_fd_sc_hd__clkbuf_8
X_19555_ _04180_ net254 _04181_ _04182_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16767_ decode.immGen._imm_T_24\[19\] _10597_ _10607_ _10934_ VGND VGND VPWR VPWR
+ _12731_ sky130_fd_sc_hd__or4_1
X_13979_ _10244_ net211 VGND VGND VPWR VPWR _10247_ sky130_fd_sc_hd__nand2_1
XFILLER_0_221_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18506_ execute.io_mem_memtoreg\[1\] execute.io_mem_memtoreg\[0\] execute.io_reg_pc\[26\]
+ _03804_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__o31a_1
XFILLER_0_158_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15718_ decode.regfile.registers_12\[10\] _10640_ _11690_ _11691_ _11704_ VGND VGND
+ VPWR VPWR _11705_ sky130_fd_sc_hd__o32a_1
X_19486_ _04409_ _04770_ _04771_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16698_ _12662_ VGND VGND VPWR VPWR _12663_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_83_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18437_ decode.io_wb_rd\[1\] _03710_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__or2b_4
XFILLER_0_186_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15649_ decode.regfile.registers_21\[8\] _11061_ _11100_ _11229_ _11637_ VGND VGND
+ VPWR VPWR _11638_ sky130_fd_sc_hd__o311a_1
XFILLER_0_173_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_140_Left_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18368_ execute.csr_read_data_out_reg\[31\] _03659_ net124 _03666_ VGND VGND VPWR
+ VPWR _03667_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17319_ _12830_ _13269_ _12835_ _13270_ VGND VGND VPWR VPWR _13271_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18299_ _03614_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_116_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20330_ _10790_ _05494_ decode.id_ex_pc_reg\[26\] VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_116_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20261_ _05445_ _05446_ _05418_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22000_ _06578_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20192_ decode.id_ex_imm_reg\[26\] decode.id_ex_pc_reg\[26\] VGND VGND VPWR VPWR
+ _05391_ sky130_fd_sc_hd__nand2_1
Xhold2402 decode.regfile.registers_18\[25\] VGND VGND VPWR VPWR net2629 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2413 decode.regfile.registers_30\[6\] VGND VGND VPWR VPWR net2640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2424 decode.regfile.registers_26\[25\] VGND VGND VPWR VPWR net2651 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2435 csr._csr_read_data_T_8\[2\] VGND VGND VPWR VPWR net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1701 fetch.bht.bhtTable_target_pc\[15\]\[14\] VGND VGND VPWR VPWR net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2446 csr._minstret_T_3\[36\] VGND VGND VPWR VPWR net2673 sky130_fd_sc_hd__dlygate4sd3_1
X_23951_ net1017 _08109_ _06156_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__mux2_1
Xhold2457 csr._csr_read_data_T_8\[26\] VGND VGND VPWR VPWR net2684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1712 decode.regfile.registers_28\[15\] VGND VGND VPWR VPWR net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1723 csr.mscratch\[18\] VGND VGND VPWR VPWR net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2468 decode.regfile.registers_0\[25\] VGND VGND VPWR VPWR net2695 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1734 decode.regfile.registers_3\[30\] VGND VGND VPWR VPWR net1961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2479 decode.regfile.registers_5\[25\] VGND VGND VPWR VPWR net2706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1745 fetch.bht.bhtTable_tag\[7\]\[22\] VGND VGND VPWR VPWR net1972 sky130_fd_sc_hd__dlygate4sd3_1
X_22902_ _06785_ _07349_ _07352_ _07035_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__or4b_1
Xhold1756 decode.id_ex_isjump_reg VGND VGND VPWR VPWR net1983 sky130_fd_sc_hd__dlygate4sd3_1
X_26670_ net2477 _09692_ _09695_ _09688_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__o211a_1
X_23882_ execute.io_target_pc\[29\] VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__buf_2
Xhold1767 decode.regfile.registers_15\[20\] VGND VGND VPWR VPWR net1994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1778 fetch.bht.bhtTable_target_pc\[0\]\[7\] VGND VGND VPWR VPWR net2005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1789 decode.id_ex_memwrite_reg VGND VGND VPWR VPWR net2016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25621_ _08920_ _09069_ VGND VGND VPWR VPWR _09078_ sky130_fd_sc_hd__nand2_1
X_22833_ _07312_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28340_ clknet_leaf_215_clock _01353_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_25552_ net673 _09024_ _09038_ _09033_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_49_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22764_ _06138_ net1869 _07265_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24503_ _08432_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21715_ csr.minstret\[27\] csr.minstret\[28\] _06404_ VGND VGND VPWR VPWR _06415_
+ sky130_fd_sc_hd__and3_1
X_28271_ clknet_leaf_61_clock _01293_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_22695_ _07209_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__buf_2
X_25483_ net926 _08995_ _08998_ _08991_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27222_ clknet_leaf_7_clock _00251_ VGND VGND VPWR VPWR decode.regfile.registers_29\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_24434_ _08062_ net1589 _08389_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21646_ csr.minstret\[10\] csr.minstret\[11\] _06349_ _06360_ VGND VGND VPWR VPWR
+ _06361_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27153_ clknet_leaf_353_clock _00182_ VGND VGND VPWR VPWR decode.regfile.registers_27\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_21577_ _06309_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__clkbuf_1
X_24365_ _08359_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_60 _10795_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_71 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_82 _12221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26104_ _09328_ VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__clkbuf_4
X_23316_ _07619_ _07573_ _07620_ _07744_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__a31o_1
X_20528_ _05526_ _05536_ _05617_ csr._csr_read_data_T_8\[12\] _05675_ VGND VGND VPWR
+ VPWR _05676_ sky130_fd_sc_hd__a221o_1
XANTENNA_93 decode.regfile.registers_12\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24296_ _08057_ net1830 _08323_ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__mux2_1
X_27084_ clknet_leaf_348_clock _00113_ VGND VGND VPWR VPWR decode.regfile.registers_24\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26035_ net2639 _09313_ _09316_ _09305_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__o211a_1
X_23247_ fetch.bht.bhtTable_target_pc\[12\]\[20\] fetch.bht.bhtTable_target_pc\[13\]\[20\]
+ fetch.bht.bhtTable_target_pc\[14\]\[20\] fetch.bht.bhtTable_target_pc\[15\]\[20\]
+ _07669_ _07100_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__mux4_1
X_20459_ _05613_ _05574_ _05586_ csr.mcycle\[4\] _05614_ VGND VGND VPWR VPWR _05615_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23178_ _07368_ _07614_ _05864_ _07345_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22129_ _06721_ _06690_ _06672_ _06723_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_140_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27986_ clknet_leaf_168_clock _01008_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29725_ clknet_leaf_312_clock _02738_ VGND VGND VPWR VPWR decode.regfile.registers_15\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_201_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ _10978_ VGND VGND VPWR VPWR _10979_ sky130_fd_sc_hd__clkbuf_4
X_26937_ _09838_ VGND VGND VPWR VPWR _09849_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_197_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ _09964_ _10200_ VGND VGND VPWR VPWR _10202_ sky130_fd_sc_hd__nand2_1
X_17670_ decode.regfile.registers_18\[22\] _12571_ _12561_ VGND VGND VPWR VPWR _03075_
+ sky130_fd_sc_hd__a21o_1
X_29656_ clknet_leaf_289_clock _02669_ VGND VGND VPWR VPWR decode.regfile.registers_12\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26868_ _09396_ _09806_ VGND VGND VPWR VPWR _09810_ sky130_fd_sc_hd__nand2_1
X_14882_ _10920_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28607_ clknet_leaf_180_clock _01620_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16621_ _12534_ VGND VGND VPWR VPWR _12586_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_193_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13833_ net2509 _10153_ _10160_ _10132_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__o211a_1
X_25819_ net2337 _09183_ _09191_ _09182_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29587_ clknet_leaf_274_clock _02600_ VGND VGND VPWR VPWR decode.regfile.registers_10\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_26799_ _09402_ _09763_ VGND VGND VPWR VPWR _09770_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19340_ _04617_ _04619_ _04622_ _04631_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__o211ai_2
X_28538_ clknet_leaf_195_clock _01551_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16552_ decode.regfile.registers_25\[0\] _12513_ _12516_ decode.regfile.registers_24\[0\]
+ VGND VGND VPWR VPWR _12517_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_97_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13764_ _10060_ memory.io_wb_aluresult\[24\] _10004_ memory.io_wb_readdata\[24\]
+ _10005_ VGND VGND VPWR VPWR _10105_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15503_ _10956_ decode.regfile.registers_22\[5\] _11093_ _10977_ _10989_ VGND VGND
+ VPWR VPWR _11495_ sky130_fd_sc_hd__o2111a_1
X_19271_ _04245_ _04303_ _04556_ _04564_ _04306_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__o311a_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28469_ clknet_leaf_139_clock _01482_ VGND VGND VPWR VPWR decode.io_id_pc\[27\] sky130_fd_sc_hd__dfxtp_1
X_16483_ _10961_ _11834_ _11944_ decode.regfile.registers_29\[30\] _12449_ VGND VGND
+ VPWR VPWR _12450_ sky130_fd_sc_hd__o221a_1
XFILLER_0_167_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13695_ _09989_ _10044_ _10045_ _10046_ VGND VGND VPWR VPWR _10047_ sky130_fd_sc_hd__a31o_4
XFILLER_0_167_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18222_ csr.mcycle\[0\] csr.mcycle\[2\] csr.mcycle\[1\] VGND VGND VPWR VPWR _03557_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_127_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15434_ _11269_ _11426_ _11427_ VGND VGND VPWR VPWR _11428_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_182_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18153_ _03495_ _10910_ _03500_ decode.io_id_pc\[31\] VGND VGND VPWR VPWR _03506_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15365_ _11207_ VGND VGND VPWR VPWR _11360_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_170_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17104_ decode.regfile.registers_3\[8\] _12836_ _10609_ _12614_ VGND VGND VPWR VPWR
+ _13061_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14316_ net547 _10434_ _10441_ _10440_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18084_ _10910_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15296_ _10627_ decode.immGen._imm_T_24\[11\] _11108_ _11056_ VGND VGND VPWR VPWR
+ _11292_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold308 decode.regfile.registers_29\[13\] VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 csr.mcycle\[31\] VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ decode.regfile.registers_22\[6\] _12527_ _12992_ _12993_ _12686_ VGND VGND
+ VPWR VPWR _12994_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14247_ net2496 _10390_ _10401_ _10398_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_229_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_140_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_140_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14178_ net2155 _10359_ _10361_ _10357_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_209_Left_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18986_ _03863_ _04254_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__or2_1
Xhold1008 fetch.bht.bhtTable_tag\[3\]\[5\] VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__dlygate4sd3_1
X_17937_ _12708_ net605 _03301_ _03335_ _03073_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__o221a_1
Xhold1019 decode.regfile.registers_6\[3\] VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_155_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_155_clock
+ sky130_fd_sc_hd__clkbuf_8
X_17868_ decode.regfile.registers_7\[27\] _12610_ _12622_ decode.regfile.registers_6\[27\]
+ _12843_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19607_ _04201_ _03938_ _04862_ _04863_ _03912_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_75_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16819_ decode.regfile.registers_3\[2\] _12629_ _12732_ VGND VGND VPWR VPWR _12782_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_177_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17799_ decode.regfile.registers_10\[25\] _12600_ _03199_ _03200_ VGND VGND VPWR
+ VPWR _03201_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_141_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19538_ _04818_ _04526_ _04452_ _04819_ _04821_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19469_ _04415_ _04737_ _04750_ _04755_ _04729_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__o311a_1
XFILLER_0_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_218_Left_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_250 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21500_ _06267_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_261 net2798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_272 _10594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22480_ _06633_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__buf_4
XFILLER_0_174_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_283 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_294 _12553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21431_ _06122_ net1594 _06230_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24150_ _08248_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21362_ _06193_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23101_ fetch.bht.bhtTable_target_pc\[8\]\[12\] fetch.bht.bhtTable_target_pc\[9\]\[12\]
+ fetch.bht.bhtTable_target_pc\[10\]\[12\] fetch.bht.bhtTable_target_pc\[11\]\[12\]
+ _07107_ _07114_ VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__mux4_1
X_20313_ _05340_ _10867_ _10798_ _05473_ _10864_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__a41o_1
X_24081_ net1029 execute.io_target_pc\[28\] _07991_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21293_ _09885_ _09890_ _09917_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__and3_4
XFILLER_0_141_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold820 decode.regfile.registers_20\[5\] VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold831 execute.csr_write_data_out_reg\[3\] VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 fetch.bht.bhtTable_target_pc\[3\]\[14\] VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__dlygate4sd3_1
X_23032_ _07108_ fetch.bht.bhtTable_target_pc\[10\]\[8\] VGND VGND VPWR VPWR _07477_
+ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_108_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_108_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold853 fetch.bht.bhtTable_target_pc\[8\]\[28\] VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__dlygate4sd3_1
X_20244_ _10704_ _10678_ _05427_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__and3_1
Xhold864 fetch.bht.bhtTable_target_pc\[15\]\[10\] VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_227_Left_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold875 decode.regfile.registers_17\[6\] VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 decode.regfile.registers_26\[12\] VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 fetch.bht.bhtTable_target_pc\[1\]\[25\] VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__dlygate4sd3_1
X_27840_ clknet_leaf_326_clock _00869_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_20175_ _05368_ _05372_ _05369_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_38_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2210 _01125_ VGND VGND VPWR VPWR net2437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2221 decode.regfile.registers_12\[26\] VGND VGND VPWR VPWR net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2232 decode.io_id_pc\[7\] VGND VGND VPWR VPWR net2459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2243 decode.regfile.registers_0\[1\] VGND VGND VPWR VPWR net2470 sky130_fd_sc_hd__dlygate4sd3_1
X_27771_ clknet_leaf_324_clock _00800_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24983_ net340 VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__clkbuf_4
Xhold2254 csr._minstret_T_3\[56\] VGND VGND VPWR VPWR net2481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1520 fetch.bht.bhtTable_target_pc\[0\]\[18\] VGND VGND VPWR VPWR net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2265 decode.regfile.registers_1\[30\] VGND VGND VPWR VPWR net2492 sky130_fd_sc_hd__dlygate4sd3_1
X_29510_ clknet_leaf_267_clock _02523_ VGND VGND VPWR VPWR decode.regfile.registers_8\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26722_ _09400_ _09720_ VGND VGND VPWR VPWR _09726_ sky130_fd_sc_hd__nand2_1
Xhold2276 decode.regfile.registers_22\[22\] VGND VGND VPWR VPWR net2503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 decode.regfile.registers_10\[17\] VGND VGND VPWR VPWR net1758 sky130_fd_sc_hd__dlygate4sd3_1
X_23934_ _08137_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__clkbuf_1
Xhold1542 fetch.bht.bhtTable_target_pc\[1\]\[1\] VGND VGND VPWR VPWR net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2287 fetch.btb.btbTable\[10\]\[1\] VGND VGND VPWR VPWR net2514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1553 fetch.bht.bhtTable_target_pc\[6\]\[31\] VGND VGND VPWR VPWR net1780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2298 decode.regfile.registers_8\[25\] VGND VGND VPWR VPWR net2525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1564 decode.regfile.registers_24\[13\] VGND VGND VPWR VPWR net1791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1575 decode.regfile.registers_15\[2\] VGND VGND VPWR VPWR net1802 sky130_fd_sc_hd__dlygate4sd3_1
X_29441_ clknet_leaf_248_clock _02454_ VGND VGND VPWR VPWR decode.regfile.registers_6\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1586 fetch.bht.bhtTable_tag\[11\]\[24\] VGND VGND VPWR VPWR net1813 sky130_fd_sc_hd__dlygate4sd3_1
X_26653_ net519 _09679_ _09685_ _09675_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__o211a_1
X_23865_ _08097_ net2050 _08079_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__mux2_1
Xhold1597 decode.regfile.registers_22\[16\] VGND VGND VPWR VPWR net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25604_ _09067_ VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__buf_2
X_22816_ _07303_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__clkbuf_1
X_29372_ clknet_leaf_256_clock _02385_ VGND VGND VPWR VPWR decode.regfile.registers_4\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_26584_ _09412_ _09645_ VGND VGND VPWR VPWR _09646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23796_ execute.io_target_pc\[1\] VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__buf_2
XFILLER_0_184_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28323_ clknet_leaf_186_clock _01336_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25535_ _08910_ _09026_ VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__nand2_1
X_22747_ _07266_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28254_ clknet_leaf_79_clock _01276_ VGND VGND VPWR VPWR csr._minstret_T_3\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_25466_ _08918_ _08980_ VGND VGND VPWR VPWR _08988_ sky130_fd_sc_hd__nand2_1
X_22678_ net2534 _07222_ _07226_ _07221_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__o211a_1
X_27205_ clknet_leaf_364_clock _00234_ VGND VGND VPWR VPWR decode.regfile.registers_28\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_24417_ net1166 execute.io_target_pc\[31\] _09911_ VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28185_ clknet_leaf_59_clock _01207_ VGND VGND VPWR VPWR csr.io_mret_vector\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_21629_ csr.minstret\[6\] csr.minstret\[7\] csr.minstret\[8\] csr.minstret\[9\] VGND
+ VGND VPWR VPWR _06349_ sky130_fd_sc_hd__and4_1
XFILLER_0_164_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25397_ _10063_ VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_124_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15150_ decode.immGen._imm_T_24\[1\] _11107_ _11041_ VGND VGND VPWR VPWR _11147_
+ sky130_fd_sc_hd__nand3_4
X_27136_ clknet_leaf_359_clock _00165_ VGND VGND VPWR VPWR decode.regfile.registers_26\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_24348_ _08350_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14101_ net2556 _10315_ _10316_ _10317_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27067_ clknet_leaf_349_clock _00096_ VGND VGND VPWR VPWR decode.regfile.registers_24\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15081_ _10960_ decode.regfile.registers_25\[0\] _11075_ _11077_ VGND VGND VPWR VPWR
+ _11078_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24279_ _08107_ net1438 _06218_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14032_ _10107_ _10268_ VGND VGND VPWR VPWR _10277_ sky130_fd_sc_hd__nand2_1
X_26018_ _08939_ _09297_ VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18840_ decode.id_ex_rs2_data_reg\[9\] net307 _03763_ _04133_ _04138_ VGND VGND VPWR
+ VPWR _04139_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_224_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_224_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_224_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_72_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_72_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18771_ _03656_ _04067_ _03670_ _04069_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__o211a_4
X_27969_ clknet_leaf_219_clock _00991_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15983_ _10649_ _10631_ _11052_ decode.regfile.registers_11\[17\] _11315_ VGND VGND
+ VPWR VPWR _11963_ sky130_fd_sc_hd__o32a_1
XFILLER_0_98_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ _11018_ _12977_ _12510_ decode.regfile.registers_8\[23\] _12892_ VGND VGND
+ VPWR VPWR _03126_ sky130_fd_sc_hd__o32a_1
X_14934_ _10948_ _10954_ _10962_ VGND VGND VPWR VPWR _10963_ sky130_fd_sc_hd__and3b_1
X_29708_ clknet_leaf_284_clock _02721_ VGND VGND VPWR VPWR decode.regfile.registers_14\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17653_ decode.regfile.registers_20\[21\] _12771_ _03057_ _03058_ _12538_ VGND VGND
+ VPWR VPWR _03059_ sky130_fd_sc_hd__a221o_1
X_14865_ fetch.bht.bhtTable_tag_MPORT_en _10907_ VGND VGND VPWR VPWR _10908_ sky130_fd_sc_hd__nor2_2
X_29639_ clknet_leaf_278_clock _02652_ VGND VGND VPWR VPWR decode.regfile.registers_12\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_87_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_87_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16604_ _12568_ VGND VGND VPWR VPWR _12569_ sky130_fd_sc_hd__buf_4
X_13816_ _09933_ VGND VGND VPWR VPWR _10149_ sky130_fd_sc_hd__clkbuf_4
X_17584_ _12697_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14796_ decode.id_ex_pc_reg\[4\] _10829_ _10838_ VGND VGND VPWR VPWR _10839_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19323_ _04227_ _04614_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16535_ _12499_ _10611_ VGND VGND VPWR VPWR _12500_ sky130_fd_sc_hd__nand2_4
XFILLER_0_156_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13747_ memory.csr_read_data_out_reg\[21\] _09987_ _10089_ _10090_ VGND VGND VPWR
+ VPWR _10091_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_175_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19254_ _04325_ net262 _04307_ _03670_ _04541_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__a41o_1
Xclkbuf_leaf_10_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_10_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16466_ decode.regfile.registers_13\[30\] _10639_ _11186_ _12431_ _12432_ VGND VGND
+ VPWR VPWR _12433_ sky130_fd_sc_hd__a32o_1
XFILLER_0_186_1320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13678_ net550 _10027_ _10032_ _10020_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18205_ _03541_ _10949_ _11000_ _03542_ _11006_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15417_ decode.regfile.registers_1\[3\] _11116_ _11137_ _11157_ VGND VGND VPWR VPWR
+ _11411_ sky130_fd_sc_hd__and4_1
XFILLER_0_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19185_ _03997_ _03998_ _04379_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_171_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16397_ _10988_ _11113_ _11119_ _12365_ VGND VGND VPWR VPWR _12366_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18136_ _03495_ _03493_ _03487_ net2190 VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15348_ _11251_ net539 _11253_ _11248_ _11343_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__o311a_1
XFILLER_0_85_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_25_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_184_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18067_ _03452_ _10916_ _03456_ _10018_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__and4b_1
XFILLER_0_223_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_184_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15279_ _10637_ _11143_ _11035_ VGND VGND VPWR VPWR _11275_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold149 io_fetch_data[1] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17018_ _12502_ VGND VGND VPWR VPWR _12977_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _04015_ _04016_ _04017_ _04019_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_143_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21980_ net881 _06587_ _06593_ _06592_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_33_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_17 _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_28 _05697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_39 _08948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20931_ _05946_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23650_ _07973_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__clkbuf_1
X_20862_ _05908_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_1092 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22601_ _07177_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_102_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23581_ _07935_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20793_ net2715 _05867_ _05868_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25320_ _08890_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22532_ _07124_ _07125_ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25251_ _08855_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__clkbuf_1
X_22463_ _06699_ _07050_ _07052_ _07057_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24202_ _08275_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21414_ _06105_ net2278 _06219_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22394_ _06673_ _06984_ _06641_ _06988_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__o211ai_1
X_25182_ _09883_ _08801_ _09881_ VGND VGND VPWR VPWR _08820_ sky130_fd_sc_hd__or3b_2
XFILLER_0_60_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24133_ net1352 execute.io_target_pc\[21\] _08232_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__mux2_1
X_21345_ _06183_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28941_ clknet_leaf_102_clock _01954_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_24064_ _08204_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__clkbuf_1
X_21276_ net921 _06143_ _06141_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__mux2_1
Xhold650 execute.csr_write_data_out_reg\[7\] VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold661 decode.regfile.registers_17\[5\] VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold672 fetch.bht.bhtTable_target_pc\[11\]\[22\] VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd3_1
X_23015_ fetch.bht.bhtTable_target_pc\[8\]\[7\] fetch.bht.bhtTable_target_pc\[9\]\[7\]
+ fetch.bht.bhtTable_target_pc\[10\]\[7\] fetch.bht.bhtTable_target_pc\[11\]\[7\]
+ _07108_ _07125_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__mux4_1
Xhold683 fetch.bht.bhtTable_tag\[11\]\[14\] VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__dlygate4sd3_1
X_20227_ _05416_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28872_ clknet_leaf_100_clock _01885_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold694 fetch.bht.bhtTable_tag\[8\]\[20\] VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27823_ clknet_leaf_317_clock _00852_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_20158_ _05358_ _05362_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_5_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2040 decode.regfile.registers_20\[21\] VGND VGND VPWR VPWR net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2051 fetch.bht.bhtTable_tag\[6\]\[2\] VGND VGND VPWR VPWR net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2062 decode.io_id_pc\[30\] VGND VGND VPWR VPWR net2289 sky130_fd_sc_hd__dlygate4sd3_1
X_27754_ clknet_leaf_321_clock _00783_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2073 decode.io_id_pc\[10\] VGND VGND VPWR VPWR net2300 sky130_fd_sc_hd__dlygate4sd3_1
X_20089_ _05295_ _05299_ _05301_ _05302_ _05296_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__o221ai_1
X_24966_ net949 _08689_ _08690_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__o21ba_1
Xhold2084 decode.regfile.registers_17\[26\] VGND VGND VPWR VPWR net2311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1350 decode.regfile.registers_24\[16\] VGND VGND VPWR VPWR net1577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2095 decode.regfile.registers_8\[18\] VGND VGND VPWR VPWR net2322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 fetch.bht.bhtTable_target_pc\[13\]\[1\] VGND VGND VPWR VPWR net1588 sky130_fd_sc_hd__dlygate4sd3_1
X_26705_ _09383_ _09710_ VGND VGND VPWR VPWR _09716_ sky130_fd_sc_hd__nand2_1
Xhold1372 fetch.bht.bhtTable_target_pc\[9\]\[4\] VGND VGND VPWR VPWR net1599 sky130_fd_sc_hd__dlygate4sd3_1
X_23917_ _08128_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__clkbuf_1
X_27685_ clknet_leaf_28_clock _00714_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1383 _01236_ VGND VGND VPWR VPWR net1610 sky130_fd_sc_hd__dlygate4sd3_1
X_24897_ _08639_ _08641_ _08645_ VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__and3_1
Xhold1394 fetch.bht.bhtTable_target_pc\[6\]\[11\] VGND VGND VPWR VPWR net1621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29424_ clknet_leaf_260_clock _02437_ VGND VGND VPWR VPWR decode.regfile.registers_5\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14650_ decode.id_ex_pc_reg\[24\] VGND VGND VPWR VPWR _10693_ sky130_fd_sc_hd__inv_2
X_26636_ _09664_ VGND VGND VPWR VPWR _09676_ sky130_fd_sc_hd__clkbuf_4
X_23848_ _08086_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13601_ _09964_ _09951_ VGND VGND VPWR VPWR _09965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29355_ clknet_leaf_228_clock _02368_ VGND VGND VPWR VPWR decode.regfile.registers_3\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26567_ _09396_ _09632_ VGND VGND VPWR VPWR _09637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14581_ _10623_ VGND VGND VPWR VPWR _10624_ sky130_fd_sc_hd__buf_4
X_23779_ _06140_ net1762 _08041_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28306_ clknet_leaf_215_clock _01319_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16320_ _11194_ decode.regfile.registers_12\[26\] decode.regfile.registers_13\[26\]
+ _11196_ _12074_ VGND VGND VPWR VPWR _12291_ sky130_fd_sc_hd__o221a_1
XFILLER_0_184_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13532_ _09908_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__clkbuf_1
X_25518_ _08968_ _08978_ VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29286_ clknet_leaf_243_clock _02299_ VGND VGND VPWR VPWR decode.regfile.registers_1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26498_ _09402_ _09589_ VGND VGND VPWR VPWR _09597_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_188_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_188_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28237_ clknet_leaf_73_clock net714 VGND VGND VPWR VPWR csr._minstret_T_3\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16251_ decode.regfile.registers_18\[24\] _10642_ _11112_ _10988_ _10976_ VGND VGND
+ VPWR VPWR _12224_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_36_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25449_ _09932_ _03672_ _08903_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__and3_1
XFILLER_0_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15202_ _11198_ VGND VGND VPWR VPWR _11199_ sky130_fd_sc_hd__clkbuf_4
X_28168_ clknet_leaf_53_clock _01190_ VGND VGND VPWR VPWR csr.io_mret_vector\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16182_ _11124_ _12155_ _12156_ VGND VGND VPWR VPWR _12157_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27119_ clknet_leaf_352_clock _00148_ VGND VGND VPWR VPWR decode.regfile.registers_26\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_15133_ _11129_ _10654_ _10623_ _10659_ VGND VGND VPWR VPWR _11130_ sky130_fd_sc_hd__or4b_1
XFILLER_0_105_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_226_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28099_ clknet_leaf_74_clock _01121_ VGND VGND VPWR VPWR csr.minstret\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1006 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15064_ _11060_ VGND VGND VPWR VPWR _11061_ sky130_fd_sc_hd__clkbuf_4
X_19941_ _05204_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14015_ _10069_ _10255_ VGND VGND VPWR VPWR _10267_ sky130_fd_sc_hd__nand2_1
X_19872_ _04297_ decode.id_ex_imm_reg\[29\] _03787_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18823_ _10014_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__inv_2
X_18754_ _03976_ _04026_ _04029_ _04039_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__o311ai_2
X_15966_ _11263_ decode.regfile.registers_22\[17\] _11404_ _11264_ _11265_ VGND VGND
+ VPWR VPWR _11946_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_106_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14917_ _10912_ _10913_ _10921_ _10946_ VGND VGND VPWR VPWR _10947_ sky130_fd_sc_hd__and4bb_1
X_17705_ _12708_ net436 _03074_ _03109_ _03073_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__o221a_1
XFILLER_0_222_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15897_ decode.regfile.registers_13\[15\] _11276_ VGND VGND VPWR VPWR _11879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18685_ net308 _03981_ decode.id_ex_immsrc_reg VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_188_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14848_ csr.io_mem_pc\[5\] net288 _10820_ VGND VGND VPWR VPWR _10891_ sky130_fd_sc_hd__a21oi_1
X_17636_ _12880_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17567_ decode.regfile.registers_17\[19\] _12580_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14779_ _10820_ _10815_ _10821_ VGND VGND VPWR VPWR _10822_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19306_ _04270_ _04332_ _04244_ _04598_ _03705_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__o221a_1
X_16518_ _11396_ _12481_ _12482_ _12483_ VGND VGND VPWR VPWR _12484_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17498_ _13183_ _13443_ _13444_ _13445_ VGND VGND VPWR VPWR _13446_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19237_ _04516_ _04465_ _04524_ _04531_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__a2bb2o_1
X_16449_ _11346_ decode.regfile.registers_30\[30\] _12095_ _12096_ _12097_ VGND VGND
+ VPWR VPWR _12416_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_136_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19168_ _09974_ _03771_ _03970_ _03969_ _04289_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18119_ _10915_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19099_ _04392_ _04316_ _04393_ _04394_ net318 VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__a32o_1
XFILLER_0_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21130_ _06057_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21061_ execute.csr_read_data_out_reg\[19\] _06014_ _06010_ VGND VGND VPWR VPWR _06017_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20012_ _05232_ _05233_ _05235_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_35_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24820_ _08597_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24751_ _08113_ net1355 _06283_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21963_ net777 _06572_ _06583_ _06579_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23702_ _08001_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20914_ _05857_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__buf_2
X_27470_ clknet_leaf_27_clock _00499_ VGND VGND VPWR VPWR csr.io_csr_address\[4\]
+ sky130_fd_sc_hd__dfxtp_4
X_24682_ _08524_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21894_ csr._mcycle_T_2\[17\] _06521_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__or2_1
X_26421_ _09402_ _09545_ VGND VGND VPWR VPWR _09552_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_169_Left_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23633_ _07964_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20845_ _03582_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__buf_2
XFILLER_0_194_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29140_ clknet_leaf_91_clock _02153_ VGND VGND VPWR VPWR csr.mcycle\[24\] sky130_fd_sc_hd__dfxtp_2
X_26352_ net1167 _09505_ _09511_ _09512_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23564_ net88 _07917_ _07926_ _05805_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20776_ _05857_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25303_ _08882_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22515_ fetch.bht.bhtTable_target_pc\[2\]\[1\] fetch.bht.bhtTable_target_pc\[3\]\[1\]
+ _07108_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__mux2_1
X_29071_ clknet_leaf_208_clock _02084_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26283_ _09412_ _09472_ VGND VGND VPWR VPWR _09473_ sky130_fd_sc_hd__nand2_1
X_23495_ net650 _07875_ _07886_ _07879_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__o211a_1
X_28022_ clknet_leaf_207_clock _01044_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25234_ _08846_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22446_ _06645_ fetch.btb.btbTable\[15\]\[1\] fetch.bht.bhtTable_valid\[15\] _06627_
+ _07040_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__a311o_1
XFILLER_0_150_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25165_ _08801_ _09880_ _09884_ VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__or3b_1
X_22377_ _06971_ _06730_ _06686_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24116_ net852 execute.io_target_pc\[13\] _08221_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__mux2_1
X_21328_ _06174_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25096_ _06113_ net1745 _08596_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28924_ clknet_leaf_182_clock _01937_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24047_ _08195_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__clkbuf_1
X_21259_ csr.io_mem_pc\[21\] VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold480 decode.regfile.registers_4\[0\] VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 decode.regfile.registers_12\[6\] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__dlygate4sd3_1
X_28855_ clknet_leaf_124_clock _01868_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15820_ decode.regfile.registers_1\[13\] _11115_ _11056_ _11108_ VGND VGND VPWR VPWR
+ _11804_ sky130_fd_sc_hd__nand4_1
XFILLER_0_102_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27806_ clknet_leaf_327_clock _00835_ VGND VGND VPWR VPWR memory.io_wb_readdata\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_28786_ clknet_leaf_106_clock _01799_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_25998_ net2742 _09286_ _09295_ _09292_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15751_ _11289_ _11735_ _11736_ VGND VGND VPWR VPWR _11737_ sky130_fd_sc_hd__o21ai_1
X_27737_ clknet_leaf_37_clock _00766_ VGND VGND VPWR VPWR decode.io_wb_rd\[0\] sky130_fd_sc_hd__dfxtp_4
X_24949_ net1109 _08678_ _08679_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1180 fetch.bht.bhtTable_tag\[0\]\[21\] VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14702_ _10705_ execute.io_target_pc\[5\] _10692_ execute.io_target_pc\[19\] _10744_
+ VGND VGND VPWR VPWR _10745_ sky130_fd_sc_hd__o221a_1
Xhold1191 _01237_ VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18470_ _09921_ _03645_ _03641_ _03643_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__nand4_4
X_15682_ decode.regfile.registers_19\[9\] _11354_ _11218_ _11669_ VGND VGND VPWR VPWR
+ _11670_ sky130_fd_sc_hd__o211a_1
X_27668_ clknet_leaf_27_clock _00697_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_219_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _13087_ decode.regfile.registers_26\[15\] _13254_ _13047_ _13088_ VGND VGND
+ VPWR VPWR _13371_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_206_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14633_ _10674_ decode.id_ex_pc_reg\[1\] _10675_ execute.io_target_pc\[16\] VGND
+ VGND VPWR VPWR _10676_ sky130_fd_sc_hd__a22oi_2
X_26619_ _10245_ _09666_ VGND VGND VPWR VPWR _09667_ sky130_fd_sc_hd__nand2_1
X_29407_ clknet_leaf_247_clock _02420_ VGND VGND VPWR VPWR decode.regfile.registers_5\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_27599_ clknet_leaf_152_clock _00628_ VGND VGND VPWR VPWR execute.io_target_pc\[8\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_68_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_215_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _12701_ decode.regfile.registers_28\[14\] _12698_ VGND VGND VPWR VPWR _13303_
+ sky130_fd_sc_hd__o21a_1
X_29338_ clknet_leaf_256_clock _02351_ VGND VGND VPWR VPWR decode.regfile.registers_3\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14564_ decode.immGen._imm_T_24\[16\] VGND VGND VPWR VPWR _10607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16303_ _11942_ net496 _12095_ _12096_ _12097_ VGND VGND VPWR VPWR _12274_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_172_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13515_ _09893_ VGND VGND VPWR VPWR _09894_ sky130_fd_sc_hd__buf_2
X_29269_ clknet_5_29__leaf_clock _02282_ VGND VGND VPWR VPWR decode.regfile.registers_0\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_17283_ decode.regfile.registers_10\[12\] _12600_ _12724_ VGND VGND VPWR VPWR _13236_
+ sky130_fd_sc_hd__a21oi_1
X_14495_ net605 _10533_ _10543_ _10535_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19022_ _04014_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16234_ decode.regfile.registers_7\[24\] _11092_ _11142_ _11169_ decode.regfile.registers_6\[24\]
+ VGND VGND VPWR VPWR _12207_ sky130_fd_sc_hd__a32o_1
XFILLER_0_180_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16165_ _12138_ _11154_ _11190_ _11148_ _12139_ VGND VGND VPWR VPWR _12140_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_144_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15116_ _11112_ VGND VGND VPWR VPWR _11113_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16096_ _11690_ _12072_ VGND VGND VPWR VPWR _12073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19924_ _05187_ _05188_ _05191_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__o21bai_1
X_15047_ _11043_ VGND VGND VPWR VPWR _11044_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_228_Right_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19855_ _05045_ _05046_ _05049_ _03852_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_78_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18806_ _04096_ _03699_ net249 decode.id_ex_rs1_data_reg\[13\] _04099_ VGND VGND
+ VPWR VPWR _04105_ sky130_fd_sc_hd__o221a_4
XTAP_TAPCELL_ROW_30_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19786_ _03838_ _03835_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_30_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16998_ _12915_ decode.regfile.registers_25\[5\] _12506_ _12812_ VGND VGND VPWR VPWR
+ _12958_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_69_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18737_ decode.id_ex_rs2_data_reg\[4\] net199 _04035_ VGND VGND VPWR VPWR _04036_
+ sky130_fd_sc_hd__o21ai_2
X_15949_ _10652_ _11112_ _11118_ _11929_ VGND VGND VPWR VPWR _11930_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_125_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18668_ net125 _03664_ _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17619_ _02986_ decode.regfile.registers_26\[20\] _13254_ _13484_ _02987_ VGND VGND
+ VPWR VPWR _03026_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_59_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18599_ _10080_ _03785_ _03897_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_50_1110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20630_ csr.mscratch\[26\] _05593_ _05625_ _05762_ _05763_ VGND VGND VPWR VPWR _05764_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20561_ _05704_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22300_ net80 _06833_ _06698_ net225 VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23280_ fetch.bht.bhtTable_target_pc\[12\]\[22\] fetch.bht.bhtTable_target_pc\[13\]\[22\]
+ fetch.bht.bhtTable_target_pc\[14\]\[22\] fetch.bht.bhtTable_target_pc\[15\]\[22\]
+ _07555_ _07710_ VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20492_ _05644_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__buf_1
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22231_ _06632_ _06825_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22162_ _06678_ _06756_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21113_ _06048_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22093_ _06683_ _06685_ _06687_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26970_ net2157 _09866_ _09868_ _09865_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_58_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout223 net81 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21044_ _06007_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__clkbuf_1
X_25921_ _08918_ _09243_ VGND VGND VPWR VPWR _09251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28640_ clknet_leaf_171_clock _01653_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25852_ net593 _09199_ _09211_ _09209_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24803_ _08588_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__clkbuf_1
X_28571_ clknet_leaf_187_clock _01584_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_25783_ _08931_ _09166_ VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__nand2_1
X_22995_ fetch.bht.bhtTable_target_pc\[12\]\[6\] fetch.bht.bhtTable_target_pc\[13\]\[6\]
+ _07439_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_177_Left_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27522_ clknet_leaf_43_clock _00551_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_2
X_24734_ _08551_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__clkbuf_1
X_21946_ _06457_ _06459_ _06470_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__and3b_2
XFILLER_0_69_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27453_ clknet_leaf_160_clock _00482_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[19\]
+ sky130_fd_sc_hd__dfxtp_2
X_24665_ net767 execute.io_target_pc\[21\] _08508_ VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21877_ _06523_ _06519_ _06520_ _06524_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26404_ net2325 _09534_ _09542_ _09540_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__o211a_1
X_23616_ _07954_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20828_ net101 _05879_ _05887_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__and3_1
X_27384_ clknet_leaf_15_clock _00413_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_24596_ _08480_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29123_ clknet_leaf_74_clock _02136_ VGND VGND VPWR VPWR csr.mcycle\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26335_ _09389_ _09502_ VGND VGND VPWR VPWR _09503_ sky130_fd_sc_hd__nand2_1
X_23547_ _03546_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20759_ _05848_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_210_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_210_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29054_ clknet_leaf_130_clock _02067_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26266_ net796 _09462_ _09463_ _09458_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__o211a_1
X_14280_ _10420_ _10245_ VGND VGND VPWR VPWR _10421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23478_ net17 _07875_ _07877_ _07865_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__o211a_2
XFILLER_0_45_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28005_ clknet_leaf_202_clock _01027_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_186_Left_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25217_ _08055_ net1527 _08837_ VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__mux2_1
X_22429_ _06790_ _07019_ _07021_ _07023_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__o22a_1
XFILLER_0_162_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26197_ _09417_ VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__buf_2
XFILLER_0_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25148_ _06281_ _08801_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25079_ _03580_ _08767_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17970_ _02986_ decode.regfile.registers_26\[29\] _13002_ _11010_ _02987_ VGND VGND
+ VPWR VPWR _03368_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_208_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28907_ clknet_leaf_93_clock _01920_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16921_ _12508_ VGND VGND VPWR VPWR _12882_ sky130_fd_sc_hd__buf_4
X_29887_ clknet_leaf_304_clock _02900_ VGND VGND VPWR VPWR decode.regfile.registers_20\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19640_ _04280_ _04282_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__or3b_1
XFILLER_0_218_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28838_ clknet_leaf_96_clock _01851_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16852_ _10928_ decode.regfile.registers_26\[2\] _12814_ _11011_ _11027_ VGND VGND
+ VPWR VPWR _12815_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_102_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_195_Left_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15803_ decode.regfile.registers_20\[12\] _11452_ _11223_ _11787_ VGND VGND VPWR
+ VPWR _11788_ sky130_fd_sc_hd__a211o_1
XFILLER_0_205_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19571_ _04408_ _04293_ _04386_ _04846_ _04853_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__o311a_2
X_16783_ decode.regfile.registers_12\[1\] _12489_ _12498_ _12540_ VGND VGND VPWR VPWR
+ _12747_ sky130_fd_sc_hd__or4_1
X_28769_ clknet_leaf_175_clock _01782_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_13995_ _10015_ _10255_ VGND VGND VPWR VPWR _10256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_217_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15734_ _11445_ _11719_ _11720_ VGND VGND VPWR VPWR _11721_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18522_ _03817_ _03819_ _03775_ _03820_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_38_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_213_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ decode.regfile.registers_1\[9\] decode.regfile.registers_0\[9\] _11300_ VGND
+ VGND VPWR VPWR _11653_ sky130_fd_sc_hd__mux2_1
X_18453_ _03711_ _03712_ _09921_ _03713_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__o211a_4
XFILLER_0_197_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_150 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_1344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14616_ decode.immGen._imm_T_24\[3\] VGND VGND VPWR VPWR _10659_ sky130_fd_sc_hd__clkbuf_4
X_17404_ _12541_ _12772_ _13352_ _13353_ VGND VGND VPWR VPWR _13354_ sky130_fd_sc_hd__o211ai_1
X_18384_ decode.id_ex_ex_rs1_reg\[0\] decode.io_wb_rd\[0\] VGND VGND VPWR VPWR _03683_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_201_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15596_ decode.regfile.registers_8\[7\] _11044_ _11174_ VGND VGND VPWR VPWR _11586_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17335_ decode.regfile.registers_21\[13\] _12681_ VGND VGND VPWR VPWR _13287_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14547_ _10589_ decode.id_ex_ex_rd_reg\[2\] VGND VGND VPWR VPWR _10590_ sky130_fd_sc_hd__xor2_1
XFILLER_0_166_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17266_ _12708_ net457 _13181_ _13218_ _13219_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__o221a_1
X_14478_ _10426_ VGND VGND VPWR VPWR _10535_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19005_ _04279_ _04019_ _04028_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__or3_2
X_16217_ decode.regfile.registers_18\[23\] _10955_ _11114_ _11094_ _10976_ VGND VGND
+ VPWR VPWR _12191_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_12_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17197_ decode.regfile.registers_10\[10\] _12598_ _13150_ _13151_ VGND VGND VPWR
+ VPWR _13152_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_183_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16148_ decode.regfile.registers_20\[21\] _11452_ _11223_ _12123_ VGND VGND VPWR
+ VPWR _12124_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16079_ decode.regfile.registers_14\[20\] _10639_ VGND VGND VPWR VPWR _12056_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_90_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19907_ _04317_ _04439_ _04410_ _04949_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1905 fetch.bht.bhtTable_tag\[5\]\[7\] VGND VGND VPWR VPWR net2132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1916 _01244_ VGND VGND VPWR VPWR net2143 sky130_fd_sc_hd__dlygate4sd3_1
X_19838_ _04492_ _05096_ _05097_ _05109_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__nor4_1
XFILLER_0_208_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1927 decode.io_id_pc\[29\] VGND VGND VPWR VPWR net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1938 decode.regfile.registers_16\[7\] VGND VGND VPWR VPWR net2165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1949 decode.regfile.registers_10\[4\] VGND VGND VPWR VPWR net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xinput1 net381 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_19769_ _04509_ _04369_ _04905_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21800_ net2626 _06467_ _06468_ _10546_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22780_ _07283_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21731_ _06426_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__buf_6
XFILLER_0_148_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24450_ _08404_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__clkbuf_1
X_21662_ _06373_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23401_ fetch.bht.bhtTable_target_pc\[0\]\[30\] fetch.bht.bhtTable_target_pc\[1\]\[30\]
+ fetch.bht.bhtTable_target_pc\[2\]\[30\] fetch.bht.bhtTable_target_pc\[3\]\[30\]
+ _07106_ _07386_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20613_ csr.mcycle\[24\] _05587_ _05575_ csr.minstret\[24\] VGND VGND VPWR VPWR _05749_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24381_ net996 execute.io_target_pc\[13\] _08367_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21593_ _06317_ csr.io_inst_retired VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__and2_1
X_26120_ _08966_ _09353_ VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23332_ _07064_ _07747_ _07748_ _07759_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20544_ csr._minstret_T_3\[46\] _05538_ _05658_ _05689_ VGND VGND VPWR VPWR _05690_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26051_ _08973_ _09285_ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__nand2_1
X_23263_ fetch.bht.bhtTable_target_pc\[6\]\[21\] fetch.bht.bhtTable_target_pc\[7\]\[21\]
+ _07068_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20475_ _03594_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25002_ _03558_ _08714_ _08701_ VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22214_ net276 VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23194_ _07626_ _07130_ _03592_ _07629_ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29810_ clknet_leaf_295_clock _02823_ VGND VGND VPWR VPWR decode.regfile.registers_17\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_22145_ _06642_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29741_ clknet_leaf_285_clock _02754_ VGND VGND VPWR VPWR decode.regfile.registers_15\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22076_ net87 _06656_ _06670_ net221 VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__a2bb2o_1
X_26953_ net649 _09853_ _09858_ _09852_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__o211a_1
X_25904_ _09930_ _10194_ _10196_ _08902_ VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__and4b_1
X_21027_ _03582_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_227_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29672_ clknet_leaf_277_clock _02685_ VGND VGND VPWR VPWR decode.regfile.registers_13\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_26884_ net2088 _09809_ _09818_ _09812_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28623_ clknet_leaf_111_clock _01636_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_25835_ _08982_ _09200_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_195_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28554_ clknet_leaf_223_clock _01567_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13780_ net1932 _10083_ _10118_ _10077_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__o211a_1
X_25766_ _08914_ _09157_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22978_ _07127_ _07421_ _07423_ _07425_ _07367_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_195_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24717_ _08078_ net1738 _08542_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__mux2_1
X_27505_ clknet_leaf_21_clock _00534_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28485_ clknet_leaf_196_clock _01498_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_21929_ _06559_ _06543_ _06544_ _06560_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25697_ net2332 _09111_ _09121_ _09115_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_191_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27436_ clknet_leaf_146_clock _00465_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15450_ _11344_ net918 _11402_ _11443_ _11249_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__o221a_1
X_24648_ net1202 execute.io_target_pc\[13\] _08497_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_191_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14401_ _10462_ VGND VGND VPWR VPWR _10490_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15381_ _11368_ _11374_ _11375_ decode.regfile.registers_4\[2\] VGND VGND VPWR VPWR
+ _11376_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_38_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27367_ clknet_leaf_30_clock _00396_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_24579_ _08471_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17120_ decode.regfile.registers_19\[8\] _11013_ _10589_ _12519_ _12544_ VGND VGND
+ VPWR VPWR _13077_ sky130_fd_sc_hd__o41a_1
XFILLER_0_93_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29106_ clknet_leaf_17_clock _02119_ VGND VGND VPWR VPWR csr._mcycle_T_3\[54\] sky130_fd_sc_hd__dfxtp_1
X_14332_ net1408 _10447_ _10450_ _10440_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__o211a_1
X_26318_ net603 _09491_ _09493_ _09484_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27298_ clknet_leaf_0_clock _00327_ VGND VGND VPWR VPWR decode.regfile.registers_31\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29037_ clknet_leaf_103_clock _02050_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_17051_ _10931_ net467 _12487_ VGND VGND VPWR VPWR _13009_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _10117_ _10400_ VGND VGND VPWR VPWR _10410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26249_ net587 _09447_ _09453_ _09440_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_150_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap209 _12638_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_1
X_16002_ _11646_ _11834_ _11944_ decode.regfile.registers_29\[17\] _11981_ VGND VGND
+ VPWR VPWR _11982_ sky130_fd_sc_hd__o221a_1
XFILLER_0_151_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14194_ _10136_ _10331_ VGND VGND VPWR VPWR _10370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29939_ clknet_leaf_340_clock _02952_ VGND VGND VPWR VPWR decode.regfile.registers_21\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_17953_ _11018_ _12977_ _12510_ decode.regfile.registers_8\[29\] _12892_ VGND VGND
+ VPWR VPWR _03351_ sky130_fd_sc_hd__o32a_1
XFILLER_0_225_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16904_ _10928_ decode.regfile.registers_26\[3\] _12814_ _11011_ _11027_ VGND VGND
+ VPWR VPWR _12866_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17884_ _12650_ _12723_ _12669_ decode.regfile.registers_14\[27\] _03283_ VGND VGND
+ VPWR VPWR _03284_ sky130_fd_sc_hd__o221a_1
XFILLER_0_228_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19623_ _04805_ _04422_ _04729_ _04883_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16835_ _12667_ _12773_ _12670_ decode.regfile.registers_14\[2\] _12797_ VGND VGND
+ VPWR VPWR _12798_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_122_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19554_ _04785_ _04836_ _04186_ _04095_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16766_ decode.regfile.registers_1\[1\] decode.regfile.registers_0\[1\] _12630_ VGND
+ VGND VPWR VPWR _12730_ sky130_fd_sc_hd__mux2_1
X_13978_ net1310 _10243_ _10246_ _10232_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18505_ execute.csr_read_data_out_reg\[26\] _03659_ net118 _03666_ VGND VGND VPWR
+ VPWR _03804_ sky130_fd_sc_hd__o22a_1
X_15717_ _11132_ _11692_ _11703_ VGND VGND VPWR VPWR _11704_ sky130_fd_sc_hd__o21a_1
X_19485_ _04409_ _04556_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__nand2_1
X_16697_ _12661_ VGND VGND VPWR VPWR _12662_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18436_ decode.io_wb_regwrite decode.id_ex_ex_use_rs2_reg VGND VGND VPWR VPWR _03735_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15648_ decode.regfile.registers_20\[8\] _11103_ _11635_ _11636_ _11222_ VGND VGND
+ VPWR VPWR _11637_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15579_ _11346_ _11253_ _11064_ decode.regfile.registers_29\[6\] _11569_ VGND VGND
+ VPWR VPWR _11570_ sky130_fd_sc_hd__o221a_1
X_18367_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17318_ decode.regfile.registers_1\[13\] decode.regfile.registers_0\[13\] _12778_
+ VGND VGND VPWR VPWR _13270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18298_ decode.id_ex_rs2_data_reg\[15\] _03605_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17249_ decode.regfile.registers_15\[11\] _12874_ _13187_ _13202_ _12576_ VGND VGND
+ VPWR VPWR _13203_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_92_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20260_ _10731_ _10680_ _10707_ _05433_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__or4b_1
XFILLER_0_4_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20191_ _00575_ _05226_ _05390_ _05239_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1086 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2403 csr._csr_read_data_T_8\[17\] VGND VGND VPWR VPWR net2630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2414 decode.regfile.registers_3\[23\] VGND VGND VPWR VPWR net2641 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2425 decode.regfile.registers_11\[27\] VGND VGND VPWR VPWR net2652 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2436 decode.regfile.registers_0\[21\] VGND VGND VPWR VPWR net2663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23950_ _08145_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__clkbuf_1
Xhold1702 csr._mcycle_T_3\[50\] VGND VGND VPWR VPWR net1929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2447 decode.regfile.registers_0\[29\] VGND VGND VPWR VPWR net2674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1713 fetch.bht.bhtTable_tag\[5\]\[20\] VGND VGND VPWR VPWR net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2458 decode.regfile.registers_25\[4\] VGND VGND VPWR VPWR net2685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1724 _01238_ VGND VGND VPWR VPWR net1951 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2469 decode.regfile.registers_11\[28\] VGND VGND VPWR VPWR net2696 sky130_fd_sc_hd__dlygate4sd3_1
X_22901_ _06976_ _07351_ _06956_ _06964_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__or4bb_1
Xhold1735 fetch.bht.bhtTable_tag\[10\]\[2\] VGND VGND VPWR VPWR net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1746 fetch.bht.bhtTable_target_pc\[5\]\[3\] VGND VGND VPWR VPWR net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23881_ _08108_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__clkbuf_1
Xhold1757 decode.io_id_pc\[28\] VGND VGND VPWR VPWR net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_323_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_323_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1768 decode.regfile.registers_21\[20\] VGND VGND VPWR VPWR net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1779 csr.mscratch\[20\] VGND VGND VPWR VPWR net2006 sky130_fd_sc_hd__dlygate4sd3_1
X_25620_ net1677 _09068_ _09077_ _09074_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__o211a_1
X_22832_ net1147 csr.io_mem_pc\[29\] _07308_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25551_ _08925_ _09036_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22763_ _07274_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24502_ _08062_ net1439 _08428_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21714_ net762 _06413_ _06414_ _06352_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__a211oi_1
X_28270_ clknet_leaf_64_clock _01292_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25482_ _08933_ _08992_ VGND VGND VPWR VPWR _08998_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_338_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_338_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22694_ _07207_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27221_ clknet_leaf_5_clock _00250_ VGND VGND VPWR VPWR decode.regfile.registers_29\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24433_ _08395_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21645_ csr.minstret\[12\] csr.minstret\[13\] VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27152_ clknet_leaf_354_clock _00181_ VGND VGND VPWR VPWR decode.regfile.registers_27\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24364_ net1381 execute.io_target_pc\[5\] _08356_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21576_ _06147_ net1376 _06306_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__mux2_1
XANTENNA_50 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_61 _10935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26103_ net2172 _09343_ _09355_ _09346_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23315_ csr._csr_read_data_T_8\[24\] _07416_ csr.io_mret_vector\[24\] _07621_ _07743_
+ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__o221a_1
X_20527_ csr.mscratch\[12\] _03718_ _05554_ _05672_ _05674_ VGND VGND VPWR VPWR _05675_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_117_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27083_ clknet_leaf_347_clock _00112_ VGND VGND VPWR VPWR decode.regfile.registers_24\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_83 _12491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24295_ _06186_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_162_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_94 execute.io_reg_pc\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26034_ _08956_ _09310_ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__nand2_1
X_23246_ fetch.bht.bhtTable_target_pc\[0\]\[20\] fetch.bht.bhtTable_target_pc\[1\]\[20\]
+ fetch.bht.bhtTable_target_pc\[2\]\[20\] fetch.bht.bhtTable_target_pc\[3\]\[20\]
+ _07669_ _07100_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__mux4_1
X_20458_ _05541_ csr.io_mret_vector\[4\] _05602_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23177_ _07612_ _07613_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20389_ _05439_ _05201_ net1810 VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_205_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22128_ _06677_ _06722_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27985_ clknet_leaf_169_clock _01007_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_201_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ _10977_ VGND VGND VPWR VPWR _10978_ sky130_fd_sc_hd__clkbuf_4
X_29724_ clknet_leaf_311_clock _02737_ VGND VGND VPWR VPWR decode.regfile.registers_15\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_22059_ _06624_ _06647_ _06632_ _06653_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_201_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26936_ net1172 _09839_ _09848_ _09836_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_197_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ net784 _10199_ _10201_ _10188_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__o211a_1
X_14881_ _10912_ _10913_ _10916_ decode.immGen._imm_T_10\[3\] VGND VGND VPWR VPWR
+ _10920_ sky130_fd_sc_hd__and4bb_1
X_29655_ clknet_leaf_281_clock _02668_ VGND VGND VPWR VPWR decode.regfile.registers_12\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_26867_ _09794_ VGND VGND VPWR VPWR _09809_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_193_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28606_ clknet_leaf_177_clock _01619_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_193_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16620_ _12584_ VGND VGND VPWR VPWR _12585_ sky130_fd_sc_hd__clkbuf_4
X_13832_ _09993_ _10154_ VGND VGND VPWR VPWR _10160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25818_ _08966_ _09179_ VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__nand2_1
X_26798_ net558 _09766_ _09769_ _09758_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__o211a_1
X_29586_ clknet_leaf_275_clock _02599_ VGND VGND VPWR VPWR decode.regfile.registers_10\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16551_ _12515_ VGND VGND VPWR VPWR _12516_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28537_ clknet_leaf_196_clock _01550_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13763_ memory.io_wb_reg_pc\[24\] _10001_ VGND VGND VPWR VPWR _10104_ sky130_fd_sc_hd__and2_1
X_25749_ _08973_ _09110_ VGND VGND VPWR VPWR _09151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15502_ _11493_ decode.regfile.registers_24\[5\] _11065_ _11072_ _10990_ VGND VGND
+ VPWR VPWR _11494_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_211_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19270_ _04052_ _04557_ _04563_ _04504_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__a22o_1
X_16482_ _11396_ _12446_ _12447_ _12448_ VGND VGND VPWR VPWR _12449_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28468_ clknet_leaf_138_clock _01481_ VGND VGND VPWR VPWR decode.io_id_pc\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13694_ memory.csr_read_data_out_reg\[13\] _09942_ VGND VGND VPWR VPWR _10046_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18221_ csr.mcycle\[14\] csr.mcycle\[16\] csr.mcycle\[15\] csr.mcycle\[17\] VGND
+ VGND VPWR VPWR _03556_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_14_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15433_ decode.regfile.registers_18\[3\] _11269_ _11271_ VGND VGND VPWR VPWR _11427_
+ sky130_fd_sc_hd__a21oi_1
X_27419_ clknet_leaf_10_clock _00448_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[28\]
+ sky130_fd_sc_hd__dfxtp_2
X_28399_ clknet_leaf_143_clock _01412_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_152_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18152_ _03505_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__clkbuf_1
X_15364_ _11123_ VGND VGND VPWR VPWR _11359_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17103_ decode.regfile.registers_2\[8\] _12634_ _13058_ _13059_ _12629_ VGND VGND
+ VPWR VPWR _13060_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_41_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14315_ _10058_ _10431_ VGND VGND VPWR VPWR _10441_ sky130_fd_sc_hd__nand2_1
X_18083_ _03466_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15295_ _11290_ VGND VGND VPWR VPWR _11291_ sky130_fd_sc_hd__buf_4
XFILLER_0_180_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17034_ decode.regfile.registers_21\[6\] _12822_ _12909_ VGND VGND VPWR VPWR _12993_
+ sky130_fd_sc_hd__o21a_1
X_14246_ _10074_ _10400_ VGND VGND VPWR VPWR _10401_ sky130_fd_sc_hd__nand2_1
Xhold309 decode.regfile.registers_30\[4\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14177_ _10092_ _10355_ VGND VGND VPWR VPWR _10361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ net189 _03781_ _04253_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__mux2_2
XFILLER_0_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17936_ _02997_ _12767_ _12965_ decode.regfile.registers_29\[28\] _03334_ VGND VGND
+ VPWR VPWR _03335_ sky130_fd_sc_hd__o221a_1
Xhold1009 fetch.bht.bhtTable_target_pc\[13\]\[21\] VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17867_ decode.regfile.registers_10\[27\] _10617_ _12776_ _10610_ _12604_ VGND VGND
+ VPWR VPWR _03267_ sky130_fd_sc_hd__o2111a_1
Xclkbuf_2_2_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_2_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19606_ _04885_ _04867_ _03938_ _04201_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_85_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16818_ decode.regfile.registers_2\[2\] _10616_ _12729_ VGND VGND VPWR VPWR _12781_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_85_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17798_ decode.regfile.registers_9\[25\] _11019_ _12504_ _12511_ _12654_ VGND VGND
+ VPWR VPWR _03200_ sky130_fd_sc_hd__o41a_1
XFILLER_0_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19537_ _03638_ _04444_ _04095_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16749_ _12712_ decode.regfile.registers_24\[1\] _10604_ _12690_ _11025_ VGND VGND
+ VPWR VPWR _12713_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19468_ _04295_ _04752_ _04362_ _04754_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_240 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_251 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_262 net2800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18419_ csr.io_csr_address\[0\] VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_44_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_273 _10660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_284 _11058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19399_ _04684_ _04685_ _04526_ _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_295 _12754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21430_ _06218_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__buf_4
XFILLER_0_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21361_ _06109_ net1896 _06188_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_886 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23100_ _07539_ _07540_ _07371_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20312_ _05484_ _05485_ _03588_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__a21oi_1
X_24080_ _08212_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__clkbuf_1
X_21292_ _06154_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__clkbuf_1
Xhold810 fetch.bht.bhtTable_target_pc\[8\]\[8\] VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold821 csr.io_inst_retired VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 decode.regfile.registers_29\[18\] VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 fetch.bht.bhtTable_target_pc\[6\]\[24\] VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__dlygate4sd3_1
X_23031_ _07108_ fetch.bht.bhtTable_target_pc\[11\]\[8\] _07111_ VGND VGND VPWR VPWR
+ _07476_ sky130_fd_sc_hd__a21bo_1
X_20243_ _05432_ _05219_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__nor2_1
Xhold854 fetch.bht.bhtTable_target_pc\[13\]\[9\] VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 fetch.bht.bhtTable_tag\[2\]\[2\] VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 fetch.bht.bhtTable_tag\[11\]\[23\] VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 fetch.bht.bhtTable_tag\[4\]\[0\] VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__dlygate4sd3_1
X_20174_ _05374_ _05375_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__nand2_1
Xhold898 decode.regfile.registers_21\[1\] VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2200 decode.regfile.registers_13\[29\] VGND VGND VPWR VPWR net2427 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2211 decode.regfile.registers_15\[3\] VGND VGND VPWR VPWR net2438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2222 decode.regfile.registers_8\[20\] VGND VGND VPWR VPWR net2449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2233 csr._minstret_T_3\[62\] VGND VGND VPWR VPWR net2460 sky130_fd_sc_hd__dlygate4sd3_1
X_24982_ net447 _08699_ _08700_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__o21ba_1
X_27770_ clknet_leaf_327_clock _00799_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2244 decode.io_id_pc\[9\] VGND VGND VPWR VPWR net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1510 fetch.bht.bhtTable_target_pc\[9\]\[27\] VGND VGND VPWR VPWR net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2255 decode.regfile.registers_22\[27\] VGND VGND VPWR VPWR net2482 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_262_clock clknet_5_22__leaf_clock VGND VGND VPWR VPWR clknet_leaf_262_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1521 decode.regfile.registers_19\[22\] VGND VGND VPWR VPWR net1748 sky130_fd_sc_hd__dlygate4sd3_1
X_23933_ net814 _08091_ _08130_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__mux2_1
Xhold2266 decode.regfile.registers_28\[21\] VGND VGND VPWR VPWR net2493 sky130_fd_sc_hd__dlygate4sd3_1
X_26721_ net516 _09723_ _09725_ _09717_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__o211a_1
Xhold1532 fetch.bht.bhtTable_target_pc\[7\]\[2\] VGND VGND VPWR VPWR net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2277 decode.regfile.registers_1\[15\] VGND VGND VPWR VPWR net2504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1543 fetch.bht.bhtTable_target_pc\[3\]\[30\] VGND VGND VPWR VPWR net1770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2288 decode.regfile.registers_22\[23\] VGND VGND VPWR VPWR net2515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 fetch.bht.bhtTable_tag\[5\]\[14\] VGND VGND VPWR VPWR net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2299 decode.regfile.registers_16\[1\] VGND VGND VPWR VPWR net2526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1565 _10692_ VGND VGND VPWR VPWR net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1576 fetch.bht.bhtTable_target_pc\[10\]\[5\] VGND VGND VPWR VPWR net1803 sky130_fd_sc_hd__dlygate4sd3_1
X_26652_ _09406_ _09676_ VGND VGND VPWR VPWR _09685_ sky130_fd_sc_hd__nand2_1
X_29440_ clknet_leaf_250_clock _02453_ VGND VGND VPWR VPWR decode.regfile.registers_6\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_23864_ execute.io_target_pc\[23\] VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_165_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1587 fetch.bht.bhtTable_target_pc\[0\]\[19\] VGND VGND VPWR VPWR net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 fetch.bht.bhtTable_target_pc\[6\]\[15\] VGND VGND VPWR VPWR net1825 sky130_fd_sc_hd__dlygate4sd3_1
X_25603_ _09066_ VGND VGND VPWR VPWR _09067_ sky130_fd_sc_hd__clkbuf_4
X_22815_ net1004 csr.io_mem_pc\[21\] _07297_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__mux2_1
X_26583_ _09621_ VGND VGND VPWR VPWR _09645_ sky130_fd_sc_hd__buf_2
X_29371_ clknet_leaf_255_clock _02384_ VGND VGND VPWR VPWR decode.regfile.registers_4\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_23795_ _08050_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_277_clock clknet_5_21__leaf_clock VGND VGND VPWR VPWR clknet_leaf_277_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28322_ clknet_leaf_201_clock _01335_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25534_ net739 _09024_ _09028_ _09017_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22746_ _06119_ net1605 _07265_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28253_ clknet_leaf_79_clock _01275_ VGND VGND VPWR VPWR csr._minstret_T_3\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25465_ net2335 _08979_ _08987_ _08972_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22677_ net806 _07223_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_200_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_200_clock
+ sky130_fd_sc_hd__clkbuf_8
X_27204_ clknet_leaf_363_clock _00233_ VGND VGND VPWR VPWR decode.regfile.registers_28\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24416_ _08385_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__clkbuf_1
X_28184_ clknet_leaf_59_clock _01206_ VGND VGND VPWR VPWR csr.io_mret_vector\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_21628_ csr._mcycle_T_2\[9\] _06321_ _06346_ csr.minstret\[8\] net2763 VGND VGND
+ VPWR VPWR _06348_ sky130_fd_sc_hd__a221oi_1
X_25396_ net2504 _08928_ _08940_ _08927_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27135_ clknet_leaf_359_clock _00164_ VGND VGND VPWR VPWR decode.regfile.registers_26\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_24347_ _08109_ net1506 _06187_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__mux2_1
X_21559_ _06130_ net1566 _06295_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14100_ _10290_ VGND VGND VPWR VPWR _10317_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_6_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_6_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27066_ clknet_leaf_349_clock _00095_ VGND VGND VPWR VPWR decode.regfile.registers_24\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_15080_ _11074_ _11076_ decode.regfile.registers_24\[0\] VGND VGND VPWR VPWR _11077_
+ sky130_fd_sc_hd__and3_1
X_24278_ _08314_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_215_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_215_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14031_ net2411 _10271_ _10276_ _10275_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26017_ net2431 _09300_ _09306_ _09305_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__o211a_1
X_23229_ _07110_ _07662_ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_224_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_224_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18770_ decode.id_ex_rs1_data_reg\[6\] _03687_ _04068_ net355 VGND VGND VPWR VPWR
+ _04069_ sky130_fd_sc_hd__o22a_1
X_27968_ clknet_leaf_237_clock _00990_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_15982_ decode.regfile.registers_10\[17\] _10638_ _11132_ _11949_ _11961_ VGND VGND
+ VPWR VPWR _11962_ sky130_fd_sc_hd__o32a_1
XFILLER_0_101_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29707_ clknet_leaf_282_clock _02720_ VGND VGND VPWR VPWR decode.regfile.registers_14\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_17721_ _12612_ _03123_ _03124_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__o21ai_2
X_26919_ _09838_ VGND VGND VPWR VPWR _09839_ sky130_fd_sc_hd__clkbuf_4
X_14933_ _10961_ VGND VGND VPWR VPWR _10962_ sky130_fd_sc_hd__buf_4
XFILLER_0_175_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27899_ clknet_leaf_18_clock _00928_ VGND VGND VPWR VPWR csr._mcycle_T_2\[20\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_215_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29638_ clknet_leaf_278_clock _02651_ VGND VGND VPWR VPWR decode.regfile.registers_12\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_17652_ decode.regfile.registers_19\[21\] _11013_ _10589_ _12519_ _12544_ VGND VGND
+ VPWR VPWR _03058_ sky130_fd_sc_hd__o41a_1
XFILLER_0_199_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14864_ _10770_ _10780_ _10785_ _10857_ _10906_ VGND VGND VPWR VPWR _10907_ sky130_fd_sc_hd__o2111a_4
XFILLER_0_188_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ _12567_ VGND VGND VPWR VPWR _12568_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_19_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13815_ net2281 _09951_ _10148_ _10132_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__o211a_1
X_14795_ _10830_ _10831_ decode.id_ex_pc_reg\[4\] _10829_ _10837_ VGND VGND VPWR VPWR
+ _10838_ sky130_fd_sc_hd__o221ai_1
X_17583_ _02990_ _13176_ decode.regfile.registers_27\[19\] _13487_ VGND VGND VPWR
+ VPWR _02991_ sky130_fd_sc_hd__or4_1
X_29569_ clknet_leaf_252_clock _02582_ VGND VGND VPWR VPWR decode.regfile.registers_10\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19322_ _04582_ _04075_ _04172_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__a21bo_1
X_16534_ _12498_ VGND VGND VPWR VPWR _12499_ sky130_fd_sc_hd__buf_4
X_13746_ _10012_ memory.io_wb_aluresult\[21\] _09981_ memory.io_wb_readdata\[21\]
+ _09995_ VGND VGND VPWR VPWR _10090_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_175_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19253_ _04322_ _04318_ _04338_ _04547_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_73_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13677_ _10031_ _10016_ VGND VGND VPWR VPWR _10032_ sky130_fd_sc_hd__nand2_1
X_16465_ _11045_ decode.regfile.registers_12\[30\] _10649_ _11051_ _10631_ VGND VGND
+ VPWR VPWR _12432_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18204_ _10943_ _10941_ decode.control.io_funct3\[2\] VGND VGND VPWR VPWR _03542_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15416_ _11367_ VGND VGND VPWR VPWR _11410_ sky130_fd_sc_hd__buf_4
XFILLER_0_112_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16396_ decode.regfile.registers_16\[28\] _11359_ _12347_ _12364_ VGND VGND VPWR
+ VPWR _12365_ sky130_fd_sc_hd__o22a_1
X_19184_ _04338_ _04377_ _04479_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_53_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18135_ _03496_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15347_ _11253_ _11254_ _11342_ VGND VGND VPWR VPWR _11343_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_113_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18066_ _10964_ _10665_ _10969_ _10965_ _03455_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__a221o_1
X_15278_ _11273_ VGND VGND VPWR VPWR _11274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_184_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14229_ net764 _10390_ _10391_ _10385_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__o211a_1
X_17017_ _12889_ _12974_ _12975_ VGND VGND VPWR VPWR _12976_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18968_ _04260_ _04247_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_143_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ decode.regfile.registers_11\[28\] _12792_ _03307_ _03317_ VGND VGND VPWR
+ VPWR _03318_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18899_ _03911_ _03935_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_33_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_18 _02192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_29 _06730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20930_ _05937_ _05945_ net50 VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20861_ net117 _05903_ _05899_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22600_ csr._minstret_T_3\[48\] csr._minstret_T_3\[47\] csr._minstret_T_3\[46\] _07172_
+ VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__and4_1
XFILLER_0_117_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23580_ _06111_ net1552 _07930_ VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20792_ _05870_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22531_ _07101_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__buf_4
XFILLER_0_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25250_ _08089_ net1424 _08848_ VGND VGND VPWR VPWR _08855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22462_ _06635_ _07054_ _07056_ _06651_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24201_ _08095_ net1763 _08266_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21413_ _06221_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25181_ _08819_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__clkbuf_1
X_22393_ _06678_ _06985_ _06627_ _06987_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24132_ net1105 VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21344_ net975 csr.io_mem_pc\[29\] _06179_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28940_ clknet_leaf_108_clock _01953_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_24063_ net1318 execute.io_target_pc\[19\] _08198_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__mux2_1
Xhold640 fetch.bht.bhtTable_target_pc\[3\]\[0\] VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__dlygate4sd3_1
X_21275_ _10760_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold651 fetch.bht.bhtTable_target_pc\[11\]\[7\] VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold662 decode.regfile.registers_13\[5\] VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__dlygate4sd3_1
X_23014_ _07457_ _07458_ _07112_ _07459_ _07076_ VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_130_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold673 fetch.bht.bhtTable_target_pc\[3\]\[15\] VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd3_1
X_20226_ _05417_ _05230_ _05419_ _05414_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28871_ clknet_leaf_115_clock _01884_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold684 fetch.bht.bhtTable_target_pc\[12\]\[19\] VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold695 fetch.bht.bhtTable_tag\[10\]\[17\] VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27822_ clknet_leaf_318_clock _00851_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_20157_ _05359_ _05360_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_5_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2030 decode.regfile.registers_11\[2\] VGND VGND VPWR VPWR net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2041 fetch.bht.bhtTable_tag\[13\]\[10\] VGND VGND VPWR VPWR net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2052 decode.regfile.registers_3\[17\] VGND VGND VPWR VPWR net2279 sky130_fd_sc_hd__dlygate4sd3_1
X_27753_ clknet_leaf_322_clock _00782_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2063 execute.csr_write_data_out_reg\[27\] VGND VGND VPWR VPWR net2290 sky130_fd_sc_hd__dlygate4sd3_1
X_24965_ csr._mcycle_T_3\[57\] csr._mcycle_T_3\[56\] _08687_ _07148_ VGND VGND VPWR
+ VPWR _08690_ sky130_fd_sc_hd__a31o_1
X_20088_ decode.id_ex_imm_reg\[13\] _10710_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__nor2_1
Xhold2074 execute.csr_write_data_out_reg\[0\] VGND VGND VPWR VPWR net2301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2085 fetch.bht.bhtTable_target_pc\[13\]\[6\] VGND VGND VPWR VPWR net2312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1340 fetch.bht.bhtTable_target_pc\[10\]\[25\] VGND VGND VPWR VPWR net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1351 fetch.bht.bhtTable_tag\[7\]\[23\] VGND VGND VPWR VPWR net1578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2096 csr._minstret_T_3\[35\] VGND VGND VPWR VPWR net2323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26704_ net2495 _09709_ _09715_ _09702_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__o211a_1
Xhold1362 fetch.bht.bhtTable_target_pc\[0\]\[6\] VGND VGND VPWR VPWR net1589 sky130_fd_sc_hd__dlygate4sd3_1
X_23916_ net981 _08074_ _08119_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__mux2_1
Xhold1373 fetch.bht.bhtTable_tag\[7\]\[15\] VGND VGND VPWR VPWR net1600 sky130_fd_sc_hd__dlygate4sd3_1
X_24896_ csr.mcycle\[20\] _03554_ _08644_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__and3_1
X_27684_ clknet_leaf_29_clock _00713_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1384 fetch.bht.bhtTable_tag\[10\]\[25\] VGND VGND VPWR VPWR net1611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 decode.regfile.registers_28\[14\] VGND VGND VPWR VPWR net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29423_ clknet_leaf_260_clock _02436_ VGND VGND VPWR VPWR decode.regfile.registers_5\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_23847_ _08085_ net1480 _08079_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__mux2_1
X_26635_ net1160 _09665_ _09674_ _09675_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13600_ net211 VGND VGND VPWR VPWR _09964_ sky130_fd_sc_hd__buf_6
XFILLER_0_68_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29354_ clknet_leaf_228_clock _02367_ VGND VGND VPWR VPWR decode.regfile.registers_3\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_14580_ decode.immGen._imm_T_24\[1\] VGND VGND VPWR VPWR _10623_ sky130_fd_sc_hd__inv_2
X_23778_ _09905_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26566_ _09621_ VGND VGND VPWR VPWR _09636_ sky130_fd_sc_hd__buf_2
XFILLER_0_156_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28305_ clknet_leaf_166_clock _01318_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13531_ net704 _09907_ VGND VGND VPWR VPWR _09908_ sky130_fd_sc_hd__or2b_1
X_22729_ _06103_ net1152 _09903_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__mux2_1
X_25517_ net2293 _09008_ _09016_ _09017_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29285_ clknet_leaf_242_clock _02298_ VGND VGND VPWR VPWR decode.regfile.registers_1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26497_ net720 _09592_ _09596_ _09595_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_188_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16250_ _12222_ decode.regfile.registers_17\[24\] _11357_ VGND VGND VPWR VPWR _12223_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28236_ clknet_leaf_77_clock _01258_ VGND VGND VPWR VPWR csr._minstret_T_3\[36\]
+ sky130_fd_sc_hd__dfxtp_2
X_25448_ net1405 _08907_ _08976_ _08972_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15201_ _11197_ VGND VGND VPWR VPWR _11198_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_209_Right_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16181_ _10988_ _11113_ _11119_ _11203_ decode.regfile.registers_16\[22\] VGND VGND
+ VPWR VPWR _12156_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28167_ clknet_leaf_53_clock _01189_ VGND VGND VPWR VPWR csr.io_mret_vector\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25379_ _10030_ VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_154_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_154_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15132_ _10645_ VGND VGND VPWR VPWR _11129_ sky130_fd_sc_hd__buf_4
X_27118_ clknet_leaf_329_clock _00147_ VGND VGND VPWR VPWR decode.regfile.registers_25\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_28098_ clknet_leaf_74_clock _01120_ VGND VGND VPWR VPWR csr.minstret\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_226_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19940_ _03581_ _05201_ net953 VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__and3b_1
X_27049_ clknet_leaf_346_clock _00078_ VGND VGND VPWR VPWR decode.regfile.registers_23\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_15063_ _11059_ VGND VGND VPWR VPWR _11060_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_147_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14014_ net1398 _10258_ _10266_ _10262_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__o211a_1
X_19871_ _04503_ _04772_ _04294_ net219 _05140_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__a41o_1
Xclkbuf_leaf_169_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_169_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18822_ _04086_ _04095_ _04107_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_207_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18753_ _04050_ _04051_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__nor2_2
XFILLER_0_218_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15965_ _11435_ decode.regfile.registers_24\[17\] _11244_ _11080_ _11079_ VGND VGND
+ VPWR VPWR _11945_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_106_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17704_ _02997_ _13262_ _12965_ decode.regfile.registers_29\[22\] _03108_ VGND VGND
+ VPWR VPWR _03109_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14916_ decode.control.io_funct3\[2\] VGND VGND VPWR VPWR _10946_ sky130_fd_sc_hd__clkbuf_4
X_18684_ _03977_ _03979_ _03982_ net353 VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__a31o_2
X_15896_ decode.regfile.registers_14\[15\] _11208_ _11274_ decode.regfile.registers_15\[15\]
+ _11202_ VGND VGND VPWR VPWR _11878_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17635_ _12732_ _03037_ _03038_ _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_177_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14847_ _10889_ _10887_ _10704_ VGND VGND VPWR VPWR _10890_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17566_ decode.regfile.registers_16\[19\] _12674_ _12901_ _02973_ VGND VGND VPWR
+ VPWR _02974_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_107_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_107_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14778_ csr.io_mem_pc\[7\] VGND VGND VPWR VPWR _10821_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_978 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19305_ _04269_ _04411_ _04597_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__a21o_1
X_16517_ _11446_ decode.regfile.registers_28\[31\] _11066_ _11037_ _11448_ VGND VGND
+ VPWR VPWR _12483_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_58_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13729_ _10074_ _10075_ VGND VGND VPWR VPWR _10076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17497_ _13087_ decode.regfile.registers_26\[17\] _13254_ _13047_ _13088_ VGND VGND
+ VPWR VPWR _13445_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19236_ _04526_ _04529_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16448_ _12133_ net445 _12382_ _12415_ _12132_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_136_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19167_ _04248_ _04460_ _04461_ _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__o31a_1
XFILLER_0_82_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16379_ decode.regfile.registers_13\[28\] _11276_ _11407_ decode.regfile.registers_12\[28\]
+ _11360_ VGND VGND VPWR VPWR _12348_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18118_ _03486_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_132_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19098_ _04263_ _04395_ _04228_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_170_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18049_ _12967_ _03442_ _03443_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__a31o_1
XFILLER_0_223_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21060_ _06016_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20011_ _05232_ _05233_ _05235_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_35_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_4__f_clock clknet_2_0_0_clock VGND VGND VPWR VPWR clknet_5_4__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_35_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24750_ _08559_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21962_ csr.mscratch\[6\] _06574_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23701_ net1883 _10872_ _07992_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20913_ _05936_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24681_ net1466 execute.io_target_pc\[29\] _07285_ VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21893_ csr.io_mret_vector\[17\] _10803_ _06515_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23632_ net1092 _10881_ _07961_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__mux2_1
X_26420_ net472 _09548_ _09551_ _09540_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__o211a_1
X_20844_ _05898_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__clkbuf_1
X_26351_ _09417_ VGND VGND VPWR VPWR _09512_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_194_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23563_ net2154 _07918_ _07915_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__or3b_1
XFILLER_0_49_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20775_ _03590_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25302_ _08880_ decode.regfile.registers_0\[12\] VGND VGND VPWR VPWR _08882_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22514_ _07107_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29070_ clknet_leaf_196_clock _02083_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26282_ _09446_ VGND VGND VPWR VPWR _09472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23494_ net2767 _07876_ _07873_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_71_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_71_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25233_ _08072_ net1032 _08837_ VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__mux2_1
X_28021_ clknet_leaf_221_clock _01043_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_22445_ _06617_ fetch.btb.btbTable\[14\]\[1\] fetch.bht.bhtTable_valid\[14\] VGND
+ VGND VPWR VPWR _07040_ sky130_fd_sc_hd__and3b_1
XFILLER_0_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25164_ _08810_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_21_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22376_ fetch.bht.bhtTable_tag\[14\]\[16\] fetch.bht.bhtTable_tag\[15\]\[16\] _06809_
+ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__mux2_1
X_24115_ _08230_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__clkbuf_1
X_21327_ net1132 csr.io_mem_pc\[21\] _06168_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_86_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_86_clock
+ sky130_fd_sc_hd__clkbuf_8
X_25095_ _08775_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24046_ net1051 execute.io_target_pc\[11\] _08187_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28923_ clknet_leaf_172_clock _01936_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_21258_ _06131_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold470 decode.regfile.registers_14\[4\] VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 csr.mcycle\[13\] VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold492 execute.csr_write_data_out_reg\[11\] VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__dlygate4sd3_1
X_20209_ _05404_ _05405_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__xnor2_1
X_28854_ clknet_leaf_123_clock _01867_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21189_ _06086_ _06082_ net405 VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27805_ clknet_leaf_328_clock _00834_ VGND VGND VPWR VPWR memory.io_wb_readdata\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_28785_ clknet_leaf_104_clock _01798_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25997_ _08918_ _09287_ VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__nand2_1
X_27736_ clknet_leaf_54_clock net418 VGND VGND VPWR VPWR fetch.bht.bhtTable_tag_MPORT_en
+ sky130_fd_sc_hd__dfxtp_4
X_15750_ decode.regfile.registers_7\[11\] _11465_ _11466_ decode.regfile.registers_6\[11\]
+ _11166_ VGND VGND VPWR VPWR _11736_ sky130_fd_sc_hd__a221oi_1
X_24948_ csr._mcycle_T_3\[51\] csr._mcycle_T_3\[50\] _08676_ _07148_ VGND VGND VPWR
+ VPWR _08679_ sky130_fd_sc_hd__a31o_1
Xhold1170 decode.regfile.registers_1\[9\] VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__dlygate4sd3_1
X_14701_ decode.id_ex_pc_reg\[29\] _10698_ _10732_ execute.io_target_pc\[23\] VGND
+ VGND VPWR VPWR _10744_ sky130_fd_sc_hd__o22a_1
Xhold1181 decode.regfile.registers_29\[22\] VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_24_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_24_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1192 decode.regfile.registers_14\[31\] VGND VGND VPWR VPWR net1419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15681_ _11106_ _11667_ _11668_ VGND VGND VPWR VPWR _11669_ sky130_fd_sc_hd__a21o_1
X_27667_ clknet_leaf_26_clock _00696_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_219_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24879_ csr.mcycle\[19\] csr.mcycle\[22\] csr.mcycle\[21\] csr.mcycle\[24\] VGND
+ VGND VPWR VPWR _08629_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_219_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17420_ _12915_ decode.regfile.registers_25\[15\] _13045_ _13294_ VGND VGND VPWR
+ VPWR _13370_ sky130_fd_sc_hd__or4_1
X_29406_ clknet_leaf_248_clock _02419_ VGND VGND VPWR VPWR decode.regfile.registers_5\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14632_ decode.id_ex_pc_reg\[16\] VGND VGND VPWR VPWR _10675_ sky130_fd_sc_hd__inv_2
X_26618_ _09664_ VGND VGND VPWR VPWR _09666_ sky130_fd_sc_hd__buf_2
X_27598_ clknet_leaf_153_clock _00627_ VGND VGND VPWR VPWR execute.io_target_pc\[7\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_184_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_215_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29337_ clknet_leaf_244_clock _02350_ VGND VGND VPWR VPWR decode.regfile.registers_2\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_17351_ _13055_ net439 _13097_ VGND VGND VPWR VPWR _13302_ sky130_fd_sc_hd__o21a_1
X_14563_ _10605_ VGND VGND VPWR VPWR _10606_ sky130_fd_sc_hd__buf_6
XFILLER_0_136_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26549_ net1533 _09622_ _09626_ _09619_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16302_ _12133_ net509 _12237_ _12273_ _12132_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13514_ csr.io_mem_pc\[2\] csr.io_mem_pc\[3\] VGND VGND VPWR VPWR _09893_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_39_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_39_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29268_ clknet_leaf_233_clock _02281_ VGND VGND VPWR VPWR decode.regfile.registers_0\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17282_ _13232_ _13233_ _13234_ VGND VGND VPWR VPWR _13235_ sky130_fd_sc_hd__a21oi_1
X_14494_ _10128_ _10505_ VGND VGND VPWR VPWR _10543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19021_ _04255_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__clkbuf_4
X_28219_ clknet_leaf_86_clock net2391 VGND VGND VPWR VPWR csr.mscratch\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16233_ decode.regfile.registers_12\[24\] _10648_ _10631_ _11051_ VGND VGND VPWR
+ VPWR _12206_ sky130_fd_sc_hd__or4_1
X_29199_ clknet_leaf_240_clock _02212_ VGND VGND VPWR VPWR fetch.btb.btbTable\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16164_ _11371_ decode.regfile.registers_0\[22\] VGND VGND VPWR VPWR _12139_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15115_ _11111_ VGND VGND VPWR VPWR _11112_ sky130_fd_sc_hd__clkbuf_4
X_16095_ decode.regfile.registers_11\[20\] _11364_ _12057_ _12071_ VGND VGND VPWR
+ VPWR _12072_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_192_Right_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19923_ _05189_ _05190_ _04505_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__o21ai_1
X_15046_ _11042_ VGND VGND VPWR VPWR _11043_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_220_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19854_ _05122_ _05101_ _03802_ _03801_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__nand4_1
XFILLER_0_120_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18805_ _04100_ _04103_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__or2_4
X_19785_ _04620_ _05058_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__nand2_2
X_16997_ _12516_ _12954_ _12955_ _12956_ VGND VGND VPWR VPWR _12957_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18736_ net308 _04032_ _03706_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_218_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15948_ _11123_ decode.regfile.registers_16\[16\] _11913_ _11928_ VGND VGND VPWR
+ VPWR _11929_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_69_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18667_ execute.csr_read_data_out_reg\[3\] _03657_ execute.io_reg_pc\[3\] _03662_
+ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__o22a_1
X_15879_ decode.regfile.registers_20\[14\] _11102_ _11327_ _11861_ VGND VGND VPWR
+ VPWR _11862_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17618_ _13407_ decode.regfile.registers_25\[20\] _13482_ _13294_ VGND VGND VPWR
+ VPWR _03025_ sky130_fd_sc_hd__or4_1
XFILLER_0_148_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18598_ net291 _03896_ decode.id_ex_rs2_data_reg\[19\] _03746_ _03727_ VGND VGND
+ VPWR VPWR _03897_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_138_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17549_ decode.regfile.registers_9\[19\] _12776_ _12604_ _12532_ _12599_ VGND VGND
+ VPWR VPWR _13495_ sky130_fd_sc_hd__a41o_1
XFILLER_0_157_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20560_ _05439_ _05703_ _03449_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_60_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19219_ _04514_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_99_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20491_ _10909_ _05643_ _09954_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__and3b_1
XFILLER_0_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22230_ fetch.bht.bhtTable_tag\[4\]\[15\] fetch.bht.bhtTable_tag\[5\]\[15\] fetch.bht.bhtTable_tag\[6\]\[15\]
+ fetch.bht.bhtTable_tag\[7\]\[15\] _06754_ _06622_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22161_ fetch.bht.bhtTable_tag\[4\]\[13\] fetch.bht.bhtTable_tag\[5\]\[13\] _06707_
+ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21112_ _05949_ _06046_ net908 VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__and3_1
XFILLER_0_218_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22092_ _06686_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__buf_4
XFILLER_0_112_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25920_ net1387 _09242_ _09249_ _09250_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__o211a_1
X_21043_ execute.csr_read_data_out_reg\[11\] _06002_ _05998_ VGND VGND VPWR VPWR _06007_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_100_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout224 net77 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25851_ _08922_ _09210_ VGND VGND VPWR VPWR _09211_ sky130_fd_sc_hd__nand2_1
X_24802_ _08095_ net1285 _08585_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__mux2_1
X_28570_ clknet_leaf_186_clock _01583_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_22994_ _07439_ fetch.bht.bhtTable_target_pc\[14\]\[6\] VGND VGND VPWR VPWR _07441_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_213_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25782_ net571 _09170_ _09171_ _09169_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27521_ clknet_leaf_43_clock _00550_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_2
X_24733_ _08095_ net1243 _08542_ VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__mux2_1
X_21945_ _06571_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_213_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24664_ _08515_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__clkbuf_1
X_27452_ clknet_leaf_150_clock _00481_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[18\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_167_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21876_ csr._mcycle_T_2\[11\] _06521_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23615_ _06145_ net2204 _07952_ VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26403_ _09383_ _09535_ VGND VGND VPWR VPWR _09542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20827_ _05889_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__clkbuf_1
X_24595_ net1356 execute.io_target_pc\[19\] _08473_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27383_ clknet_leaf_15_clock _00412_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[24\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_154_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29122_ clknet_leaf_68_clock _02135_ VGND VGND VPWR VPWR csr.mcycle\[6\] sky130_fd_sc_hd__dfxtp_2
X_23546_ net80 _07903_ _07916_ _07907_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26334_ _09490_ VGND VGND VPWR VPWR _09502_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20758_ _03452_ _05201_ csr.io_csr_address\[6\] VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_210_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29053_ clknet_leaf_178_clock _02066_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_210_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26265_ _09396_ _09459_ VGND VGND VPWR VPWR _09463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23477_ _10994_ _07876_ _07873_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__or3b_1
XFILLER_0_165_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20689_ _05809_ decode.id_ex_rs1_data_reg\[6\] _05798_ VGND VGND VPWR VPWR _05811_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28004_ clknet_leaf_198_clock _01026_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_25216_ _09905_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__clkbuf_8
X_22428_ _07022_ _06690_ _06627_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26196_ _10130_ VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25147_ _10568_ _09887_ VGND VGND VPWR VPWR _08801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22359_ _06952_ _06953_ _00002_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25078_ csr._mcycle_T_2\[29\] _08710_ _08765_ _08766_ VGND VGND VPWR VPWR _08767_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_103_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_208_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28906_ clknet_leaf_98_clock _01919_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_208_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24029_ net1451 execute.io_target_pc\[3\] _08014_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__mux2_1
X_16920_ decode.regfile.registers_4\[4\] _12618_ _12620_ decode.regfile.registers_5\[4\]
+ _12623_ VGND VGND VPWR VPWR _12881_ sky130_fd_sc_hd__a221oi_1
X_29886_ clknet_leaf_304_clock _02899_ VGND VGND VPWR VPWR decode.regfile.registers_20\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28837_ clknet_leaf_139_clock _01850_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16851_ _12759_ VGND VGND VPWR VPWR _12814_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15802_ decode.regfile.registers_19\[12\] _11453_ _11454_ _11786_ VGND VGND VPWR
+ VPWR _11787_ sky130_fd_sc_hd__o211a_1
X_19570_ _04409_ _04302_ _04851_ _04852_ _04515_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__o311a_1
X_28768_ clknet_leaf_170_clock _01781_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_16782_ _12724_ _12743_ _12744_ _12745_ VGND VGND VPWR VPWR _12746_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_217_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13994_ _10242_ VGND VGND VPWR VPWR _10255_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18521_ decode.id_ex_rs1_data_reg\[27\] _03689_ _10121_ _03772_ VGND VGND VPWR VPWR
+ _03820_ sky130_fd_sc_hd__a2bb2o_1
X_15733_ _11489_ decode.regfile.registers_28\[10\] decode.regfile.registers_29\[10\]
+ _11255_ _11246_ VGND VGND VPWR VPWR _11720_ sky130_fd_sc_hd__o221a_1
XFILLER_0_38_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27719_ clknet_leaf_20_clock _00748_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_217_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28699_ clknet_leaf_173_clock _01712_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _03718_ _03642_ _03748_ _03749_ _03750_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__o2111a_4
XTAP_TAPCELL_ROW_64_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _10647_ _11097_ decode.regfile.registers_5\[9\] VGND VGND VPWR VPWR _11652_
+ sky130_fd_sc_hd__or3b_1
XANTENNA_140 _12882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _12498_ _12504_ _12649_ decode.regfile.registers_11\[15\] VGND VGND VPWR
+ VPWR _13353_ sky130_fd_sc_hd__or4b_1
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14615_ _10657_ decode.id_ex_ex_rd_reg\[2\] VGND VGND VPWR VPWR _10658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_213_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18383_ _03680_ _09929_ _03681_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__a21oi_2
X_15595_ _11084_ _11297_ _11534_ decode.regfile.registers_6\[7\] _11584_ VGND VGND
+ VPWR VPWR _11585_ sky130_fd_sc_hd__o221a_1
XFILLER_0_200_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17334_ decode.regfile.registers_19\[13\] _12679_ _13264_ _13285_ _12545_ VGND VGND
+ VPWR VPWR _13286_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14546_ _10588_ VGND VGND VPWR VPWR _10589_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17265_ _12704_ VGND VGND VPWR VPWR _13219_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14477_ _10087_ _10530_ VGND VGND VPWR VPWR _10534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19004_ _04302_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16216_ _12189_ decode.regfile.registers_17\[23\] _11357_ VGND VGND VPWR VPWR _12190_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17196_ decode.regfile.registers_9\[10\] _11017_ _12503_ _12509_ _12652_ VGND VGND
+ VPWR VPWR _13151_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_168_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16147_ decode.regfile.registers_19\[21\] _11453_ _11454_ _12122_ VGND VGND VPWR
+ VPWR _12123_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16078_ decode.regfile.registers_23\[20\] _11087_ _11074_ _11049_ VGND VGND VPWR
+ VPWR _12055_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_90_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_22__f_clock clknet_2_2_0_clock VGND VGND VPWR VPWR clknet_5_22__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_220_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19906_ _04443_ _04415_ _05174_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__a21oi_1
X_15029_ _11033_ _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_127_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1906 decode.regfile.registers_16\[14\] VGND VGND VPWR VPWR net2133 sky130_fd_sc_hd__dlygate4sd3_1
X_19837_ _05099_ _05108_ _04589_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__a21oi_2
Xhold1917 fetch.bht.bhtTable_tag\[15\]\[17\] VGND VGND VPWR VPWR net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1928 decode.regfile.registers_27\[21\] VGND VGND VPWR VPWR net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1939 decode.regfile.registers_10\[13\] VGND VGND VPWR VPWR net2166 sky130_fd_sc_hd__dlygate4sd3_1
X_19768_ _04949_ _05039_ _05040_ _05042_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__o31a_1
XFILLER_0_127_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 net382 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_224_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18719_ decode.id_ex_imm_reg\[2\] VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19699_ _04973_ _04975_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21730_ _09885_ _09892_ _09916_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__and3_4
XFILLER_0_189_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21661_ _10019_ _06371_ _06372_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23400_ fetch.bht.bhtTable_target_pc\[4\]\[30\] fetch.bht.bhtTable_target_pc\[5\]\[30\]
+ fetch.bht.bhtTable_target_pc\[6\]\[30\] fetch.bht.bhtTable_target_pc\[7\]\[30\]
+ _07106_ _07070_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20612_ net770 _05537_ _05748_ _05454_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24380_ _09910_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21592_ _06320_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23331_ execute.io_target_pc\[25\] _07090_ _07089_ _07758_ _06032_ VGND VGND VPWR
+ VPWR _07759_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20543_ csr._csr_read_data_T_8\[14\] _05617_ _05686_ _05688_ _05616_ VGND VGND VPWR
+ VPWR _05689_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26050_ net2023 _09313_ _09324_ _09318_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__o211a_1
X_23262_ _07110_ _07693_ VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__or2b_1
XFILLER_0_144_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20474_ net1446 _05593_ _05625_ _05626_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__o32a_1
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25001_ csr.mcycle\[4\] csr.mcycle\[3\] _03557_ csr.mcycle\[5\] VGND VGND VPWR VPWR
+ _08714_ sky130_fd_sc_hd__a31oi_1
X_22213_ net69 _06794_ _06656_ _06795_ _06807_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__a221oi_2
X_23193_ _07627_ _07628_ _07391_ _07392_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22144_ _06635_ _06724_ _06728_ _06738_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__o31a_4
XFILLER_0_11_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29740_ clknet_leaf_284_clock _02753_ VGND VGND VPWR VPWR decode.regfile.registers_15\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_22075_ _06658_ _06663_ _06665_ _06669_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__a2bb2o_2
X_26952_ _10052_ _09849_ VGND VGND VPWR VPWR _09858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25903_ net2447 _09200_ _09239_ _09235_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__o211a_1
X_21026_ _05997_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__clkbuf_1
X_29671_ clknet_leaf_277_clock _02684_ VGND VGND VPWR VPWR decode.regfile.registers_13\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_26883_ _09410_ _09806_ VGND VGND VPWR VPWR _09818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_203_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28622_ clknet_leaf_112_clock _01635_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_25834_ net2199 _09199_ _09201_ _09194_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28553_ clknet_leaf_216_clock _01566_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_22977_ _07075_ _07424_ _07084_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25765_ net1246 _09156_ _09161_ _09153_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_195_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_195_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_27_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27504_ clknet_leaf_28_clock _00533_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dfxtp_1
X_24716_ _06282_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__clkbuf_8
X_28484_ clknet_leaf_202_clock _01497_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_21928_ csr._mcycle_T_2\[27\] _06545_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25696_ _08920_ _09112_ VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27435_ clknet_leaf_55_clock _00464_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24647_ _08506_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__clkbuf_1
X_21859_ csr.io_mret_vector\[7\] _10821_ _06040_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14400_ net454 _10477_ _10489_ _10481_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15380_ _10645_ _10627_ decode.immGen._imm_T_24\[11\] _11082_ VGND VGND VPWR VPWR
+ _11375_ sky130_fd_sc_hd__or4_4
XFILLER_0_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27366_ clknet_leaf_33_clock _00395_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_24578_ net1286 execute.io_target_pc\[11\] _08462_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29105_ clknet_leaf_17_clock _02118_ VGND VGND VPWR VPWR csr._mcycle_T_3\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14331_ _10097_ _10444_ VGND VGND VPWR VPWR _10450_ sky130_fd_sc_hd__nand2_1
X_26317_ _09025_ _09492_ VGND VGND VPWR VPWR _09493_ sky130_fd_sc_hd__nand2_1
X_23529_ net225 _07903_ _07906_ _07907_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27297_ clknet_leaf_0_clock _00326_ VGND VGND VPWR VPWR decode.regfile.registers_31\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29036_ clknet_leaf_108_clock _02049_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14262_ net779 _10403_ _10409_ _10398_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17050_ _13006_ _13007_ _12704_ _13008_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26248_ _09379_ _09448_ VGND VGND VPWR VPWR _09453_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16001_ _11403_ _11978_ _11979_ _11980_ VGND VGND VPWR VPWR _11981_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_36_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14193_ net675 _10359_ _10368_ _10369_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26179_ _09404_ _09390_ VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_1193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29938_ clknet_leaf_340_clock _02951_ VGND VGND VPWR VPWR decode.regfile.registers_21\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_17952_ _03348_ _03349_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16903_ _10939_ decode.regfile.registers_25\[3\] _12506_ _12812_ VGND VGND VPWR VPWR
+ _12865_ sky130_fd_sc_hd__or4_1
XFILLER_0_206_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17883_ _12658_ _03280_ _03281_ _03282_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__a31o_1
X_29869_ clknet_leaf_301_clock _02882_ VGND VGND VPWR VPWR decode.regfile.registers_19\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_19622_ _04546_ _04428_ _04692_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__a31o_1
XFILLER_0_219_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16834_ decode.regfile.registers_13\[2\] _12775_ _12795_ _12796_ _12664_ VGND VGND
+ VPWR VPWR _12797_ sky130_fd_sc_hd__a221o_1
XFILLER_0_206_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19553_ net283 _04103_ _04119_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__o21ai_1
X_16765_ _12728_ VGND VGND VPWR VPWR _12729_ sky130_fd_sc_hd__clkbuf_4
X_13977_ _10244_ _10245_ VGND VGND VPWR VPWR _10246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18504_ _03801_ _03802_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__nand2_2
XFILLER_0_38_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15716_ _11693_ _11701_ _11702_ VGND VGND VPWR VPWR _11703_ sky130_fd_sc_hd__o21ai_1
X_19484_ _04673_ _04769_ _04541_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16696_ _10598_ _10588_ _10610_ _12597_ VGND VGND VPWR VPWR _12661_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18435_ _03730_ _03731_ _03732_ _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__nand4_2
XFILLER_0_201_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15647_ decode.regfile.registers_19\[8\] _11049_ _11215_ _11217_ _11219_ VGND VGND
+ VPWR VPWR _11636_ sky130_fd_sc_hd__o41a_1
XFILLER_0_69_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18366_ _03664_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_173_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15578_ _11403_ _11566_ _11567_ _11568_ VGND VGND VPWR VPWR _11569_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17317_ _12882_ decode.regfile.registers_2\[13\] VGND VGND VPWR VPWR _13269_ sky130_fd_sc_hd__and2b_1
XFILLER_0_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14529_ _10572_ VGND VGND VPWR VPWR _10573_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_21_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18297_ _03613_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17248_ _10604_ _10619_ _12773_ _13188_ _13201_ VGND VGND VPWR VPWR _13202_ sky130_fd_sc_hd__o32a_1
XFILLER_0_142_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17179_ _12701_ decode.regfile.registers_28\[9\] _13093_ VGND VGND VPWR VPWR _13135_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20190_ _05389_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__inv_2
XFILLER_0_179_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2404 _01301_ VGND VGND VPWR VPWR net2631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2415 decode.regfile.registers_16\[24\] VGND VGND VPWR VPWR net2642 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2426 decode.regfile.registers_21\[26\] VGND VGND VPWR VPWR net2653 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2437 decode.regfile.registers_1\[16\] VGND VGND VPWR VPWR net2664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 fetch.bht.bhtTable_target_pc\[14\]\[3\] VGND VGND VPWR VPWR net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 fetch.btb.btbTable\[9\]\[1\] VGND VGND VPWR VPWR net2675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 fetch.bht.bhtTable_tag\[1\]\[19\] VGND VGND VPWR VPWR net1941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2459 decode.regfile.registers_8\[24\] VGND VGND VPWR VPWR net2686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1725 decode.regfile.registers_10\[26\] VGND VGND VPWR VPWR net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22900_ _06718_ _06717_ _07048_ _07058_ _07350_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__o2111ai_1
XTAP_TAPCELL_ROW_146_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23880_ _08107_ net1908 _07940_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__mux2_1
Xhold1736 fetch.bht.bhtTable_tag\[14\]\[14\] VGND VGND VPWR VPWR net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1747 fetch.bht.bhtTable_tag\[15\]\[13\] VGND VGND VPWR VPWR net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1758 fetch.bht.bhtTable_target_pc\[6\]\[7\] VGND VGND VPWR VPWR net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1769 fetch.bht.bhtTable_target_pc\[5\]\[23\] VGND VGND VPWR VPWR net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22831_ _07311_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22762_ _06136_ net922 _07265_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25550_ net471 _09024_ _09037_ _09033_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24501_ _08431_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__clkbuf_1
X_21713_ csr._mcycle_T_2\[28\] _06321_ _06413_ csr.minstret\[28\] VGND VGND VPWR VPWR
+ _06414_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_49_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25481_ net674 _08995_ _08997_ _08991_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__o211a_1
X_22693_ net2569 _07222_ _07233_ _07234_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27220_ clknet_leaf_7_clock _00249_ VGND VGND VPWR VPWR decode.regfile.registers_29\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_24432_ _08060_ net1584 _08389_ VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__mux2_1
X_21644_ net2444 _06357_ _06359_ _10546_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24363_ _08358_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27151_ clknet_leaf_352_clock _00180_ VGND VGND VPWR VPWR decode.regfile.registers_27\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_21575_ _06308_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_40 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_51 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23314_ _07089_ _07738_ _07739_ _07742_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_62 _10935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26102_ _08948_ _09353_ VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20526_ csr.minstret\[12\] _05571_ _05561_ csr.mcycle\[12\] _05673_ VGND VGND VPWR
+ VPWR _05674_ sky130_fd_sc_hd__a221o_1
X_27082_ clknet_leaf_346_clock _00111_ VGND VGND VPWR VPWR decode.regfile.registers_24\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_73 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24294_ _08322_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_84 _12491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_95 execute.io_reg_pc\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23245_ fetch.bht.bhtTable_target_pc\[4\]\[20\] fetch.bht.bhtTable_target_pc\[5\]\[20\]
+ fetch.bht.bhtTable_target_pc\[6\]\[20\] fetch.bht.bhtTable_target_pc\[7\]\[20\]
+ _07068_ _07656_ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__mux4_1
X_26033_ net2351 _09313_ _09315_ _09305_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__o211a_1
X_20457_ csr.minstret\[4\] VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__buf_2
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23176_ net74 net73 _07582_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__and3_2
X_20388_ _05549_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_205_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22127_ fetch.bht.bhtTable_tag\[8\]\[4\] fetch.bht.bhtTable_tag\[9\]\[4\] _06706_
+ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27984_ clknet_leaf_188_clock _01006_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29723_ clknet_leaf_312_clock _02736_ VGND VGND VPWR VPWR decode.regfile.registers_15\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22058_ _06648_ _06652_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__or2b_1
X_26935_ _10007_ _09840_ VGND VGND VPWR VPWR _09848_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_201_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13900_ _09950_ _10200_ VGND VGND VPWR VPWR _10201_ sky130_fd_sc_hd__nand2_1
X_21009_ _05988_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__clkbuf_1
X_29654_ clknet_leaf_281_clock _02667_ VGND VGND VPWR VPWR decode.regfile.registers_12\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_26866_ net544 _09795_ _09808_ _09799_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14880_ _10919_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__clkbuf_1
X_28605_ clknet_leaf_178_clock _01618_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_193_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13831_ net1520 _10153_ _10159_ _10132_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__o211a_1
X_25817_ net2579 _09183_ _09190_ _09182_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_3_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29585_ clknet_leaf_275_clock _02598_ VGND VGND VPWR VPWR decode.regfile.registers_10\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_26797_ _09400_ _09763_ VGND VGND VPWR VPWR _09769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28536_ clknet_leaf_196_clock _01549_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16550_ _12514_ VGND VGND VPWR VPWR _12515_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13762_ net2515 _10083_ _10103_ _10077_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__o211a_1
X_25748_ net2580 _09139_ _09150_ _09142_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15501_ _10956_ VGND VGND VPWR VPWR _11493_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28467_ clknet_leaf_139_clock _01480_ VGND VGND VPWR VPWR decode.io_id_pc\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_156_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16481_ _11446_ decode.regfile.registers_28\[30\] _11871_ _11037_ _11448_ VGND VGND
+ VPWR VPWR _12448_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_214_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13693_ _09943_ memory.io_wb_aluresult\[13\] _09981_ memory.io_wb_readdata\[13\]
+ VGND VGND VPWR VPWR _10045_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_85_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25679_ _09110_ VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__clkbuf_4
X_18220_ csr.mcycle\[22\] VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15432_ decode.regfile.registers_17\[3\] _11357_ _11425_ VGND VGND VPWR VPWR _11426_
+ sky130_fd_sc_hd__a21oi_1
X_27418_ clknet_leaf_10_clock _00447_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[27\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_14_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28398_ clknet_leaf_144_clock _01411_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18151_ _03495_ _03493_ _03500_ net2289 VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_155_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27349_ clknet_leaf_45_clock _00378_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[22\]
+ sky130_fd_sc_hd__dfxtp_2
X_15363_ decode.regfile.registers_17\[2\] _11357_ VGND VGND VPWR VPWR _11358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17102_ _12882_ _12933_ _12932_ decode.regfile.registers_0\[8\] VGND VGND VPWR VPWR
+ _13059_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14314_ net851 _10434_ _10439_ _10440_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__o211a_1
X_18082_ _03463_ _03464_ _03465_ decode.io_id_pc\[0\] VGND VGND VPWR VPWR _03466_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_29_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15294_ _11116_ _11091_ _11137_ VGND VGND VPWR VPWR _11290_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29019_ clknet_leaf_174_clock _02032_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17033_ decode.regfile.registers_20\[6\] _12771_ _12990_ _12991_ _12538_ VGND VGND
+ VPWR VPWR _12992_ sky130_fd_sc_hd__a221o_1
X_14245_ _10375_ VGND VGND VPWR VPWR _10400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14176_ net561 _10359_ _10360_ _10357_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_111_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_182_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _12967_ _03331_ _03332_ _03333_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__a31o_1
XFILLER_0_178_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17866_ decode.regfile.registers_15\[27\] _10611_ _10618_ _12588_ _12672_ VGND VGND
+ VPWR VPWR _03266_ sky130_fd_sc_hd__a41o_1
XFILLER_0_178_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16817_ decode.regfile.registers_1\[2\] _12778_ _12634_ _12779_ VGND VGND VPWR VPWR
+ _12780_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_1_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19605_ _04867_ _04885_ _04202_ _04526_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17797_ _03197_ _03198_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_85_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19536_ _04454_ _04818_ _04819_ _04496_ _04445_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__a221oi_1
X_16748_ _10926_ VGND VGND VPWR VPWR _12712_ sky130_fd_sc_hd__buf_2
XFILLER_0_221_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19467_ _04245_ _04542_ _04346_ _04753_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16679_ _11016_ _10597_ _10935_ _12637_ VGND VGND VPWR VPWR _12644_ sky130_fd_sc_hd__or4_1
XFILLER_0_192_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_230 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_241 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_252 net200 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18418_ execute.io_mem_rd\[4\] csr.io_csr_address\[4\] VGND VGND VPWR VPWR _03717_
+ sky130_fd_sc_hd__xnor2_2
XFILLER_0_174_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_263 _03728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19398_ _04168_ _04686_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__xor2_1
XINSDIODE1_274 _10660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_285 _11318_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_296 _12952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18349_ execute.io_mem_rd\[1\] decode.id_ex_ex_rs1_reg\[1\] VGND VGND VPWR VPWR _03648_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21360_ _06192_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20311_ _05355_ _05412_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21291_ net1425 _06153_ _06141_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__mux2_1
Xinput60 io_memory_read_data[4] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_1
XFILLER_0_31_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold800 decode.regfile.registers_20\[4\] VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 fetch.bht.bhtTable_tag\[2\]\[18\] VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23030_ _07076_ _07474_ _07084_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__a21o_1
Xhold822 _01131_ VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 fetch.bht.bhtTable_target_pc\[3\]\[18\] VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__dlygate4sd3_1
X_20242_ _05418_ _05259_ _05430_ _05431_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_114_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold844 fetch.bht.bhtTable_tag\[12\]\[8\] VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold855 fetch.bht.bhtTable_target_pc\[1\]\[10\] VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold866 csr._mcycle_T_2\[22\] VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold877 fetch.bht.bhtTable_target_pc\[4\]\[20\] VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 fetch.bht.bhtTable_target_pc\[14\]\[20\] VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20173_ decode.id_ex_imm_reg\[25\] _10790_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__nand2_1
Xhold899 decode.regfile.registers_6\[4\] VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2201 decode.regfile.registers_14\[29\] VGND VGND VPWR VPWR net2428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2212 decode.regfile.registers_10\[6\] VGND VGND VPWR VPWR net2439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2223 decode.regfile.registers_2\[20\] VGND VGND VPWR VPWR net2450 sky130_fd_sc_hd__dlygate4sd3_1
X_24981_ csr._mcycle_T_3\[63\] csr._mcycle_T_3\[62\] csr._mcycle_T_3\[61\] _08696_
+ _03579_ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__a41o_1
Xhold2234 decode.regfile.registers_7\[22\] VGND VGND VPWR VPWR net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1500 fetch.bht.bhtTable_target_pc\[7\]\[23\] VGND VGND VPWR VPWR net1727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2245 decode.regfile.registers_15\[14\] VGND VGND VPWR VPWR net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 fetch.bht.bhtTable_target_pc\[13\]\[14\] VGND VGND VPWR VPWR net1738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2256 csr._mcycle_T_2\[7\] VGND VGND VPWR VPWR net2483 sky130_fd_sc_hd__clkbuf_2
X_26720_ _09398_ _09720_ VGND VGND VPWR VPWR _09725_ sky130_fd_sc_hd__nand2_1
Xhold1522 fetch.bht.bhtTable_target_pc\[3\]\[25\] VGND VGND VPWR VPWR net1749 sky130_fd_sc_hd__dlygate4sd3_1
X_23932_ _08136_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__clkbuf_1
Xhold2267 decode.regfile.registers_4\[22\] VGND VGND VPWR VPWR net2494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 fetch.bht.bhtTable_tag\[11\]\[12\] VGND VGND VPWR VPWR net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2278 execute.io_reg_pc\[5\] VGND VGND VPWR VPWR net2505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1544 decode.regfile.registers_13\[19\] VGND VGND VPWR VPWR net1771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2289 decode.regfile.registers_7\[24\] VGND VGND VPWR VPWR net2516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 fetch.bht.bhtTable_tag\[9\]\[11\] VGND VGND VPWR VPWR net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1566 fetch.bht.bhtTable_tag\[14\]\[16\] VGND VGND VPWR VPWR net1793 sky130_fd_sc_hd__dlygate4sd3_1
X_26651_ net644 _09679_ _09684_ _09675_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__o211a_1
X_23863_ _08096_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__clkbuf_1
Xhold1577 fetch.bht.bhtTable_tag\[11\]\[21\] VGND VGND VPWR VPWR net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1588 fetch.bht.bhtTable_tag\[14\]\[13\] VGND VGND VPWR VPWR net1815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1599 fetch.bht.bhtTable_target_pc\[0\]\[9\] VGND VGND VPWR VPWR net1826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25602_ _10373_ _08903_ _09935_ _10196_ VGND VGND VPWR VPWR _09066_ sky130_fd_sc_hd__and4_1
X_22814_ _07302_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__clkbuf_1
X_29370_ clknet_leaf_255_clock _02383_ VGND VGND VPWR VPWR decode.regfile.registers_4\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_26582_ net738 _09636_ _09644_ _09635_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23794_ _08049_ net1422 _07952_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28321_ clknet_leaf_199_clock _01334_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25533_ _08982_ _09026_ VGND VGND VPWR VPWR _09028_ sky130_fd_sc_hd__nand2_1
X_22745_ _09901_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_183_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28252_ clknet_leaf_79_clock _01274_ VGND VGND VPWR VPWR csr._minstret_T_3\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22676_ net2633 _07222_ _07225_ _07221_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__o211a_1
X_25464_ _08916_ _08980_ VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27203_ clknet_leaf_363_clock _00232_ VGND VGND VPWR VPWR decode.regfile.registers_28\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_24415_ net1164 execute.io_target_pc\[30\] _09911_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__mux2_1
X_21627_ csr.minstret\[8\] _06346_ _06347_ _06331_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_192_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28183_ clknet_leaf_59_clock _01205_ VGND VGND VPWR VPWR csr.io_mret_vector\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25395_ _08939_ _08923_ VGND VGND VPWR VPWR _08940_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27134_ clknet_leaf_360_clock _00163_ VGND VGND VPWR VPWR decode.regfile.registers_26\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_24346_ _08349_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__clkbuf_1
X_21558_ _06299_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20509_ csr._minstret_T_3\[42\] _05578_ _05617_ csr._csr_read_data_T_8\[10\] _05559_
+ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24277_ _08105_ net1144 _06218_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27065_ clknet_leaf_345_clock _00094_ VGND VGND VPWR VPWR decode.regfile.registers_24\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_21489_ _06261_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__clkbuf_1
X_14030_ _10102_ _10268_ VGND VGND VPWR VPWR _10276_ sky130_fd_sc_hd__nand2_1
X_23228_ fetch.bht.bhtTable_target_pc\[8\]\[19\] fetch.bht.bhtTable_target_pc\[9\]\[19\]
+ _07067_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26016_ _08937_ _09297_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23159_ net280 _07596_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_224_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27967_ clknet_leaf_239_clock _00989_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ decode.regfile.registers_8\[17\] _11285_ _11287_ _11960_ VGND VGND VPWR VPWR
+ _11961_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_8_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29706_ clknet_leaf_282_clock _02719_ VGND VGND VPWR VPWR decode.regfile.registers_14\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17720_ decode.regfile.registers_7\[23\] _12612_ _12889_ VGND VGND VPWR VPWR _03124_
+ sky130_fd_sc_hd__a21oi_1
X_26918_ _09837_ VGND VGND VPWR VPWR _09838_ sky130_fd_sc_hd__clkbuf_4
X_14932_ _10960_ VGND VGND VPWR VPWR _10961_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27898_ clknet_leaf_69_clock _00927_ VGND VGND VPWR VPWR csr._mcycle_T_2\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_145_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17651_ decode.regfile.registers_18\[21\] _12572_ _12562_ _03056_ VGND VGND VPWR
+ VPWR _03057_ sky130_fd_sc_hd__a211o_1
X_29637_ clknet_leaf_276_clock _02650_ VGND VGND VPWR VPWR decode.regfile.registers_12\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14863_ decode.id_ex_pc_reg\[26\] _10769_ _10858_ _10860_ _10905_ VGND VGND VPWR
+ VPWR _10906_ sky130_fd_sc_hd__o311a_1
X_26849_ net2276 _09795_ _09798_ _09799_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16602_ _12559_ VGND VGND VPWR VPWR _12567_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_19_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ _10147_ _09937_ VGND VGND VPWR VPWR _10148_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17582_ _10939_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__clkbuf_2
X_29568_ clknet_leaf_312_clock _02581_ VGND VGND VPWR VPWR decode.regfile.registers_10\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14794_ _10832_ _10833_ _10835_ _10836_ VGND VGND VPWR VPWR _10837_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19321_ _04171_ _04173_ _04611_ _04590_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__or4_1
X_28519_ clknet_leaf_194_clock _01532_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_16533_ _12497_ VGND VGND VPWR VPWR _12498_ sky130_fd_sc_hd__clkbuf_4
X_13745_ _09943_ _09940_ memory.io_wb_reg_pc\[21\] VGND VGND VPWR VPWR _10089_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_80_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29499_ clknet_leaf_251_clock _02512_ VGND VGND VPWR VPWR decode.regfile.registers_8\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19252_ _04054_ _03971_ _04233_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16464_ decode.regfile.registers_10\[30\] _11509_ _12419_ _12430_ VGND VGND VPWR
+ VPWR _12431_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13676_ _10030_ VGND VGND VPWR VPWR _10031_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18203_ decode.control.io_funct3\[2\] _10943_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15415_ decode.regfile.registers_5\[3\] _10637_ _11139_ VGND VGND VPWR VPWR _11409_
+ sky130_fd_sc_hd__and3_1
X_19183_ _04255_ _04062_ _04324_ _04478_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_1344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16395_ _12348_ _12362_ _12363_ VGND VGND VPWR VPWR _12364_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18134_ _03495_ _03493_ _03487_ net2171 VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_170_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15346_ decode.regfile.registers_29\[1\] _11255_ _11256_ _11341_ _11246_ VGND VGND
+ VPWR VPWR _11342_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_113_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_322_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_322_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18065_ _10943_ _10941_ _10581_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_78_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15277_ _11272_ VGND VGND VPWR VPWR _11273_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_184_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17016_ decode.regfile.registers_8\[6\] _12889_ _12607_ VGND VGND VPWR VPWR _12975_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_229_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14228_ _10031_ _10387_ VGND VGND VPWR VPWR _10391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14159_ net631 _10346_ _10350_ _10344_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_337_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_337_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18967_ net190 _04253_ _04264_ _04265_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _12602_ decode.regfile.registers_9\[28\] _12653_ _03316_ VGND VGND VPWR VPWR
+ _03317_ sky130_fd_sc_hd__o211a_2
X_18898_ _03890_ decode.id_ex_imm_reg\[17\] _03906_ _03907_ _03934_ VGND VGND VPWR
+ VPWR _04197_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_217_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_19 _02192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17849_ decode.regfile.registers_21\[26\] _12682_ _03226_ _03249_ _12806_ VGND VGND
+ VPWR VPWR _03250_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_33_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20860_ _05907_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19519_ _04729_ _04797_ _04800_ _04803_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_102_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20791_ execute.io_mem_rd\[1\] _05867_ _05868_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_102_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22530_ fetch.bht.bhtTable_target_pc\[6\]\[1\] fetch.bht.bhtTable_target_pc\[7\]\[1\]
+ _07123_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22461_ fetch.btb.btbTable\[1\]\[1\] _06674_ fetch.bht.bhtTable_valid\[1\] _07055_
+ _00002_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__a311o_1
XFILLER_0_228_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24200_ _08274_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__clkbuf_1
X_21412_ _06103_ net1358 _06219_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25180_ _10573_ net2690 _08818_ VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22392_ _06684_ _06986_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24131_ net1104 execute.io_target_pc\[20\] _08232_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__mux2_1
X_21343_ _06182_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24062_ net1061 VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__clkbuf_1
X_21274_ _06142_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__clkbuf_1
Xhold630 _08202_ VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold641 fetch.bht.bhtTable_target_pc\[11\]\[30\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23013_ fetch.bht.bhtTable_target_pc\[12\]\[7\] fetch.bht.bhtTable_target_pc\[13\]\[7\]
+ _07439_ VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__mux2_1
Xhold652 fetch.bht.bhtTable_tag\[8\]\[0\] VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold663 fetch.bht.bhtTable_target_pc\[1\]\[9\] VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__dlygate4sd3_1
X_20225_ decode.id_ex_pc_reg\[1\] _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__or2_1
X_28870_ clknet_leaf_96_clock _01883_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold674 decode.regfile.registers_14\[11\] VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 fetch.bht.bhtTable_target_pc\[12\]\[12\] VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold696 csr._csr_read_data_T_8\[11\] VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__buf_1
XFILLER_0_228_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27821_ clknet_leaf_325_clock _00850_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_20156_ decode.id_ex_imm_reg\[21\] _10798_ _05357_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2020 decode.regfile.registers_9\[16\] VGND VGND VPWR VPWR net2247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2031 decode.regfile.registers_18\[0\] VGND VGND VPWR VPWR net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2042 execute.csr_write_enable_out_reg VGND VGND VPWR VPWR net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2053 decode.io_id_pc\[1\] VGND VGND VPWR VPWR net2280 sky130_fd_sc_hd__dlygate4sd3_1
X_27752_ clknet_leaf_323_clock _00781_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20087_ decode.id_ex_imm_reg\[13\] _10710_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__and2_1
X_24964_ csr._mcycle_T_3\[56\] csr._mcycle_T_3\[55\] _08685_ VGND VGND VPWR VPWR _08689_
+ sky130_fd_sc_hd__and3_1
Xhold2064 csr._minstret_T_3\[39\] VGND VGND VPWR VPWR net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1330 fetch.bht.bhtTable_tag\[3\]\[19\] VGND VGND VPWR VPWR net1557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2075 decode.regfile.registers_3\[26\] VGND VGND VPWR VPWR net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 fetch.bht.bhtTable_tag\[6\]\[16\] VGND VGND VPWR VPWR net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2086 decode.regfile.registers_24\[14\] VGND VGND VPWR VPWR net2313 sky130_fd_sc_hd__dlygate4sd3_1
X_26703_ _09381_ _09710_ VGND VGND VPWR VPWR _09715_ sky130_fd_sc_hd__nand2_1
X_23915_ _08127_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__clkbuf_1
Xhold1352 fetch.bht.bhtTable_target_pc\[7\]\[10\] VGND VGND VPWR VPWR net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2097 decode.regfile.registers_24\[4\] VGND VGND VPWR VPWR net2324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1363 csr.mscratch\[10\] VGND VGND VPWR VPWR net1590 sky130_fd_sc_hd__dlygate4sd3_1
X_27683_ clknet_leaf_30_clock _00712_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24895_ net341 _08643_ _03556_ csr.mcycle\[18\] VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__and4_1
Xhold1374 fetch.bht.bhtTable_target_pc\[0\]\[12\] VGND VGND VPWR VPWR net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1385 fetch.bht.bhtTable_target_pc\[9\]\[15\] VGND VGND VPWR VPWR net1612 sky130_fd_sc_hd__dlygate4sd3_1
X_29422_ clknet_leaf_262_clock _02435_ VGND VGND VPWR VPWR decode.regfile.registers_5\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1396 fetch.bht.bhtTable_tag\[8\]\[13\] VGND VGND VPWR VPWR net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26634_ _09566_ VGND VGND VPWR VPWR _09675_ sky130_fd_sc_hd__clkbuf_4
X_23846_ execute.io_target_pc\[17\] VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__buf_2
XFILLER_0_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29353_ clknet_leaf_228_clock _02366_ VGND VGND VPWR VPWR decode.regfile.registers_3\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26565_ net575 _09622_ _09634_ _09635_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__o211a_1
X_23777_ _08040_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__clkbuf_1
X_20989_ execute.io_reg_pc\[19\] _05977_ _05973_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__and3_1
XFILLER_0_200_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28304_ clknet_leaf_155_clock _01317_ VGND VGND VPWR VPWR decode.id_ex_aluop_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13530_ _09906_ VGND VGND VPWR VPWR _09907_ sky130_fd_sc_hd__buf_4
X_25516_ _08990_ VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22728_ _07256_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__clkbuf_1
X_29284_ clknet_leaf_231_clock _02297_ VGND VGND VPWR VPWR decode.regfile.registers_1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26496_ _09400_ _09589_ VGND VGND VPWR VPWR _09596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28235_ clknet_leaf_72_clock _01257_ VGND VGND VPWR VPWR csr._minstret_T_3\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_188_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25447_ _08975_ _08905_ VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_188_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22659_ net2702 _07208_ _07215_ _07164_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15200_ _11191_ _10624_ _11051_ VGND VGND VPWR VPWR _11197_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_213_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28166_ clknet_leaf_53_clock _01188_ VGND VGND VPWR VPWR csr.io_mret_vector\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16180_ decode.regfile.registers_14\[22\] _11208_ _12153_ _11199_ _12154_ VGND VGND
+ VPWR VPWR _12155_ sky130_fd_sc_hd__a221o_1
X_25378_ _08905_ VGND VGND VPWR VPWR _08928_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15131_ _11127_ VGND VGND VPWR VPWR _11128_ sky130_fd_sc_hd__clkbuf_4
X_27117_ clknet_leaf_329_clock _00146_ VGND VGND VPWR VPWR decode.regfile.registers_25\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_24329_ _08091_ net1184 _08334_ VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28097_ clknet_leaf_70_clock _01119_ VGND VGND VPWR VPWR csr.minstret\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27048_ clknet_leaf_346_clock _00077_ VGND VGND VPWR VPWR decode.regfile.registers_23\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15062_ _11058_ VGND VGND VPWR VPWR _11059_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14013_ _10064_ _10255_ VGND VGND VPWR VPWR _10266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19870_ _04392_ _05136_ _05139_ _04492_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18821_ _04116_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__nor2_2
X_28999_ clknet_leaf_111_clock _02012_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_207_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18752_ _04044_ _04049_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__and2_2
X_15964_ _11063_ VGND VGND VPWR VPWR _11944_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_216_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ _13221_ _03105_ _03106_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__a31o_1
X_14915_ _10945_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18683_ net202 _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__nand2_2
X_15895_ _11435_ decode.regfile.registers_22\[15\] _11450_ _10979_ _10991_ VGND VGND
+ VPWR VPWR _11877_ sky130_fd_sc_hd__o2111a_1
X_17634_ _03039_ _10602_ _10593_ _12522_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_177_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ csr.io_mem_pc\[5\] net287 VGND VGND VPWR VPWR _10889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_177_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17565_ _12874_ _02971_ _02972_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a21oi_1
X_14777_ csr.io_mem_pc\[6\] VGND VGND VPWR VPWR _10820_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19304_ _04324_ _04276_ net245 _04418_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__o211a_1
X_16516_ _11076_ decode.regfile.registers_27\[31\] _11257_ VGND VGND VPWR VPWR _12482_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13728_ _09937_ VGND VGND VPWR VPWR _10075_ sky130_fd_sc_hd__buf_2
X_17496_ _13407_ decode.regfile.registers_25\[17\] _13045_ _13294_ VGND VGND VPWR
+ VPWR _13444_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19235_ _04500_ _04464_ _04039_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16447_ _11445_ _12413_ _12414_ VGND VGND VPWR VPWR _12415_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13659_ _09937_ VGND VGND VPWR VPWR _10016_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_136_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19166_ _04373_ _04255_ _04231_ _04352_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_261_clock clknet_5_22__leaf_clock VGND VGND VPWR VPWR clknet_leaf_261_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16378_ decode.regfile.registers_15\[28\] _11036_ _11205_ _11202_ VGND VGND VPWR
+ VPWR _12347_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_76_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18117_ _03482_ _03480_ _03474_ decode.io_id_pc\[15\] VGND VGND VPWR VPWR _03486_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_83_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15329_ _11218_ VGND VGND VPWR VPWR _11325_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19097_ _03816_ _04000_ _04005_ _04001_ _03998_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_152_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18048_ _10929_ decode.regfile.registers_28\[31\] _12697_ VGND VGND VPWR VPWR _03444_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_276_clock clknet_5_21__leaf_clock VGND VGND VPWR VPWR clknet_leaf_276_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20010_ _04261_ decode.id_ex_pc_reg\[1\] _05234_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19999_ _05222_ _03587_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__nor2_4
XFILLER_0_158_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21961_ net1370 _06572_ _06582_ _06579_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23700_ _08000_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20912_ _05925_ _05933_ net41 VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__and3_1
X_24680_ _08523_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__clkbuf_1
X_21892_ _06533_ _06519_ _06520_ _06534_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_5_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_5_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_214_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_214_clock
+ sky130_fd_sc_hd__clkbuf_8
X_23631_ _07963_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__clkbuf_1
X_20843_ net108 _05891_ _05887_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26350_ _09406_ _09502_ VGND VGND VPWR VPWR _09511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23562_ _06795_ _07917_ _07925_ _05805_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__o211a_1
X_20774_ _10018_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25301_ _08881_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22513_ _07106_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__clkbuf_8
X_23493_ net25 _07875_ _07885_ _07879_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__o211a_1
X_26281_ net1697 _09462_ _09470_ _09471_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28020_ clknet_leaf_237_clock _01042_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25232_ _08845_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22444_ _06618_ fetch.btb.btbTable\[11\]\[1\] fetch.bht.bhtTable_valid\[11\] _07038_
+ _06631_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__a311o_1
XFILLER_0_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22375_ _06730_ _06969_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__and2b_1
XFILLER_0_190_998 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25163_ _10573_ net2760 _08809_ VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24114_ net1328 execute.io_target_pc\[12\] _08221_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__mux2_1
X_21326_ _06173_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__clkbuf_1
X_25094_ _06111_ net2102 _08596_ VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28922_ clknet_leaf_128_clock _01935_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24045_ _08194_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__clkbuf_1
X_21257_ net1234 _06130_ _06120_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__mux2_1
Xhold460 decode.regfile.registers_22\[14\] VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 decode.regfile.registers_29\[6\] VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap190 _03956_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
Xhold482 execute.csr_write_data_out_reg\[30\] VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20208_ decode.id_ex_imm_reg\[30\] decode.id_ex_pc_reg\[30\] VGND VGND VPWR VPWR
+ _05405_ sky130_fd_sc_hd__xor2_1
Xhold493 decode.regfile.registers_15\[12\] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28853_ clknet_leaf_114_clock _01866_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21188_ _06089_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27804_ clknet_leaf_328_clock _00833_ VGND VGND VPWR VPWR memory.io_wb_readdata\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_20139_ decode.id_ex_imm_reg\[17\] _10806_ _05334_ _05336_ VGND VGND VPWR VPWR _05346_
+ sky130_fd_sc_hd__o211ai_1
X_28784_ clknet_leaf_121_clock _01797_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_25996_ net2659 _09286_ _09294_ _09292_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27735_ clknet_leaf_38_clock _00764_ VGND VGND VPWR VPWR decode.id_ex_ex_use_rs2_reg
+ sky130_fd_sc_hd__dfxtp_1
X_24947_ csr._mcycle_T_3\[50\] csr._mcycle_T_3\[49\] _08674_ VGND VGND VPWR VPWR _08678_
+ sky130_fd_sc_hd__and3_1
Xhold1160 decode.regfile.registers_8\[5\] VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14700_ decode.id_ex_pc_reg\[28\] VGND VGND VPWR VPWR _10743_ sky130_fd_sc_hd__inv_2
Xhold1171 decode.regfile.registers_25\[16\] VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 fetch.bht.bhtTable_tag\[1\]\[11\] VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__dlygate4sd3_1
X_15680_ decode.regfile.registers_18\[9\] _10642_ _11112_ _10652_ _10633_ VGND VGND
+ VPWR VPWR _11668_ sky130_fd_sc_hd__o2111a_1
X_27666_ clknet_leaf_29_clock _00695_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_219_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24878_ csr.mcycle\[16\] csr.mcycle\[15\] _08626_ _08627_ VGND VGND VPWR VPWR _08628_
+ sky130_fd_sc_hd__and4_1
Xhold1193 decode.regfile.registers_19\[6\] VGND VGND VPWR VPWR net1420 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_219_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29405_ clknet_leaf_247_clock _02418_ VGND VGND VPWR VPWR decode.regfile.registers_5\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_219_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ execute.io_target_pc\[1\] VGND VGND VPWR VPWR _10674_ sky130_fd_sc_hd__inv_2
X_26617_ _09664_ VGND VGND VPWR VPWR _09665_ sky130_fd_sc_hd__buf_2
X_23829_ _08073_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27597_ clknet_leaf_153_clock _00626_ VGND VGND VPWR VPWR execute.io_target_pc\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_169_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29336_ clknet_leaf_243_clock _02349_ VGND VGND VPWR VPWR decode.regfile.registers_2\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17350_ _12708_ net409 _13261_ _13301_ _13219_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_215_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ decode.immGen._imm_T_24\[18\] VGND VGND VPWR VPWR _10605_ sky130_fd_sc_hd__clkinv_4
X_26548_ _09377_ _09623_ VGND VGND VPWR VPWR _09626_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_215_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16301_ _11646_ _11834_ _11944_ decode.regfile.registers_29\[25\] _12272_ VGND VGND
+ VPWR VPWR _12273_ sky130_fd_sc_hd__o221a_1
XFILLER_0_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13513_ _09881_ _09884_ _09885_ _09892_ net391 VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__a41o_1
X_29267_ clknet_leaf_224_clock _02280_ VGND VGND VPWR VPWR decode.regfile.registers_0\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_17281_ decode.regfile.registers_8\[12\] _12776_ _12549_ _12604_ _12606_ VGND VGND
+ VPWR VPWR _13234_ sky130_fd_sc_hd__a41o_1
XFILLER_0_222_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26479_ _09383_ _09579_ VGND VGND VPWR VPWR _09586_ sky130_fd_sc_hd__nand2_1
X_14493_ net518 _10533_ _10542_ _10535_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19020_ net314 _04307_ _04249_ _04318_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28218_ clknet_leaf_84_clock net2007 VGND VGND VPWR VPWR csr.mscratch\[20\] sky130_fd_sc_hd__dfxtp_1
X_16232_ decode.regfile.registers_14\[24\] _11207_ _11273_ decode.regfile.registers_15\[24\]
+ _11361_ VGND VGND VPWR VPWR _12205_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29198_ clknet_leaf_240_clock _02211_ VGND VGND VPWR VPWR fetch.btb.btbTable\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28149_ clknet_leaf_190_clock _01171_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16163_ decode.regfile.registers_1\[22\] VGND VGND VPWR VPWR _12138_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15114_ _11110_ VGND VGND VPWR VPWR _11111_ sky130_fd_sc_hd__buf_4
XFILLER_0_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16094_ _12069_ _12070_ VGND VGND VPWR VPWR _12071_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_71_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19922_ _03854_ _03862_ _05164_ _04496_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__o31ai_1
X_15045_ _11041_ VGND VGND VPWR VPWR _11042_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_166_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19853_ _03803_ _05123_ _04526_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18804_ _03889_ decode.id_ex_imm_reg\[13\] _04101_ _04102_ VGND VGND VPWR VPWR _04103_
+ sky130_fd_sc_hd__a22oi_4
X_16996_ _10927_ decode.regfile.registers_24\[5\] _10933_ _12759_ _12862_ VGND VGND
+ VPWR VPWR _12956_ sky130_fd_sc_hd__o2111a_1
X_19784_ _05044_ _05055_ _03835_ _05057_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_207_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15947_ decode.regfile.registers_14\[16\] _11360_ _11927_ _11198_ VGND VGND VPWR
+ VPWR _11928_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18735_ decode.id_ex_rs1_data_reg\[4\] _03687_ _04030_ _03699_ _04033_ VGND VGND
+ VPWR VPWR _04034_ sky130_fd_sc_hd__o221a_4
XTAP_TAPCELL_ROW_69_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18666_ _03888_ _03893_ _03872_ _03881_ _03964_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__o221a_1
X_15878_ decode.regfile.registers_19\[14\] _11354_ _11837_ _11860_ _11325_ VGND VGND
+ VPWR VPWR _11861_ sky130_fd_sc_hd__o221a_1
X_14829_ csr.io_mem_pc\[14\] VGND VGND VPWR VPWR _10872_ sky130_fd_sc_hd__clkbuf_8
X_17617_ _13339_ _03021_ _03022_ _03023_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18597_ execute.csr_read_data_out_reg\[19\] _03659_ net110 _03665_ _03895_ VGND VGND
+ VPWR VPWR _03896_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_138_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17548_ decode.regfile.registers_13\[19\] _12534_ _12589_ _12664_ VGND VGND VPWR
+ VPWR _13494_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17479_ _13425_ _13426_ VGND VGND VPWR VPWR _13427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19218_ _03638_ _04241_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20490_ csr.mcycle\[7\] _05552_ _05636_ _05642_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19149_ _04445_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_225_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22160_ fetch.bht.bhtTable_tag\[0\]\[13\] fetch.bht.bhtTable_tag\[1\]\[13\] fetch.bht.bhtTable_tag\[2\]\[13\]
+ fetch.bht.bhtTable_tag\[3\]\[13\] _06754_ _06622_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21111_ _06047_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_1253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22091_ _06626_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_160_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21042_ _06006_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout225 net71 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25850_ _09198_ VGND VGND VPWR VPWR _09210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24801_ _08587_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25781_ _08929_ _09166_ VGND VGND VPWR VPWR _09171_ sky130_fd_sc_hd__nand2_1
X_22993_ _07439_ fetch.bht.bhtTable_target_pc\[15\]\[6\] _07125_ VGND VGND VPWR VPWR
+ _07440_ sky130_fd_sc_hd__a21bo_1
X_27520_ clknet_leaf_54_clock _00549_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_4
X_24732_ _08550_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_153_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_153_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21944_ _06570_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27451_ clknet_leaf_149_clock _00480_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_24663_ net1035 execute.io_target_pc\[20\] _08508_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21875_ csr.io_mret_vector\[11\] _10812_ _06515_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__mux2_1
X_26402_ net697 _09534_ _09541_ _09540_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23614_ _07953_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__clkbuf_1
X_20826_ net131 _05879_ _05887_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__and3_1
X_27382_ clknet_leaf_15_clock _00411_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[23\]
+ sky130_fd_sc_hd__dfxtp_2
X_24594_ net1182 VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29121_ clknet_leaf_68_clock _02134_ VGND VGND VPWR VPWR csr.mcycle\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_168_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_168_clock
+ sky130_fd_sc_hd__clkbuf_8
X_26333_ net585 _09491_ _09501_ _09499_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23545_ net2236 _07904_ _07915_ VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__or3b_1
XFILLER_0_147_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20757_ _05847_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__buf_1
XFILLER_0_65_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29052_ clknet_leaf_181_clock _02065_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_210_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26264_ _09446_ VGND VGND VPWR VPWR _09462_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23476_ _10670_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__buf_2
X_20688_ _05801_ _05808_ net2588 _05810_ _00692_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__a32o_1
XFILLER_0_208_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28003_ clknet_leaf_194_clock _01025_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_25215_ _08836_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22427_ fetch.bht.bhtTable_tag\[6\]\[12\] fetch.bht.bhtTable_tag\[7\]\[12\] _06691_
+ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26195_ _09415_ _09413_ VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__nand2_1
X_25146_ net94 _07343_ _07344_ _07432_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__o31a_2
XFILLER_0_103_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22358_ fetch.bht.bhtTable_tag\[12\]\[14\] fetch.bht.bhtTable_tag\[13\]\[14\] fetch.bht.bhtTable_tag\[14\]\[14\]
+ fetch.bht.bhtTable_tag\[15\]\[14\] _06679_ _06620_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__mux4_1
X_21309_ _06164_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22289_ fetch.bht.bhtTable_tag\[12\]\[11\] fetch.bht.bhtTable_tag\[13\]\[11\] fetch.bht.bhtTable_tag\[14\]\[11\]
+ fetch.bht.bhtTable_tag\[15\]\[11\] _06674_ _06650_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__mux4_1
X_25077_ csr.mcycle\[28\] csr.mcycle\[27\] csr.mcycle\[29\] _08759_ VGND VGND VPWR
+ VPWR _08766_ sky130_fd_sc_hd__and4_1
XFILLER_0_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_208_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_106_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_106_clock
+ sky130_fd_sc_hd__clkbuf_8
X_24028_ _08185_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__clkbuf_1
X_28905_ clknet_leaf_88_clock _01918_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_208_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold290 decode.regfile.registers_29\[16\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
X_29885_ clknet_leaf_304_clock _02898_ VGND VGND VPWR VPWR decode.regfile.registers_20\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16850_ _10939_ decode.regfile.registers_25\[2\] _12506_ _12812_ VGND VGND VPWR VPWR
+ _12813_ sky130_fd_sc_hd__or4_1
X_28836_ clknet_leaf_130_clock _01849_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15801_ decode.regfile.registers_18\[12\] _11455_ _11784_ _11785_ _11456_ VGND VGND
+ VPWR VPWR _11786_ sky130_fd_sc_hd__a221o_1
X_28767_ clknet_leaf_180_clock _01780_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16781_ _12590_ VGND VGND VPWR VPWR _12745_ sky130_fd_sc_hd__clkbuf_4
X_13993_ net2286 _10243_ _10254_ _10249_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__o211a_1
X_25979_ net2603 _09243_ _09283_ _09277_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18520_ net119 _03666_ _03818_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15732_ _11251_ _11259_ decode.regfile.registers_27\[10\] _11686_ _11718_ VGND VGND
+ VPWR VPWR _11719_ sky130_fd_sc_hd__o32a_1
X_27718_ clknet_leaf_16_clock _00747_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28698_ clknet_leaf_177_clock _01711_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18451_ _03741_ execute.io_mem_rd\[2\] VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__nand2_1
X_27649_ clknet_leaf_49_clock _00678_ VGND VGND VPWR VPWR execute.io_reg_pc\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ decode.regfile.registers_7\[9\] _11465_ _11466_ decode.regfile.registers_6\[9\]
+ _11281_ VGND VGND VPWR VPWR _11651_ sky130_fd_sc_hd__a221o_1
XANTENNA_130 _10660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_141 csr._minstret_T_3\[42\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ decode.regfile.registers_10\[15\] _12790_ _13341_ _13351_ _12792_ VGND VGND
+ VPWR VPWR _13352_ sky130_fd_sc_hd__o221ai_2
XANTENNA_152 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14614_ _10655_ VGND VGND VPWR VPWR _10657_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_120_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ decode.io_wb_regwrite decode.id_ex_ex_use_rs1_reg VGND VGND VPWR VPWR _03681_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15594_ _11290_ _11582_ _11583_ VGND VGND VPWR VPWR _11584_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_200_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29319_ clknet_leaf_228_clock _02332_ VGND VGND VPWR VPWR decode.regfile.registers_2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_17333_ _13265_ _13284_ _12566_ VGND VGND VPWR VPWR _13285_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14545_ decode.immGen._imm_T_24\[17\] VGND VGND VPWR VPWR _10588_ sky130_fd_sc_hd__buf_4
XFILLER_0_166_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17264_ _13099_ _12768_ _13182_ decode.regfile.registers_29\[11\] _13217_ VGND VGND
+ VPWR VPWR _13218_ sky130_fd_sc_hd__o221a_1
X_14476_ _10505_ VGND VGND VPWR VPWR _10533_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19003_ _04297_ decode.id_ex_imm_reg\[4\] _04035_ _04298_ _04301_ VGND VGND VPWR
+ VPWR _04302_ sky130_fd_sc_hd__a221o_2
XFILLER_0_102_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16215_ decode.regfile.registers_16\[23\] _11359_ _12172_ _12188_ VGND VGND VPWR
+ VPWR _12189_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17195_ _13148_ _13149_ VGND VGND VPWR VPWR _13150_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_168_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16146_ decode.regfile.registers_18\[21\] _11455_ _12120_ _12121_ _11456_ VGND VGND
+ VPWR VPWR _12122_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_94_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16077_ _11942_ decode.regfile.registers_30\[20\] _11722_ _11723_ _11724_ VGND VGND
+ VPWR VPWR _12054_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_224_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15028_ _10994_ VGND VGND VPWR VPWR _11033_ sky130_fd_sc_hd__buf_4
X_19905_ _04425_ _05169_ _04794_ _04879_ _05173_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__a221o_1
XFILLER_0_220_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19836_ _05103_ _05104_ _05107_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__a21bo_1
Xhold1907 decode.regfile.registers_27\[18\] VGND VGND VPWR VPWR net2134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1918 fetch.bht.bhtTable_tag\[13\]\[5\] VGND VGND VPWR VPWR net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_70_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1929 csr._minstret_T_3\[52\] VGND VGND VPWR VPWR net2156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19767_ _04805_ _04654_ _04729_ _05041_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__a31o_1
X_16979_ _12936_ _12937_ _12938_ VGND VGND VPWR VPWR _12939_ sky130_fd_sc_hd__a21oi_1
Xinput3 net640 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_88_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18718_ net207 net206 net203 _09969_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__o211ai_4
X_19698_ _04974_ _04972_ _04957_ _04454_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18649_ _03944_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_85_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_85_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21660_ net2648 _06370_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20611_ _05588_ _05747_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__or2_2
XFILLER_0_4_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21591_ _06319_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__buf_2
XFILLER_0_117_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23330_ _07751_ _07757_ _07084_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__mux2_1
X_20542_ csr.minstret\[14\] _05572_ _05582_ csr.mcycle\[14\] _05687_ VGND VGND VPWR
+ VPWR _05688_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23261_ fetch.bht.bhtTable_target_pc\[4\]\[21\] fetch.bht.bhtTable_target_pc\[5\]\[21\]
+ _07106_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__mux2_1
X_20473_ _05627_ csr.io_mret_vector\[5\] _05603_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25000_ csr.mcycle\[4\] net1888 _08709_ _08713_ _06336_ VGND VGND VPWR VPWR _02133_
+ sky130_fd_sc_hd__a311oi_1
X_22212_ net90 _06806_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__xnor2_1
X_23192_ _06887_ _07613_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_23_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22143_ _06672_ _06731_ _06733_ _06737_ _06640_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__a311o_1
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22074_ _06661_ _06666_ _06633_ _06668_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_199_1151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26951_ net909 _09853_ _09857_ _09852_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1082 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25902_ _08975_ _09198_ VGND VGND VPWR VPWR _09239_ sky130_fd_sc_hd__nand2_1
X_21025_ execute.csr_read_data_out_reg\[3\] _05989_ _05985_ VGND VGND VPWR VPWR _05997_
+ sky130_fd_sc_hd__and3_1
X_29670_ clknet_leaf_281_clock _02683_ VGND VGND VPWR VPWR decode.regfile.registers_13\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26882_ net1743 _09809_ _09817_ _09812_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_38_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_38_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28621_ clknet_leaf_101_clock _01634_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25833_ _09025_ _09200_ VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28552_ clknet_leaf_214_clock _01565_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25764_ _08912_ _09157_ VGND VGND VPWR VPWR _09161_ sky130_fd_sc_hd__nand2_1
X_22976_ fetch.bht.bhtTable_target_pc\[12\]\[5\] fetch.bht.bhtTable_target_pc\[13\]\[5\]
+ fetch.bht.bhtTable_target_pc\[14\]\[5\] fetch.bht.bhtTable_target_pc\[15\]\[5\]
+ _07068_ _07110_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_195_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27503_ clknet_leaf_30_clock _00532_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dfxtp_1
X_24715_ _08541_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_195_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21927_ csr.io_mret_vector\[27\] _10759_ _06539_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__mux2_1
X_28483_ clknet_leaf_208_clock _01496_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_25695_ net2572 _09111_ _09120_ _09115_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27434_ clknet_leaf_54_clock _00463_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_191_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24646_ net912 execute.io_target_pc\[12\] _08497_ VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__mux2_1
X_21858_ _06509_ _06494_ _06495_ _06510_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20809_ net111 _05879_ _05875_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__and3_1
X_27365_ clknet_leaf_27_clock _00394_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24577_ _08470_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21789_ csr.io_csr_write_address\[1\] _06315_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__nor2_4
X_29104_ clknet_leaf_17_clock _02117_ VGND VGND VPWR VPWR csr._mcycle_T_3\[52\] sky130_fd_sc_hd__dfxtp_1
X_14330_ net1000 _10447_ _10449_ _10440_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__o211a_1
X_26316_ _09490_ VGND VGND VPWR VPWR _09492_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23528_ _04459_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_154_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27296_ clknet_leaf_1_clock _00325_ VGND VGND VPWR VPWR decode.regfile.registers_31\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29035_ clknet_leaf_93_clock _02048_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14261_ _10112_ _10400_ VGND VGND VPWR VPWR _10409_ sky130_fd_sc_hd__nand2_1
X_26247_ net609 _09447_ _09452_ _09440_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__o211a_1
X_23459_ net8 _07861_ _07866_ _07865_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_150_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16000_ _11756_ decode.regfile.registers_28\[17\] _11871_ _11681_ _11440_ VGND VGND
+ VPWR VPWR _11980_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_180_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14192_ _10290_ VGND VGND VPWR VPWR _10369_ sky130_fd_sc_hd__clkbuf_4
X_26178_ _10052_ VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25129_ _06147_ net1526 _08562_ VGND VGND VPWR VPWR _08793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29937_ clknet_leaf_340_clock _02950_ VGND VGND VPWR VPWR decode.regfile.registers_21\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_17951_ decode.regfile.registers_7\[29\] _12611_ _12889_ VGND VGND VPWR VPWR _03349_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16902_ _12516_ _12860_ _12861_ _12863_ VGND VGND VPWR VPWR _12864_ sky130_fd_sc_hd__a31o_1
X_17882_ decode.regfile.registers_13\[27\] _12533_ _12582_ _12662_ VGND VGND VPWR
+ VPWR _03282_ sky130_fd_sc_hd__a31o_1
X_29868_ clknet_leaf_300_clock _02881_ VGND VGND VPWR VPWR decode.regfile.registers_19\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19621_ _04509_ _04428_ _04898_ _04901_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__a31o_1
X_28819_ clknet_leaf_140_clock _01832_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_16833_ _11020_ _12490_ _12512_ decode.regfile.registers_12\[2\] _12591_ VGND VGND
+ VPWR VPWR _12796_ sky130_fd_sc_hd__o32a_1
X_29799_ clknet_leaf_297_clock _02812_ VGND VGND VPWR VPWR decode.regfile.registers_17\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16764_ _12557_ _10591_ _10607_ VGND VGND VPWR VPWR _12728_ sky130_fd_sc_hd__and3_1
X_19552_ _04740_ _04120_ _04834_ _04107_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__nand4_2
X_13976_ _09949_ VGND VGND VPWR VPWR _10245_ sky130_fd_sc_hd__buf_4
XFILLER_0_219_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15715_ decode.regfile.registers_9\[10\] _11547_ _10638_ _11132_ VGND VGND VPWR VPWR
+ _11702_ sky130_fd_sc_hd__o2bb2a_1
X_18503_ _03795_ _03800_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__nand2_2
XFILLER_0_220_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16695_ decode.regfile.registers_12\[0\] _12591_ _12596_ _12656_ _12659_ VGND VGND
+ VPWR VPWR _12660_ sky130_fd_sc_hd__o221a_1
X_19483_ _04768_ _04704_ _04352_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15646_ _11613_ _11633_ _11634_ VGND VGND VPWR VPWR _11635_ sky130_fd_sc_hd__o21ai_1
X_18434_ csr.io_csr_address\[0\] decode.io_wb_rd\[0\] VGND VGND VPWR VPWR _03733_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18365_ _03663_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__clkbuf_4
X_15577_ _10960_ decode.regfile.registers_28\[6\] _11067_ _11038_ _11440_ VGND VGND
+ VPWR VPWR _11568_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_113_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17316_ decode.regfile.registers_3\[13\] _10616_ _12729_ _12838_ VGND VGND VPWR VPWR
+ _13268_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14528_ _10565_ _10564_ _10571_ VGND VGND VPWR VPWR _10572_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18296_ decode.id_ex_rs2_data_reg\[14\] _03605_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17247_ decode.regfile.registers_12\[11\] _12591_ _13189_ _13200_ _12659_ VGND VGND
+ VPWR VPWR _13201_ sky130_fd_sc_hd__o221a_1
X_14459_ _10042_ _10517_ VGND VGND VPWR VPWR _10524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17178_ _13091_ _12706_ decode.regfile.registers_27\[9\] _13050_ VGND VGND VPWR VPWR
+ _13134_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16129_ decode.regfile.registers_1\[21\] _11539_ _12104_ VGND VGND VPWR VPWR _12105_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2405 csr._csr_read_data_T_8\[30\] VGND VGND VPWR VPWR net2632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2416 csr.mcycle\[11\] VGND VGND VPWR VPWR net2643 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2427 csr._csr_read_data_T_8\[4\] VGND VGND VPWR VPWR net2654 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2438 decode.regfile.registers_11\[19\] VGND VGND VPWR VPWR net2665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1704 fetch.bht.bhtTable_target_pc\[14\]\[10\] VGND VGND VPWR VPWR net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2449 csr._mcycle_T_2\[6\] VGND VGND VPWR VPWR net2676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1715 fetch.bht.bhtTable_target_pc\[10\]\[0\] VGND VGND VPWR VPWR net1942 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19819_ net188 _03812_ _04254_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__mux2_1
Xhold1726 decode.regfile.registers_20\[22\] VGND VGND VPWR VPWR net1953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1737 fetch.bht.bhtTable_tag\[13\]\[23\] VGND VGND VPWR VPWR net1964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1748 fetch.bht.bhtTable_tag\[7\]\[21\] VGND VGND VPWR VPWR net1975 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1759 fetch.bht.bhtTable_target_pc\[14\]\[7\] VGND VGND VPWR VPWR net1986 sky130_fd_sc_hd__dlygate4sd3_1
X_22830_ net1274 _10771_ _07308_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22761_ _07273_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24500_ _08060_ net1803 _08428_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21712_ csr.minstret\[27\] _06410_ _06317_ _06412_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_49_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25480_ _08931_ _08992_ VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22692_ _06578_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_192_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24431_ _08394_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21643_ net2444 _06358_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27150_ clknet_leaf_351_clock _00179_ VGND VGND VPWR VPWR decode.regfile.registers_26\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_24362_ net1628 execute.io_target_pc\[4\] _08356_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21574_ _06145_ net1904 _06306_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_30 _08939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26101_ net1836 _09343_ _09354_ _09346_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__o211a_1
XANTENNA_52 _10598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23313_ _07740_ _07063_ _07741_ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_63 _10935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20525_ _03721_ csr.io_mret_vector\[12\] _05565_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__o21a_1
X_27081_ clknet_leaf_347_clock _00110_ VGND VGND VPWR VPWR decode.regfile.registers_24\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24293_ _08055_ net1319 _06210_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__mux2_1
XANTENNA_74 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _12559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_96 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26032_ _08954_ _09310_ VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__nand2_1
X_23244_ net79 _07651_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__nand2_1
X_20456_ net1569 _05592_ _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23175_ net73 _07582_ net74 VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__a21oi_1
X_20387_ _05439_ _05201_ net455 VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__and3b_1
XFILLER_0_113_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_205_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22126_ fetch.bht.bhtTable_tag\[10\]\[4\] fetch.bht.bhtTable_tag\[11\]\[4\] _06680_
+ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__mux2_1
X_27983_ clknet_leaf_167_clock _01005_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26934_ net679 _09839_ _09847_ _09836_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__o211a_1
X_29722_ clknet_leaf_289_clock _02735_ VGND VGND VPWR VPWR decode.regfile.registers_15\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_201_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22057_ _06651_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_201_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21008_ execute.io_reg_pc\[28\] _05977_ _05985_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_197_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29653_ clknet_leaf_281_clock _02666_ VGND VGND VPWR VPWR decode.regfile.registers_12\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_26865_ _09392_ _09806_ VGND VGND VPWR VPWR _09808_ sky130_fd_sc_hd__nand2_1
X_28604_ clknet_leaf_181_clock _01617_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13830_ _09984_ _10154_ VGND VGND VPWR VPWR _10159_ sky130_fd_sc_hd__nand2_1
X_25816_ _08964_ _09179_ VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29584_ clknet_leaf_274_clock _02597_ VGND VGND VPWR VPWR decode.regfile.registers_10\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26796_ net520 _09766_ _09768_ _09758_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_3_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28535_ clknet_leaf_215_clock _01548_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13761_ _10102_ _10075_ VGND VGND VPWR VPWR _10103_ sky130_fd_sc_hd__nand2_1
X_25747_ _08970_ _09110_ VGND VGND VPWR VPWR _09150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22959_ fetch.bht.bhtTable_target_pc\[4\]\[4\] fetch.bht.bhtTable_target_pc\[5\]\[4\]
+ fetch.bht.bhtTable_target_pc\[6\]\[4\] fetch.bht.bhtTable_target_pc\[7\]\[4\] _07407_
+ _07115_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15500_ _10962_ decode.regfile.registers_30\[5\] _11039_ _11032_ _11033_ VGND VGND
+ VPWR VPWR _11492_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28466_ clknet_leaf_138_clock _01479_ VGND VGND VPWR VPWR decode.io_id_pc\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_156_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16480_ _11076_ decode.regfile.registers_27\[30\] _11869_ VGND VGND VPWR VPWR _12447_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_195_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13692_ _09977_ _09978_ memory.io_wb_reg_pc\[13\] VGND VGND VPWR VPWR _10044_ sky130_fd_sc_hd__o21ai_2
X_25678_ _09109_ VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15431_ _11124_ decode.regfile.registers_16\[3\] _11127_ _11424_ VGND VGND VPWR VPWR
+ _11425_ sky130_fd_sc_hd__o211a_1
X_27417_ clknet_leaf_15_clock _00446_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[26\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24629_ _07284_ VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_14_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28397_ clknet_leaf_143_clock _01410_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_14_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18150_ _03504_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_152_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27348_ clknet_leaf_45_clock _00377_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[21\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15362_ _11356_ VGND VGND VPWR VPWR _11357_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17101_ decode.regfile.registers_1\[8\] _12636_ _12531_ VGND VGND VPWR VPWR _13058_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_81_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14313_ _10426_ VGND VGND VPWR VPWR _10440_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18081_ _10915_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__buf_2
XFILLER_0_81_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27279_ clknet_leaf_328_clock _00308_ VGND VGND VPWR VPWR decode.regfile.registers_31\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_15293_ _11288_ VGND VGND VPWR VPWR _11289_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29018_ clknet_leaf_129_clock _02031_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_17032_ decode.regfile.registers_19\[6\] _10599_ _10589_ _12518_ _12544_ VGND VGND
+ VPWR VPWR _12991_ sky130_fd_sc_hd__o41a_1
XFILLER_0_180_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14244_ net652 _10390_ _10399_ _10398_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14175_ _10087_ _10355_ VGND VGND VPWR VPWR _10360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18983_ _04019_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_182_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17934_ _10929_ decode.regfile.registers_28\[28\] _02992_ VGND VGND VPWR VPWR _03333_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_175_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17865_ decode.regfile.registers_17\[27\] _11021_ _12559_ _12534_ VGND VGND VPWR
+ VPWR _03265_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19604_ _03911_ _03935_ _04865_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__o21a_1
X_16816_ _12531_ _10592_ _12558_ decode.regfile.registers_0\[2\] VGND VGND VPWR VPWR
+ _12779_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_85_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17796_ decode.regfile.registers_8\[25\] _12889_ _12607_ VGND VGND VPWR VPWR _03198_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_85_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19535_ _04081_ _04085_ _04786_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_191_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_187_Right_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13959_ _10117_ _10223_ VGND VGND VPWR VPWR _10234_ sky130_fd_sc_hd__nand2_1
X_16747_ _10930_ decode.regfile.registers_28\[1\] _12698_ VGND VGND VPWR VPWR _12711_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19466_ _04291_ _04535_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__or2_1
X_16678_ decode.regfile.registers_6\[0\] _10603_ _12615_ _12624_ _12642_ VGND VGND
+ VPWR VPWR _12643_ sky130_fd_sc_hd__o32a_1
XFILLER_0_9_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_220 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_231 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_242 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18417_ execute.io_mem_rd\[2\] csr.io_csr_address\[2\] VGND VGND VPWR VPWR _03716_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15629_ decode.regfile.registers_3\[8\] _11614_ _11367_ _10636_ VGND VGND VPWR VPWR
+ _11618_ sky130_fd_sc_hd__o2bb2a_1
XINSDIODE1_253 net200 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_264 _04982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19397_ _04645_ _04144_ _04670_ _04659_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__o211ai_1
XINSDIODE1_275 _10662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_286 _11381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_297 _13399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18348_ decode.id_ex_ex_rs1_reg\[1\] execute.io_mem_rd\[1\] VGND VGND VPWR VPWR _03647_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_228_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18279_ decode.id_ex_rs2_data_reg\[6\] _03596_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20310_ _05411_ _05482_ _05483_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__or3b_1
X_21290_ csr.io_mem_pc\[31\] VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__buf_2
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput50 io_memory_read_data[24] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 io_memory_read_data[5] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
Xhold801 fetch.bht.bhtTable_target_pc\[1\]\[18\] VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold812 fetch.bht.bhtTable_tag\[2\]\[6\] VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold823 fetch.bht.bhtTable_tag\[3\]\[25\] VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__dlygate4sd3_1
X_20241_ _10704_ _05427_ _05416_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold834 _08203_ VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold845 fetch.bht.bhtTable_target_pc\[1\]\[22\] VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold856 fetch.bht.bhtTable_target_pc\[1\]\[3\] VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold867 _01242_ VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 _08239_ VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20172_ decode.id_ex_imm_reg\[25\] _10790_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__or2_1
Xhold889 decode.regfile.registers_16\[4\] VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2202 decode.regfile.registers_5\[1\] VGND VGND VPWR VPWR net2429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24980_ _06331_ _08698_ _08699_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__nor3_1
Xhold2213 decode.regfile.registers_16\[5\] VGND VGND VPWR VPWR net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2224 decode.regfile.registers_19\[24\] VGND VGND VPWR VPWR net2451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2235 decode.regfile.registers_19\[27\] VGND VGND VPWR VPWR net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1501 fetch.bht.bhtTable_target_pc\[13\]\[0\] VGND VGND VPWR VPWR net1728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2246 fetch.bht.bhtTable_target_pc\[0\]\[30\] VGND VGND VPWR VPWR net2473 sky130_fd_sc_hd__dlygate4sd3_1
X_23931_ net1180 _08089_ _08130_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__mux2_1
Xhold1512 fetch.bht.bhtTable_tag\[12\]\[3\] VGND VGND VPWR VPWR net1739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2257 decode.regfile.registers_16\[30\] VGND VGND VPWR VPWR net2484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1523 fetch.bht.bhtTable_tag\[5\]\[23\] VGND VGND VPWR VPWR net1750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2268 decode.regfile.registers_18\[4\] VGND VGND VPWR VPWR net2495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1534 decode.regfile.registers_1\[17\] VGND VGND VPWR VPWR net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2279 decode.regfile.registers_7\[23\] VGND VGND VPWR VPWR net2506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1545 fetch.bht.bhtTable_target_pc\[13\]\[16\] VGND VGND VPWR VPWR net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 fetch.bht.bhtTable_target_pc\[6\]\[16\] VGND VGND VPWR VPWR net1783 sky130_fd_sc_hd__dlygate4sd3_1
X_26650_ _09404_ _09676_ VGND VGND VPWR VPWR _09684_ sky130_fd_sc_hd__nand2_1
Xhold1567 fetch.bht.bhtTable_target_pc\[10\]\[29\] VGND VGND VPWR VPWR net1794 sky130_fd_sc_hd__dlygate4sd3_1
X_23862_ _08095_ net1211 _08079_ VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__mux2_1
Xhold1578 fetch.bht.bhtTable_tag\[13\]\[24\] VGND VGND VPWR VPWR net1805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1589 fetch.bht.bhtTable_target_pc\[14\]\[8\] VGND VGND VPWR VPWR net1816 sky130_fd_sc_hd__dlygate4sd3_1
X_25601_ net717 _09026_ _09065_ _09059_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22813_ net2320 _10795_ _07297_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26581_ _09410_ _09632_ VGND VGND VPWR VPWR _09644_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23793_ execute.io_target_pc\[0\] VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28320_ clknet_leaf_193_clock _01333_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25532_ net637 _09024_ _09027_ _09017_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__o211a_1
X_22744_ _07264_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28251_ clknet_leaf_79_clock _01273_ VGND VGND VPWR VPWR csr._minstret_T_3\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_25463_ net2128 _08979_ _08986_ _08972_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22675_ net881 _07223_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27202_ clknet_leaf_363_clock _00231_ VGND VGND VPWR VPWR decode.regfile.registers_28\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_24414_ _08384_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28182_ clknet_leaf_59_clock _01204_ VGND VGND VPWR VPWR csr.io_mret_vector\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_21626_ net2436 _06329_ _06346_ csr.minstret\[8\] VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_75_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_205_Left_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25394_ _10057_ VGND VGND VPWR VPWR _08939_ sky130_fd_sc_hd__buf_6
XFILLER_0_69_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27133_ clknet_leaf_357_clock _00162_ VGND VGND VPWR VPWR decode.regfile.registers_26\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_24345_ _08107_ net2161 _06187_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21557_ _06128_ net1823 _06295_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20508_ _05534_ _05562_ _05536_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__or3b_4
XFILLER_0_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27064_ clknet_leaf_350_clock _00093_ VGND VGND VPWR VPWR decode.regfile.registers_24\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_24276_ _08313_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__clkbuf_1
X_21488_ _06117_ net1675 _06252_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26015_ net1298 _09300_ _09304_ _09305_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23227_ _07660_ _07071_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20439_ csr.minstret\[2\] _05594_ _05595_ csr._minstret_T_3\[34\] _05596_ VGND VGND
+ VPWR VPWR _05597_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23158_ _07592_ _07593_ _07594_ _07595_ _07371_ _07127_ VGND VGND VPWR VPWR _07596_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_224_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22109_ _06701_ _06623_ _06673_ _06703_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_224_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15980_ _11950_ _11959_ _11284_ VGND VGND VPWR VPWR _11960_ sky130_fd_sc_hd__nand3b_1
XPHY_EDGE_ROW_214_Left_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23089_ net69 _07504_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__nor2_1
X_27966_ clknet_leaf_218_clock _00988_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29705_ clknet_leaf_282_clock _02718_ VGND VGND VPWR VPWR decode.regfile.registers_14\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14931_ _10959_ VGND VGND VPWR VPWR _10960_ sky130_fd_sc_hd__clkbuf_4
X_26917_ net331 _10240_ _09935_ _10149_ VGND VGND VPWR VPWR _09837_ sky130_fd_sc_hd__and4_1
XFILLER_0_175_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27897_ clknet_leaf_19_clock _00926_ VGND VGND VPWR VPWR csr._mcycle_T_2\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_76_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14862_ decode.id_ex_pc_reg\[24\] _10861_ _10862_ _10904_ VGND VGND VPWR VPWR _10905_
+ sky130_fd_sc_hd__o211a_1
X_17650_ _12901_ _03054_ _03055_ _12826_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__o211a_1
X_29636_ clknet_leaf_276_clock _02649_ VGND VGND VPWR VPWR decode.regfile.registers_12\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_26848_ _09701_ VGND VGND VPWR VPWR _09799_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16601_ _12565_ VGND VGND VPWR VPWR _12566_ sky130_fd_sc_hd__clkbuf_4
X_13813_ _10146_ VGND VGND VPWR VPWR _10147_ sky130_fd_sc_hd__buf_4
X_17581_ _13183_ _02984_ _02985_ _02988_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__a31o_1
X_14793_ csr.io_mem_pc\[2\] _10834_ VGND VGND VPWR VPWR _10836_ sky130_fd_sc_hd__or2_1
X_26779_ _09381_ _09753_ VGND VGND VPWR VPWR _09759_ sky130_fd_sc_hd__nand2_1
X_29567_ clknet_leaf_252_clock _02580_ VGND VGND VPWR VPWR decode.regfile.registers_10\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16532_ _11016_ VGND VGND VPWR VPWR _12497_ sky130_fd_sc_hd__clkbuf_4
X_19320_ _04171_ _04173_ _04611_ _04590_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__o22ai_4
X_28518_ clknet_leaf_187_clock _01531_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_13744_ net2660 _10083_ _10088_ _10077_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29498_ clknet_leaf_252_clock _02511_ VGND VGND VPWR VPWR decode.regfile.registers_8\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19251_ _04409_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16463_ _12420_ _12428_ _12429_ VGND VGND VPWR VPWR _12430_ sky130_fd_sc_hd__o21a_1
X_28449_ clknet_leaf_144_clock _01462_ VGND VGND VPWR VPWR decode.io_id_pc\[7\] sky130_fd_sc_hd__dfxtp_1
X_13675_ memory.csr_read_data_out_reg\[10\] _09988_ _10028_ _10029_ VGND VGND VPWR
+ VPWR _10030_ sky130_fd_sc_hd__o22ai_4
XPHY_EDGE_ROW_223_Left_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18202_ _03535_ _03536_ _03537_ _03539_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15414_ decode.regfile.registers_7\[3\] _11378_ _11170_ decode.regfile.registers_6\[3\]
+ _11134_ VGND VGND VPWR VPWR _11408_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_117_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19182_ _04230_ _04126_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__or2_1
X_16394_ decode.regfile.registers_14\[28\] _11047_ _11053_ _11318_ VGND VGND VPWR
+ VPWR _12363_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18133_ _10575_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__buf_2
XFILLER_0_143_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15345_ _11250_ decode.regfile.registers_27\[1\] _11259_ _11238_ _11340_ VGND VGND
+ VPWR VPWR _11341_ sky130_fd_sc_hd__o311a_1
XFILLER_0_171_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18064_ _03454_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15276_ _10660_ _10655_ _11167_ VGND VGND VPWR VPWR _11272_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_78_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17015_ decode.regfile.registers_7\[6\] _12612_ _12623_ decode.regfile.registers_6\[6\]
+ _12973_ VGND VGND VPWR VPWR _12974_ sky130_fd_sc_hd__a221oi_2
XTAP_TAPCELL_ROW_184_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14227_ _10375_ VGND VGND VPWR VPWR _10390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_1075 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14158_ _10048_ _10342_ VGND VGND VPWR VPWR _10350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14089_ _10064_ _10299_ VGND VGND VPWR VPWR _10310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18966_ _03986_ _03985_ _03984_ _03987_ _03944_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__a311o_2
XFILLER_0_225_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _12726_ _03314_ _03315_ _12606_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_143_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18897_ _04190_ _04193_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__and3_1
XFILLER_0_206_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17848_ decode.regfile.registers_19\[26\] _12679_ _03227_ _03248_ _12545_ VGND VGND
+ VPWR VPWR _03249_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_33_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17779_ _10929_ decode.regfile.registers_28\[24\] _02992_ VGND VGND VPWR VPWR _03182_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19518_ _04386_ _04360_ _04799_ _04294_ _04802_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20790_ _05869_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19449_ _04735_ _04550_ _04409_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22460_ _06809_ fetch.bht.bhtTable_valid\[0\] fetch.btb.btbTable\[0\]\[1\] VGND VGND
+ VPWR VPWR _07055_ sky130_fd_sc_hd__and3b_1
XFILLER_0_147_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_228_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21411_ _06220_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22391_ fetch.bht.bhtTable_tag\[12\]\[9\] fetch.bht.bhtTable_tag\[13\]\[9\] _06706_
+ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24130_ _08238_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21342_ net1108 _10771_ _06179_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24061_ net1060 execute.io_target_pc\[18\] _08198_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__mux2_1
X_21273_ net1200 _06140_ _06141_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold620 decode.regfile.registers_4\[5\] VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 fetch.bht.bhtTable_target_pc\[11\]\[28\] VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold642 fetch.bht.bhtTable_target_pc\[0\]\[1\] VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlygate4sd3_1
X_23012_ _07439_ fetch.bht.bhtTable_target_pc\[14\]\[7\] VGND VGND VPWR VPWR _07458_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold653 decode.regfile.registers_29\[20\] VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20224_ decode.id_ex_rdsel_reg VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold664 decode.regfile.registers_29\[27\] VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold675 decode.regfile.registers_27\[17\] VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 fetch.bht.bhtTable_target_pc\[4\]\[1\] VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _05670_ VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_223_Right_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_217_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20155_ decode.id_ex_imm_reg\[20\] _10867_ _10798_ decode.id_ex_imm_reg\[21\] VGND
+ VGND VPWR VPWR _05360_ sky130_fd_sc_hd__a22oi_2
X_27820_ clknet_leaf_321_clock _00849_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2010 decode.regfile.registers_7\[17\] VGND VGND VPWR VPWR net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2021 decode.regfile.registers_16\[23\] VGND VGND VPWR VPWR net2248 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2032 decode.regfile.registers_16\[31\] VGND VGND VPWR VPWR net2259 sky130_fd_sc_hd__dlygate4sd3_1
X_20086_ _00560_ _05227_ _05300_ _05267_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__a2bb2oi_1
X_27751_ clknet_leaf_323_clock _00780_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2043 decode.regfile.registers_15\[4\] VGND VGND VPWR VPWR net2270 sky130_fd_sc_hd__dlygate4sd3_1
X_24963_ net940 _08687_ _08688_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__o21ba_1
Xhold2054 decode.regfile.registers_22\[31\] VGND VGND VPWR VPWR net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2065 fetch.bht.bhtTable_tag\[11\]\[17\] VGND VGND VPWR VPWR net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1320 fetch.bht.bhtTable_tag\[2\]\[1\] VGND VGND VPWR VPWR net1547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1331 decode.regfile.registers_2\[1\] VGND VGND VPWR VPWR net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2076 fetch.bht.bhtTable_tag\[0\]\[22\] VGND VGND VPWR VPWR net2303 sky130_fd_sc_hd__dlygate4sd3_1
X_23914_ net1156 _08072_ _08119_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__mux2_1
X_26702_ net2295 _09709_ _09714_ _09702_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__o211a_1
Xhold1342 csr.mscratch\[4\] VGND VGND VPWR VPWR net1569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2087 csr._mcycle_T_3\[47\] VGND VGND VPWR VPWR net2314 sky130_fd_sc_hd__dlygate4sd3_1
X_27682_ clknet_leaf_21_clock _00711_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_24894_ csr.mcycle\[11\] _03559_ _08642_ VGND VGND VPWR VPWR _08643_ sky130_fd_sc_hd__and3_1
Xhold1353 decode.regfile.registers_4\[30\] VGND VGND VPWR VPWR net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2098 decode.regfile.registers_14\[5\] VGND VGND VPWR VPWR net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 _01230_ VGND VGND VPWR VPWR net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 fetch.bht.bhtTable_tag\[0\]\[4\] VGND VGND VPWR VPWR net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 fetch.bht.bhtTable_target_pc\[10\]\[10\] VGND VGND VPWR VPWR net1613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26633_ _09387_ _09666_ VGND VGND VPWR VPWR _09674_ sky130_fd_sc_hd__nand2_1
X_29421_ clknet_leaf_260_clock _02434_ VGND VGND VPWR VPWR decode.regfile.registers_5\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23845_ _08084_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1397 fetch.bht.bhtTable_tag\[3\]\[20\] VGND VGND VPWR VPWR net1624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29352_ clknet_leaf_258_clock _02365_ VGND VGND VPWR VPWR decode.regfile.registers_3\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_26564_ _09566_ VGND VGND VPWR VPWR _09635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23776_ _06138_ net1873 _08030_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20988_ _05866_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__buf_2
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25515_ _08966_ _09005_ VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__nand2_1
X_28303_ clknet_leaf_45_clock net172 VGND VGND VPWR VPWR decode.id_ex_aluop_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_71_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22727_ _06101_ net1196 _09903_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__mux2_1
X_29283_ clknet_leaf_241_clock _02296_ VGND VGND VPWR VPWR decode.regfile.registers_1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_26495_ net939 _09592_ _09594_ _09595_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28234_ clknet_leaf_72_clock _01256_ VGND VGND VPWR VPWR csr._minstret_T_3\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_25446_ _10146_ VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_188_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22658_ net777 _07210_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_188_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_213_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21609_ _06323_ _06333_ net2705 _06331_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__a211oi_1
X_28165_ clknet_leaf_67_clock _01187_ VGND VGND VPWR VPWR csr._csr_read_data_T_9\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25377_ net1397 _08906_ _08926_ _08927_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_170_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22589_ csr._minstret_T_3\[44\] _07168_ _07169_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone53 net281 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__buf_4
XFILLER_0_106_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27116_ clknet_leaf_347_clock _00145_ VGND VGND VPWR VPWR decode.regfile.registers_25\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15130_ _11126_ VGND VGND VPWR VPWR _11127_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24328_ _08340_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone75 net303 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__buf_4
XFILLER_0_161_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28096_ clknet_leaf_69_clock net1065 VGND VGND VPWR VPWR csr.minstret\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_226_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27047_ clknet_leaf_342_clock _00076_ VGND VGND VPWR VPWR decode.regfile.registers_23\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15061_ _11057_ VGND VGND VPWR VPWR _11058_ sky130_fd_sc_hd__clkbuf_8
X_24259_ _08087_ net1795 _08300_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_226_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14012_ net780 _10258_ _10265_ _10262_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18820_ _04117_ _04118_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28998_ clknet_leaf_97_clock _02011_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_18751_ _04045_ _04049_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__nor2_4
X_27949_ clknet_leaf_205_clock _00971_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_15963_ _11942_ decode.regfile.registers_30\[17\] _11722_ _11723_ _11724_ VGND VGND
+ VPWR VPWR _11943_ sky130_fd_sc_hd__o2111a_1
X_17702_ _10929_ decode.regfile.registers_28\[22\] _02992_ VGND VGND VPWR VPWR _03107_
+ sky130_fd_sc_hd__o21a_1
X_14914_ _10912_ _10913_ _10921_ _10944_ VGND VGND VPWR VPWR _10945_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_106_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15894_ _11446_ decode.regfile.registers_26\[15\] _11447_ _11348_ _10993_ VGND VGND
+ VPWR VPWR _11876_ sky130_fd_sc_hd__o2111a_1
X_18682_ _03662_ execute.io_reg_pc\[0\] net100 _03663_ _03980_ VGND VGND VPWR VPWR
+ _03981_ sky130_fd_sc_hd__o221a_2
XFILLER_0_203_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29619_ clknet_leaf_280_clock _02632_ VGND VGND VPWR VPWR decode.regfile.registers_11\[25\]
+ sky130_fd_sc_hd__dfxtp_2
X_17633_ decode.regfile.registers_4\[21\] decode.regfile.registers_5\[21\] _12508_
+ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_177_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14845_ _10705_ _10815_ _10887_ VGND VGND VPWR VPWR _10888_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_177_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14776_ _10814_ decode.id_ex_pc_reg\[11\] VGND VGND VPWR VPWR _10819_ sky130_fd_sc_hd__nand2_1
X_17564_ decode.regfile.registers_15\[19\] _12874_ _12576_ VGND VGND VPWR VPWR _02972_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_67_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19303_ _04443_ _04589_ _04590_ _04594_ _04595_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__a32o_1
X_16515_ _12479_ _11236_ _12480_ VGND VGND VPWR VPWR _12481_ sky130_fd_sc_hd__a21o_1
X_13727_ _10073_ VGND VGND VPWR VPWR _10074_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17495_ _13441_ _13442_ VGND VGND VPWR VPWR _13443_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19234_ _04527_ _04528_ _04500_ _04464_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_184_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16446_ _11489_ decode.regfile.registers_28\[29\] decode.regfile.registers_29\[29\]
+ _11063_ _11245_ VGND VGND VPWR VPWR _12414_ sky130_fd_sc_hd__o221a_1
X_13658_ _10014_ VGND VGND VPWR VPWR _10015_ sky130_fd_sc_hd__buf_4
XFILLER_0_186_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_16__f_clock clknet_2_2_0_clock VGND VGND VPWR VPWR clknet_5_16__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_170_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19165_ _03971_ _04254_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__nor2_1
X_16377_ _11346_ decode.regfile.registers_30\[28\] _12095_ _12096_ _12097_ VGND VGND
+ VPWR VPWR _12346_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13589_ _09953_ VGND VGND VPWR VPWR _09954_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_186_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18116_ _03485_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15328_ decode.regfile.registers_18\[1\] _11269_ _11271_ _11323_ VGND VGND VPWR VPWR
+ _11324_ sky130_fd_sc_hd__a211o_1
XFILLER_0_171_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19096_ _03635_ decode.id_ex_aluop_reg\[2\] _03633_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_2_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18047_ _10939_ _03068_ decode.regfile.registers_27\[31\] _12506_ VGND VGND VPWR
+ VPWR _03443_ sky130_fd_sc_hd__or4_1
X_15259_ _11063_ VGND VGND VPWR VPWR _11255_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19998_ _05223_ _05224_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__nor2_1
X_18949_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_129_Left_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_1330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21960_ net1446 _06574_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20911_ _05935_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__clkbuf_1
X_21891_ csr._mcycle_T_2\[16\] _06521_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23630_ net1547 _10821_ _07961_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20842_ _05897_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23561_ net1984 _07918_ _07915_ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__or3b_1
X_20773_ _05855_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25300_ _08880_ net2753 VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22512_ _07066_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__buf_4
X_26280_ _09417_ VGND VGND VPWR VPWR _09471_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23492_ decode.control.io_funct7\[6\] _07876_ _07873_ VGND VGND VPWR VPWR _07885_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_107_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25231_ _08070_ net2075 _08837_ VGND VGND VPWR VPWR _08845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22443_ _06754_ fetch.btb.btbTable\[10\]\[1\] fetch.bht.bhtTable_valid\[10\] VGND
+ VGND VPWR VPWR _07038_ sky130_fd_sc_hd__and3b_1
XFILLER_0_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25162_ net419 _08809_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22374_ fetch.bht.bhtTable_tag\[12\]\[16\] fetch.bht.bhtTable_tag\[13\]\[16\] _06643_
+ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24113_ _08229_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__clkbuf_1
X_21325_ net1216 _10795_ _06168_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__mux2_1
X_25093_ _08774_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28921_ clknet_leaf_127_clock _01934_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_24044_ net1448 execute.io_target_pc\[10\] _08187_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21256_ _10795_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__buf_2
Xhold450 decode.control.io_funct7\[3\] VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 decode.regfile.registers_28\[6\] VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold472 csr._mcycle_T_3\[60\] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap191 _10127_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_221_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20207_ _05399_ _05402_ _05400_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__o21bai_1
Xhold483 decode.regfile.registers_26\[3\] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28852_ clknet_leaf_117_clock _01865_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold494 decode.regfile.registers_29\[25\] VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21187_ _06086_ _06082_ net1456 VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__and3_1
XFILLER_0_229_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_147_Left_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27803_ clknet_leaf_331_clock _00832_ VGND VGND VPWR VPWR memory.io_wb_readdata\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_20138_ decode.id_ex_imm_reg\[20\] _10867_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__xor2_2
XFILLER_0_216_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28783_ clknet_leaf_110_clock _01796_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_25995_ _08916_ _09287_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__nand2_1
X_20069_ decode.id_ex_imm_reg\[9\] _10706_ _05285_ _05279_ VGND VGND VPWR VPWR _05286_
+ sky130_fd_sc_hd__a2bb2o_1
X_27734_ clknet_leaf_65_clock _00763_ VGND VGND VPWR VPWR execute.csr_write_enable_out_reg
+ sky130_fd_sc_hd__dfxtp_1
X_24946_ net1929 _08676_ _08677_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__o21a_1
Xhold1150 decode.io_id_pc\[3\] VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1161 fetch.bht.bhtTable_tag\[4\]\[12\] VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 fetch.bht.bhtTable_tag\[9\]\[15\] VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 fetch.bht.bhtTable_target_pc\[4\]\[0\] VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__dlygate4sd3_1
X_24877_ csr.mcycle\[10\] csr.mcycle\[9\] csr.mcycle\[12\] csr.mcycle\[11\] VGND VGND
+ VPWR VPWR _08627_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_321_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_321_clock
+ sky130_fd_sc_hd__clkbuf_8
X_27665_ clknet_leaf_27_clock _00694_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1194 decode.regfile.registers_28\[28\] VGND VGND VPWR VPWR net1421 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_219_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _10672_ VGND VGND VPWR VPWR _10673_ sky130_fd_sc_hd__clkbuf_4
X_29404_ clknet_leaf_247_clock _02417_ VGND VGND VPWR VPWR decode.regfile.registers_5\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_23828_ _08072_ net2227 _08058_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_219_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26616_ _09663_ VGND VGND VPWR VPWR _09664_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_213_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27596_ clknet_leaf_147_clock _00625_ VGND VGND VPWR VPWR execute.io_target_pc\[5\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29335_ clknet_leaf_226_clock _02348_ VGND VGND VPWR VPWR decode.regfile.registers_2\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_26547_ net2526 _09622_ _09625_ _09619_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__o211a_1
X_14561_ _10603_ VGND VGND VPWR VPWR _10604_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_215_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23759_ _08031_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_172_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_156_Left_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13512_ _09891_ _09888_ VGND VGND VPWR VPWR _09892_ sky130_fd_sc_hd__nor2_4
X_16300_ _11396_ _12269_ _12270_ _12271_ VGND VGND VPWR VPWR _12272_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17280_ _12497_ _12539_ _12503_ decode.regfile.registers_7\[12\] _12645_ VGND VGND
+ VPWR VPWR _13233_ sky130_fd_sc_hd__o32a_1
XFILLER_0_95_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29266_ clknet_leaf_224_clock _02279_ VGND VGND VPWR VPWR decode.regfile.registers_0\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26478_ net2270 _09578_ _09585_ _09582_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__o211a_1
X_14492_ _10122_ _10530_ VGND VGND VPWR VPWR _10542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16231_ _11263_ decode.regfile.registers_22\[24\] _11404_ _11264_ _11265_ VGND VGND
+ VPWR VPWR _12204_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_36_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28217_ clknet_leaf_84_clock net1207 VGND VGND VPWR VPWR csr.mscratch\[19\] sky130_fd_sc_hd__dfxtp_1
X_25429_ net2263 _08951_ _08963_ _08950_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29197_ clknet_leaf_163_clock _02210_ VGND VGND VPWR VPWR fetch.btb.btbTable\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16162_ decode.regfile.registers_17\[22\] _11128_ _11106_ VGND VGND VPWR VPWR _12137_
+ sky130_fd_sc_hd__o21ai_1
X_28148_ clknet_leaf_192_clock _01170_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15113_ _11109_ VGND VGND VPWR VPWR _11110_ sky130_fd_sc_hd__clkbuf_4
X_28079_ clknet_leaf_204_clock _01101_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16093_ decode.regfile.registers_8\[20\] _11285_ _11365_ decode.regfile.registers_9\[20\]
+ _11381_ VGND VGND VPWR VPWR _12070_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15044_ decode.immGen._imm_T_24\[11\] VGND VGND VPWR VPWR _11041_ sky130_fd_sc_hd__inv_2
X_19921_ _03862_ _05164_ _03854_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_165_Left_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19852_ _05101_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18803_ decode.id_ex_rs2_data_reg\[13\] net199 _04096_ _03763_ VGND VGND VPWR VPWR
+ _04102_ sky130_fd_sc_hd__o22a_4
X_19783_ _05056_ decode.id_ex_imm_reg\[25\] _04388_ _03837_ VGND VGND VPWR VPWR _05057_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16995_ _11015_ _10937_ decode.regfile.registers_23\[5\] _12520_ VGND VGND VPWR VPWR
+ _12955_ sky130_fd_sc_hd__or4_1
XFILLER_0_218_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18734_ _03816_ _04032_ net353 VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_30_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15946_ decode.regfile.registers_13\[16\] _10639_ _11186_ _11925_ _11926_ VGND VGND
+ VPWR VPWR _11927_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_69_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18665_ _03894_ _03958_ _03963_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15877_ _11225_ _11125_ _11104_ _11859_ VGND VGND VPWR VPWR _11860_ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17616_ _13250_ decode.regfile.registers_24\[20\] _13170_ _13083_ _13367_ VGND VGND
+ VPWR VPWR _03023_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_59_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14828_ csr.io_mem_pc\[13\] VGND VGND VPWR VPWR _10871_ sky130_fd_sc_hd__clkbuf_8
X_18596_ execute.io_mem_memtoreg\[1\] execute.io_mem_memtoreg\[0\] execute.io_reg_pc\[19\]
+ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17547_ _13451_ net2794 _13492_ VGND VGND VPWR VPWR _13493_ sky130_fd_sc_hd__o21a_1
X_14759_ _10801_ decode.id_ex_pc_reg\[19\] VGND VGND VPWR VPWR _10802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17478_ decode.regfile.registers_4\[17\] _12548_ _13145_ decode.regfile.registers_5\[17\]
+ _12625_ VGND VGND VPWR VPWR _13426_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19217_ _04508_ _04512_ _04491_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_60_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16429_ decode.regfile.registers_11\[29\] _11071_ _11204_ _11407_ VGND VGND VPWR
+ VPWR _12397_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_99_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19148_ _04444_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__buf_4
XFILLER_0_229_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19079_ _04376_ _04160_ _04254_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21110_ _05949_ _06046_ net626 VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22090_ _06684_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21041_ execute.csr_read_data_out_reg\[10\] _06002_ _05998_ VGND VGND VPWR VPWR _06006_
+ sky130_fd_sc_hd__and3_1
Xfanout226 net70 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24800_ _08093_ net1329 _08585_ VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25780_ _09155_ VGND VGND VPWR VPWR _09170_ sky130_fd_sc_hd__clkbuf_4
X_22992_ _07069_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24731_ _08093_ net1236 _08542_ VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21943_ csr.io_csr_write_address\[1\] _06457_ _06315_ _06470_ VGND VGND VPWR VPWR
+ _06570_ sky130_fd_sc_hd__or4b_1
XFILLER_0_96_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27450_ clknet_leaf_149_clock _00479_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_24662_ _08514_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21874_ _06518_ _06519_ _06520_ _06522_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26401_ _09381_ _09535_ VGND VGND VPWR VPWR _09541_ sky130_fd_sc_hd__nand2_1
X_23613_ _06143_ net1698 _07952_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20825_ _05888_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__clkbuf_1
X_27381_ clknet_leaf_10_clock _00410_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[22\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_210_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24593_ net1181 execute.io_target_pc\[18\] _08473_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29120_ clknet_leaf_68_clock _02133_ VGND VGND VPWR VPWR csr.mcycle\[4\] sky130_fd_sc_hd__dfxtp_2
X_26332_ _09387_ _09492_ VGND VGND VPWR VPWR _09501_ sky130_fd_sc_hd__nand2_1
X_23544_ decode.id_ex_memread_reg VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_212_1282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20756_ _05439_ _05201_ csr.io_csr_address\[5\] VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__and3b_1
XFILLER_0_37_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29051_ clknet_leaf_172_clock _02064_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_210_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26263_ net598 _09447_ _09461_ _09458_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_210_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23475_ _03546_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20687_ _05809_ decode.id_ex_rs1_data_reg\[5\] _05798_ VGND VGND VPWR VPWR _05810_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_210_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25214_ _08053_ net2112 _08041_ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__mux2_1
X_28002_ clknet_leaf_205_clock _01024_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_22426_ _06622_ _07020_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26194_ net201 VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25145_ net93 _06248_ _10916_ _07415_ _05856_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__o311a_2
X_22357_ fetch.bht.bhtTable_tag\[8\]\[14\] fetch.bht.bhtTable_tag\[9\]\[14\] fetch.bht.bhtTable_tag\[10\]\[14\]
+ fetch.bht.bhtTable_tag\[11\]\[14\] net302 _06620_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21308_ net1625 csr.io_mem_pc\[12\] _06157_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25076_ csr.mcycle\[28\] csr.mcycle\[27\] _08759_ csr.mcycle\[29\] VGND VGND VPWR
+ VPWR _08765_ sky130_fd_sc_hd__a31oi_1
X_22288_ _06673_ _06882_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__nor2_1
X_28904_ clknet_leaf_100_clock _01917_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24027_ net965 execute.io_target_pc\[2\] _08014_ VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_208_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21239_ _06118_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__clkbuf_1
Xhold280 decode.regfile.registers_1\[24\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_208_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29884_ clknet_leaf_305_clock _02897_ VGND VGND VPWR VPWR decode.regfile.registers_20\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold291 decode.regfile.registers_31\[27\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__buf_1
X_28835_ clknet_leaf_130_clock _01848_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15800_ _11225_ _11125_ _11216_ decode.regfile.registers_17\[12\] _11128_ VGND VGND
+ VPWR VPWR _11785_ sky130_fd_sc_hd__o32a_1
XFILLER_0_176_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28766_ clknet_leaf_176_clock _01779_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_16780_ _12497_ _12503_ _12637_ decode.regfile.registers_11\[1\] VGND VGND VPWR VPWR
+ _12744_ sky130_fd_sc_hd__or4b_1
X_13992_ _10008_ _10244_ VGND VGND VPWR VPWR _10254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25978_ _08975_ _09241_ VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_260_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_260_clock
+ sky130_fd_sc_hd__clkbuf_8
X_15731_ _11250_ decode.regfile.registers_25\[10\] _11090_ _11486_ _11717_ VGND VGND
+ VPWR VPWR _11718_ sky130_fd_sc_hd__o311a_1
X_27717_ clknet_leaf_20_clock _00746_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_24929_ net468 _08665_ _08666_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__o21a_1
X_28697_ clknet_leaf_122_clock _01710_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18450_ execute.io_mem_rd\[2\] csr.io_csr_address\[2\] VGND VGND VPWR VPWR _03749_
+ sky130_fd_sc_hd__or2b_1
XANTENNA_120 _10556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27648_ clknet_leaf_48_clock net170 VGND VGND VPWR VPWR execute.io_reg_pc\[25\] sky130_fd_sc_hd__dfxtp_1
X_15662_ decode.regfile.registers_11\[9\] _11180_ _11509_ decode.regfile.registers_10\[9\]
+ _11186_ VGND VGND VPWR VPWR _11650_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_131 _10662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17401_ decode.regfile.registers_8\[15\] _12892_ _12602_ _13350_ VGND VGND VPWR VPWR
+ _13351_ sky130_fd_sc_hd__o211a_1
XANTENNA_142 decode.id_ex_rs1_data_reg\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_153 _10662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _10655_ decode.id_ex_ex_rd_reg\[2\] VGND VGND VPWR VPWR _10656_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_120_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18381_ decode.id_ex_ex_rs1_reg\[2\] VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__inv_2
X_15593_ decode.regfile.registers_5\[7\] _11290_ _10635_ _11135_ VGND VGND VPWR VPWR
+ _11583_ sky130_fd_sc_hd__o2bb2a_1
X_27579_ clknet_leaf_171_clock _00608_ VGND VGND VPWR VPWR csr.io_mem_pc\[20\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_275_clock clknet_5_21__leaf_clock VGND VGND VPWR VPWR clknet_leaf_275_clock
+ sky130_fd_sc_hd__clkbuf_8
X_29318_ clknet_leaf_228_clock _02331_ VGND VGND VPWR VPWR decode.regfile.registers_2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14544_ _10578_ _10579_ decode.control.io_funct3\[2\] _10582_ _10586_ VGND VGND VPWR
+ VPWR _10587_ sky130_fd_sc_hd__o221a_4
X_17332_ decode.regfile.registers_16\[13\] _12576_ _12579_ _13283_ VGND VGND VPWR
+ VPWR _13284_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29249_ clknet_leaf_233_clock _02262_ VGND VGND VPWR VPWR decode.regfile.registers_0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_17263_ _12496_ _13213_ _13214_ _13216_ VGND VGND VPWR VPWR _13217_ sky130_fd_sc_hd__a31o_1
X_14475_ net443 _10520_ _10532_ _10522_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19002_ _04300_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16214_ _12173_ _12186_ _12187_ VGND VGND VPWR VPWR _12188_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17194_ decode.regfile.registers_8\[10\] _12888_ _12606_ VGND VGND VPWR VPWR _13149_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16145_ _11225_ _11125_ _11216_ decode.regfile.registers_17\[21\] _11128_ VGND VGND
+ VPWR VPWR _12121_ sky130_fd_sc_hd__o32a_1
XFILLER_0_3_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_173_Left_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_4_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16076_ _11761_ net443 _12015_ _12053_ _11760_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_213_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_213_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_90_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15027_ _10662_ _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__a31o_1
X_19904_ _04436_ _05072_ _05172_ _04392_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19835_ _05105_ _04401_ _05106_ _04504_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_127_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1908 decode.regfile.registers_4\[29\] VGND VGND VPWR VPWR net2135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1919 csr._minstret_T_3\[49\] VGND VGND VPWR VPWR net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19766_ _04442_ _04245_ _04386_ _04806_ _04728_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__o311a_4
Xclkbuf_leaf_228_clock clknet_5_22__leaf_clock VGND VGND VPWR VPWR clknet_leaf_228_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16978_ decode.regfile.registers_3\[5\] _12628_ _12732_ VGND VGND VPWR VPWR _12938_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 net383 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
X_18717_ decode.id_ex_rs2_data_reg\[2\] _03758_ net235 VGND VGND VPWR VPWR _04016_
+ sky130_fd_sc_hd__nand3b_2
X_15929_ _11571_ net402 _11722_ _11723_ _11724_ VGND VGND VPWR VPWR _11910_ sky130_fd_sc_hd__o2111a_1
X_19697_ _04189_ _03894_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_88_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_182_Left_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18648_ _03707_ decode.id_ex_imm_reg\[21\] _03945_ _03946_ VGND VGND VPWR VPWR _03947_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_94_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_31__f_clock clknet_2_3_0_clock VGND VGND VPWR VPWR clknet_5_31__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_18579_ decode.io_wb_rd\[0\] _03721_ _03755_ _10194_ _03732_ VGND VGND VPWR VPWR
+ _03878_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20610_ csr.minstret\[23\] _05658_ _05556_ csr._minstret_T_3\[55\] _05746_ VGND VGND
+ VPWR VPWR _05747_ sky130_fd_sc_hd__o221a_1
XFILLER_0_191_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21590_ csr.io_csr_write_address\[11\] net216 _06314_ _06316_ VGND VGND VPWR VPWR
+ _06319_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20541_ _05540_ csr.io_mret_vector\[14\] _05565_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23260_ _07122_ _07691_ VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__nor2_1
X_20472_ _05541_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_191_Left_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22211_ _06642_ _06801_ _06805_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23191_ net74 net73 _07582_ _06887_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22142_ _06734_ _06677_ _00002_ _06736_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_113_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22073_ _06667_ _06624_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__or2b_1
X_26950_ _10047_ _09849_ VGND VGND VPWR VPWR _09857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25901_ net2174 _09200_ _09238_ _09235_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__o211a_1
X_21024_ _05996_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26881_ _09408_ _09806_ VGND VGND VPWR VPWR _09817_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_203_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28620_ clknet_leaf_87_clock _01633_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_203_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25832_ _09198_ VGND VGND VPWR VPWR _09200_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28551_ clknet_leaf_182_clock _01564_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_22975_ _07422_ _07371_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__and2_1
X_25763_ net1870 _09156_ _09160_ _09153_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_195_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27502_ clknet_leaf_29_clock _00531_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dfxtp_1
X_24714_ _08076_ net1225 _08531_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_195_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21926_ _06557_ _06543_ _06544_ _06558_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__o211a_1
X_28482_ clknet_leaf_206_clock _01495_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_25694_ _08918_ _09112_ VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24645_ _08505_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27433_ clknet_leaf_41_clock _00462_ VGND VGND VPWR VPWR decode.id_ex_immsrc_reg
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_171_1082 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21857_ net777 _06497_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20808_ _05866_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__buf_2
X_24576_ net1118 execute.io_target_pc\[10\] _08462_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27364_ clknet_leaf_31_clock _00393_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_21788_ csr.io_csr_write_address\[10\] csr.io_csr_write_address\[11\] csr.io_csr_write_address\[9\]
+ csr.io_csr_write_address\[8\] VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_93_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29103_ clknet_leaf_17_clock _02116_ VGND VGND VPWR VPWR csr._mcycle_T_3\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23527_ net1955 _07904_ _07901_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__or3b_1
XFILLER_0_19_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26315_ _09490_ VGND VGND VPWR VPWR _09491_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27295_ clknet_leaf_1_clock _00324_ VGND VGND VPWR VPWR decode.regfile.registers_31\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20739_ _05831_ _05813_ decode.id_ex_rs1_data_reg\[26\] _05840_ _00713_ VGND VGND
+ VPWR VPWR _00745_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_154_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29034_ clknet_leaf_98_clock _02047_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14260_ net774 _10403_ _10408_ _10398_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__o211a_1
X_26246_ _09377_ _09448_ VGND VGND VPWR VPWR _09452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23458_ _11011_ _07862_ _07859_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__or3b_1
XFILLER_0_190_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22409_ _07001_ _07003_ _06790_ _06640_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_150_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14191_ _10128_ _10331_ VGND VGND VPWR VPWR _10368_ sky130_fd_sc_hd__nand2_1
X_26177_ net2511 _09395_ _09403_ _09394_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23389_ net88 _06795_ _07783_ VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25128_ _08792_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25059_ csr._mcycle_T_2\[24\] _08710_ _08751_ csr.mcycle\[24\] VGND VGND VPWR VPWR
+ _08753_ sky130_fd_sc_hd__a211oi_1
X_29936_ clknet_leaf_341_clock _02949_ VGND VGND VPWR VPWR decode.regfile.registers_21\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_17950_ _12649_ _12615_ _12880_ decode.regfile.registers_6\[29\] _03347_ VGND VGND
+ VPWR VPWR _03348_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_130_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16901_ _10927_ decode.regfile.registers_24\[3\] _10933_ _12759_ _12862_ VGND VGND
+ VPWR VPWR _12863_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_218_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17881_ decode.regfile.registers_12\[27\] _12489_ _12498_ _12540_ VGND VGND VPWR
+ VPWR _03281_ sky130_fd_sc_hd__or4_1
X_29867_ clknet_leaf_300_clock _02880_ VGND VGND VPWR VPWR decode.regfile.registers_19\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19620_ _04225_ _04242_ _04425_ _04899_ _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__a221o_1
X_28818_ clknet_leaf_106_clock _01831_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_16832_ decode.regfile.registers_11\[2\] _12595_ _12789_ _12793_ _12794_ VGND VGND
+ VPWR VPWR _12795_ sky130_fd_sc_hd__a221o_1
XFILLER_0_228_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29798_ clknet_leaf_296_clock _02811_ VGND VGND VPWR VPWR decode.regfile.registers_17\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19551_ _04186_ _04095_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__nor2_1
X_28749_ clknet_leaf_99_clock _01762_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16763_ decode.regfile.registers_4\[1\] _12617_ _12619_ decode.regfile.registers_5\[1\]
+ VGND VGND VPWR VPWR _12727_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13975_ _10242_ VGND VGND VPWR VPWR _10244_ sky130_fd_sc_hd__buf_2
X_18502_ _03795_ _03800_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__or2_1
XFILLER_0_214_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15714_ _11136_ _11699_ _11700_ VGND VGND VPWR VPWR _11701_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19482_ _04112_ net285 _04274_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__mux2_1
X_16694_ _12658_ VGND VGND VPWR VPWR _12659_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_213_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18433_ csr.io_csr_address\[4\] decode.io_wb_rd\[4\] VGND VGND VPWR VPWR _03732_
+ sky130_fd_sc_hd__or2b_1
X_15645_ decode.regfile.registers_18\[8\] _11455_ _11456_ VGND VGND VPWR VPWR _11634_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18364_ _03657_ _03662_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__nand2_1
X_15576_ _11250_ decode.regfile.registers_27\[6\] _11258_ VGND VGND VPWR VPWR _11567_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17315_ decode.regfile.registers_7\[13\] _12611_ _12623_ decode.regfile.registers_6\[13\]
+ _12888_ VGND VGND VPWR VPWR _13267_ sky130_fd_sc_hd__a221oi_1
X_14527_ _10566_ _10565_ _10564_ VGND VGND VPWR VPWR _10571_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18295_ _03612_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17246_ _12499_ _12504_ _12650_ _13199_ VGND VGND VPWR VPWR _13200_ sky130_fd_sc_hd__o31a_1
XFILLER_0_189_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14458_ net457 _10520_ _10523_ _10522_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17177_ _12695_ _13130_ _13131_ _13132_ VGND VGND VPWR VPWR _13133_ sky130_fd_sc_hd__a31o_1
X_14389_ net439 _10477_ _10483_ _10481_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_152_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_152_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16128_ _11190_ _11148_ _11154_ decode.regfile.registers_0\[21\] VGND VGND VPWR VPWR
+ _12104_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_110_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16059_ _12018_ _12036_ VGND VGND VPWR VPWR _12037_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2406 csr._csr_read_data_T_8\[13\] VGND VGND VPWR VPWR net2633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2417 _02141_ VGND VGND VPWR VPWR net2644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_167_clock clknet_5_25__leaf_clock VGND VGND VPWR VPWR clknet_leaf_167_clock
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2428 decode.regfile.registers_9\[28\] VGND VGND VPWR VPWR net2655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2439 decode.regfile.registers_0\[24\] VGND VGND VPWR VPWR net2666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1705 decode.regfile.registers_22\[26\] VGND VGND VPWR VPWR net1932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1716 fetch.bht.bhtTable_target_pc\[5\]\[18\] VGND VGND VPWR VPWR net1943 sky130_fd_sc_hd__dlygate4sd3_1
X_19818_ _03819_ _03817_ _03775_ _03820_ _03825_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_208_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1727 decode.regfile.registers_19\[9\] VGND VGND VPWR VPWR net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1738 decode.regfile.registers_11\[29\] VGND VGND VPWR VPWR net1965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1749 decode.regfile.registers_2\[6\] VGND VGND VPWR VPWR net1976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19749_ _05022_ _05023_ _04190_ _04195_ _04193_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_194_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22760_ _06134_ net1705 _07265_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21711_ csr.minstret\[23\] csr.minstret\[24\] _06411_ VGND VGND VPWR VPWR _06412_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22691_ csr._mcycle_T_2\[21\] _07223_ VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24430_ _08057_ net1660 _08389_ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21642_ csr.minstret\[12\] _06338_ _06355_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_105_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_105_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24361_ _08357_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21573_ _06307_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 _05621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 _08956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26100_ _08945_ _09353_ VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__nand2_1
X_23312_ net222 net223 _07716_ net221 VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__a31o_1
XANTENNA_42 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20524_ _05540_ _03741_ _05528_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__or3b_2
XFILLER_0_105_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27080_ clknet_leaf_346_clock _00109_ VGND VGND VPWR VPWR decode.regfile.registers_24\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_53 _10598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24292_ _08321_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_64 _11011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _11092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_86 _13475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26031_ net2488 _09313_ _09314_ _09305_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__o211a_1
X_23243_ net224 net76 _06887_ _07613_ net79 VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__a41o_1
XFILLER_0_160_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_97 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20455_ _05554_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23174_ _07085_ _07604_ _07610_ net280 VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__a211o_1
XFILLER_0_162_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20386_ _05533_ _05547_ _05548_ _05414_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__o31a_1
X_22125_ _06671_ _06719_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27982_ clknet_leaf_166_clock _01004_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput160 net160 VGND VGND VPWR VPWR io_memory_write_data[31] sky130_fd_sc_hd__clkbuf_4
X_29721_ clknet_leaf_311_clock _02734_ VGND VGND VPWR VPWR decode.regfile.registers_14\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22056_ _06650_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__buf_4
X_26933_ _09998_ _09840_ VGND VGND VPWR VPWR _09847_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_201_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_197_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21007_ _05987_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_197_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29652_ clknet_leaf_279_clock _02665_ VGND VGND VPWR VPWR decode.regfile.registers_12\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_197_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26864_ net651 _09795_ _09807_ _09799_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__o211a_1
X_28603_ clknet_leaf_170_clock _01616_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25815_ net2582 _09183_ _09189_ _09182_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__o211a_1
X_29583_ clknet_leaf_274_clock _02596_ VGND VGND VPWR VPWR decode.regfile.registers_10\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26795_ _09398_ _09763_ VGND VGND VPWR VPWR _09768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28534_ clknet_leaf_216_clock _01547_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13760_ _10101_ VGND VGND VPWR VPWR _10102_ sky130_fd_sc_hd__buf_6
X_22958_ _07119_ VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__buf_4
XFILLER_0_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25746_ net2359 _09139_ _09149_ _09142_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21909_ csr.io_mret_vector\[21\] csr.io_mem_pc\[21\] _06539_ VGND VGND VPWR VPWR
+ _06547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28465_ clknet_leaf_138_clock _01478_ VGND VGND VPWR VPWR decode.io_id_pc\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13691_ net589 _10027_ _10043_ _10020_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22889_ _07341_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_156_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25677_ _10373_ _10240_ _08903_ _09935_ VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_156_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15430_ decode.regfile.registers_14\[3\] _11208_ _11422_ _11199_ _11423_ VGND VGND
+ VPWR VPWR _11424_ sky130_fd_sc_hd__a221o_1
X_27416_ clknet_leaf_15_clock _00445_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[25\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_214_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24628_ _08496_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__clkbuf_1
X_28396_ clknet_leaf_142_clock _01409_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_14_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15361_ _11355_ VGND VGND VPWR VPWR _11356_ sky130_fd_sc_hd__clkbuf_4
X_24559_ net915 execute.io_target_pc\[2\] _07335_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__mux2_1
X_27347_ clknet_leaf_45_clock _00376_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[20\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17100_ decode.regfile.registers_7\[8\] _12610_ _12737_ decode.regfile.registers_6\[8\]
+ _12843_ VGND VGND VPWR VPWR _13057_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14312_ _10053_ _10431_ VGND VGND VPWR VPWR _10439_ sky130_fd_sc_hd__nand2_1
X_18080_ _10910_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_124_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15292_ _11091_ _11057_ _10628_ VGND VGND VPWR VPWR _11288_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27278_ clknet_leaf_11_clock _00307_ VGND VGND VPWR VPWR decode.regfile.registers_30\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29017_ clknet_leaf_127_clock _02030_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14243_ _10069_ _10387_ VGND VGND VPWR VPWR _10399_ sky130_fd_sc_hd__nand2_1
X_17031_ decode.regfile.registers_18\[6\] _12572_ _12561_ _12989_ VGND VGND VPWR VPWR
+ _12990_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_115_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26229_ _09417_ VGND VGND VPWR VPWR _09440_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14174_ _10331_ VGND VGND VPWR VPWR _10359_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_186_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_84_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18982_ _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _02990_ _03068_ decode.regfile.registers_27\[28\] _12506_ VGND VGND VPWR
+ VPWR _03332_ sky130_fd_sc_hd__or4_1
X_29919_ clknet_leaf_335_clock _02932_ VGND VGND VPWR VPWR decode.regfile.registers_21\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17864_ decode.regfile.registers_18\[27\] _12571_ _12560_ VGND VGND VPWR VPWR _03264_
+ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_99_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_99_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19603_ _04872_ _04874_ _04882_ _04884_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__o31a_1
XFILLER_0_205_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16815_ _12630_ VGND VGND VPWR VPWR _12778_ sky130_fd_sc_hd__buf_4
X_17795_ _12612_ _03195_ _03196_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_85_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19534_ _04186_ _04782_ _04795_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_141_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16746_ _10931_ net665 _12487_ VGND VGND VPWR VPWR _12710_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_141_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13958_ net2318 _10226_ _10233_ _10232_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19465_ _04408_ _03705_ _04305_ _04751_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_22_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_124_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16677_ _10610_ _12626_ _12629_ decode.regfile.registers_3\[0\] _12641_ VGND VGND
+ VPWR VPWR _12642_ sky130_fd_sc_hd__o221a_1
X_13889_ _10142_ _10152_ VGND VGND VPWR VPWR _10192_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_210 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_221 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_232 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18416_ net208 VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__clkbuf_4
X_15628_ decode.regfile.registers_2\[8\] _11369_ _11615_ _11616_ VGND VGND VPWR VPWR
+ _11617_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_124_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_243 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_254 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19396_ _04683_ _04663_ _04167_ _04165_ _04401_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__a41o_1
XFILLER_0_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_265 _06250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_276 _11012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_287 _12504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18347_ decode.id_ex_ex_rs1_reg\[2\] execute.io_mem_rd\[2\] VGND VGND VPWR VPWR _03646_
+ sky130_fd_sc_hd__or2b_1
XINSDIODE1_298 csr._minstret_T_3\[51\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15559_ decode.regfile.registers_10\[6\] _10637_ _11131_ _11315_ VGND VGND VPWR VPWR
+ _11550_ sky130_fd_sc_hd__o31a_1
XFILLER_0_86_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_37_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18278_ _03603_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_204_Right_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17229_ _12694_ VGND VGND VPWR VPWR _13183_ sky130_fd_sc_hd__buf_2
Xinput40 io_memory_read_data[15] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
XFILLER_0_71_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 io_memory_read_data[25] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_1
Xhold802 fetch.bht.bhtTable_target_pc\[3\]\[28\] VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput62 io_memory_read_data[6] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_163_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold813 fetch.bht.bhtTable_target_pc\[12\]\[5\] VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__dlygate4sd3_1
X_20240_ _10834_ _10747_ decode.id_ex_pc_reg\[4\] _10704_ VGND VGND VPWR VPWR _05430_
+ sky130_fd_sc_hd__and4_1
Xhold824 fetch.bht.bhtTable_target_pc\[3\]\[11\] VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 fetch.bht.bhtTable_tag\[4\]\[24\] VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 fetch.bht.bhtTable_target_pc\[15\]\[20\] VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 fetch.bht.bhtTable_target_pc\[11\]\[9\] VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold868 fetch.bht.bhtTable_target_pc\[5\]\[15\] VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__dlygate4sd3_1
X_20171_ _00572_ _05226_ _05373_ _05239_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold879 fetch.bht.bhtTable_target_pc\[12\]\[18\] VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2203 decode.regfile.registers_7\[6\] VGND VGND VPWR VPWR net2430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2214 decode.regfile.registers_11\[0\] VGND VGND VPWR VPWR net2441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2225 decode.regfile.registers_5\[27\] VGND VGND VPWR VPWR net2452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2236 decode.regfile.registers_21\[25\] VGND VGND VPWR VPWR net2463 sky130_fd_sc_hd__dlygate4sd3_1
X_23930_ _08135_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2247 decode.regfile.registers_23\[2\] VGND VGND VPWR VPWR net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1502 decode.regfile.registers_16\[0\] VGND VGND VPWR VPWR net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 fetch.bht.bhtTable_target_pc\[5\]\[7\] VGND VGND VPWR VPWR net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2258 decode.regfile.registers_24\[27\] VGND VGND VPWR VPWR net2485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2269 decode.regfile.registers_28\[18\] VGND VGND VPWR VPWR net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 decode.regfile.registers_22\[1\] VGND VGND VPWR VPWR net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 fetch.bht.bhtTable_tag\[9\]\[19\] VGND VGND VPWR VPWR net1762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23861_ execute.io_target_pc\[22\] VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__buf_2
Xhold1546 decode.regfile.registers_5\[13\] VGND VGND VPWR VPWR net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 fetch.bht.bhtTable_tag\[11\]\[19\] VGND VGND VPWR VPWR net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1568 fetch.bht.bhtTable_target_pc\[6\]\[18\] VGND VGND VPWR VPWR net1795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1579 fetch.bht.bhtTable_target_pc\[11\]\[3\] VGND VGND VPWR VPWR net1806 sky130_fd_sc_hd__dlygate4sd3_1
X_22812_ _07301_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__clkbuf_1
X_25600_ _08975_ _09023_ VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_192_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23792_ _08048_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26580_ net1968 _09636_ _09643_ _09635_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22743_ _06117_ net1192 _09903_ VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__mux2_1
X_25531_ _09025_ _09026_ VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28250_ clknet_leaf_78_clock _01272_ VGND VGND VPWR VPWR csr._minstret_T_3\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_25462_ _08914_ _08980_ VGND VGND VPWR VPWR _08986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22674_ net2096 _07222_ _07224_ _07221_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__o211a_1
X_24413_ net833 execute.io_target_pc\[29\] _09911_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__mux2_1
X_27201_ clknet_leaf_364_clock _00230_ VGND VGND VPWR VPWR decode.regfile.registers_28\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_21625_ _06317_ _06342_ csr.minstret\[6\] csr.minstret\[7\] VGND VGND VPWR VPWR _06346_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_118_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28181_ clknet_leaf_59_clock _01203_ VGND VGND VPWR VPWR csr.io_mret_vector\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_25393_ net2048 _08928_ _08938_ _08927_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24344_ _08348_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27132_ clknet_leaf_357_clock _00161_ VGND VGND VPWR VPWR decode.regfile.registers_26\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_21556_ _06298_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27063_ clknet_leaf_350_clock _00092_ VGND VGND VPWR VPWR decode.regfile.registers_24\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20507_ _05657_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__clkbuf_1
X_24275_ _08103_ net1309 _06218_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21487_ _06260_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26014_ _09263_ VGND VGND VPWR VPWR _09305_ sky130_fd_sc_hd__buf_2
X_23226_ fetch.bht.bhtTable_target_pc\[10\]\[19\] fetch.bht.bhtTable_target_pc\[11\]\[19\]
+ _07067_ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20438_ csr.minstret\[2\] _05573_ _05563_ csr._csr_read_data_T_9\[2\] VGND VGND VPWR
+ VPWR _05596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23157_ fetch.bht.bhtTable_target_pc\[8\]\[15\] fetch.bht.bhtTable_target_pc\[9\]\[15\]
+ fetch.bht.bhtTable_target_pc\[10\]\[15\] fetch.bht.bhtTable_target_pc\[11\]\[15\]
+ _07555_ _07114_ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20369_ decode.csr_write_reg _05531_ net474 VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__a21oi_1
X_22108_ _06678_ _06702_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_224_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_224_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27965_ clknet_leaf_214_clock _00987_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_23088_ net69 net68 net98 _07472_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_8_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29704_ clknet_leaf_283_clock _02717_ VGND VGND VPWR VPWR decode.regfile.registers_14\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22039_ fetch.bht.bhtTable_tag\[12\]\[22\] fetch.bht.bhtTable_tag\[13\]\[22\] fetch.bht.bhtTable_tag\[14\]\[22\]
+ fetch.bht.bhtTable_tag\[15\]\[22\] _06619_ _06624_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__mux4_1
X_14930_ _10958_ VGND VGND VPWR VPWR _10959_ sky130_fd_sc_hd__buf_2
X_26916_ net1014 _09796_ _09835_ _09836_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27896_ clknet_leaf_18_clock _00925_ VGND VGND VPWR VPWR csr._mcycle_T_2\[17\] sky130_fd_sc_hd__dfxtp_2
X_29635_ clknet_leaf_287_clock _02648_ VGND VGND VPWR VPWR decode.regfile.registers_12\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_14861_ decode.id_ex_pc_reg\[24\] _10861_ _10863_ _10864_ _10903_ VGND VGND VPWR
+ VPWR _10904_ sky130_fd_sc_hd__a221oi_1
X_26847_ _09450_ _09796_ VGND VGND VPWR VPWR _09798_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16600_ _12564_ VGND VGND VPWR VPWR _12565_ sky130_fd_sc_hd__clkbuf_4
X_13812_ memory.csr_read_data_out_reg\[31\] _09988_ _10144_ _10145_ VGND VGND VPWR
+ VPWR _10146_ sky130_fd_sc_hd__o22ai_4
X_17580_ _02986_ decode.regfile.registers_26\[19\] _13254_ _13484_ _02987_ VGND VGND
+ VPWR VPWR _02988_ sky130_fd_sc_hd__o2111a_1
X_29566_ clknet_leaf_252_clock _02579_ VGND VGND VPWR VPWR decode.regfile.registers_10\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14792_ _09891_ _10834_ VGND VGND VPWR VPWR _10835_ sky130_fd_sc_hd__nand2_1
X_26778_ net615 _09752_ _09757_ _09758_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28517_ clknet_leaf_200_clock _01530_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_16531_ _12495_ VGND VGND VPWR VPWR _12496_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13743_ _10087_ _10075_ VGND VGND VPWR VPWR _10088_ sky130_fd_sc_hd__nand2_1
X_25729_ net2356 _09139_ _09140_ _09129_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__o211a_1
X_29497_ clknet_leaf_249_clock _02510_ VGND VGND VPWR VPWR decode.regfile.registers_7\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19250_ _04439_ _04540_ _04544_ _04346_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__a2bb2o_2
X_28448_ clknet_leaf_145_clock _01461_ VGND VGND VPWR VPWR decode.io_id_pc\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16462_ decode.regfile.registers_8\[30\] _11284_ _11287_ decode.regfile.registers_9\[30\]
+ _11131_ VGND VGND VPWR VPWR _12429_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13674_ _10012_ memory.io_wb_aluresult\[10\] _09981_ memory.io_wb_readdata\[10\]
+ _09977_ VGND VGND VPWR VPWR _10029_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_175_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18201_ decode.control.io_funct7\[0\] net214 _03538_ decode.control.io_funct7\[2\]
+ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_117_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15413_ _11278_ VGND VGND VPWR VPWR _11407_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19181_ _04295_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_117_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28379_ clknet_leaf_186_clock _01392_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16393_ _11364_ decode.regfile.registers_11\[28\] _12349_ _12361_ _11690_ VGND VGND
+ VPWR VPWR _12362_ sky130_fd_sc_hd__o221a_1
XFILLER_0_66_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18132_ _03494_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15344_ _11260_ _11331_ _11337_ _11339_ VGND VGND VPWR VPWR _11340_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18063_ _03452_ _10916_ _03453_ _10018_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__and4b_1
XFILLER_0_123_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15275_ _11270_ VGND VGND VPWR VPWR _11271_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_78_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17014_ _12969_ _12971_ _12972_ VGND VGND VPWR VPWR _12973_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14226_ net629 _10376_ _10389_ _10385_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1087 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14157_ net630 _10346_ _10349_ _10344_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14088_ net756 _10302_ _10309_ _10304_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__o211a_1
X_18965_ _03709_ _04261_ _04263_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_37_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ decode.regfile.registers_8\[28\] _12592_ _10593_ _12549_ VGND VGND VPWR VPWR
+ _03315_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_143_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18896_ _04194_ _03882_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_143_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17847_ decode.regfile.registers_17\[26\] _12580_ _03228_ _03247_ _12566_ VGND VGND
+ VPWR VPWR _03248_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_33_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17778_ _02990_ _03068_ decode.regfile.registers_27\[24\] _13487_ VGND VGND VPWR
+ VPWR _03181_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19517_ _04291_ _04598_ _04345_ _04801_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16729_ _11012_ _10926_ _12500_ _10606_ VGND VGND VPWR VPWR _12694_ sky130_fd_sc_hd__or4_4
XFILLER_0_159_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19448_ _04648_ _04734_ _04541_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19379_ _04446_ _04661_ _04666_ _04668_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__o31a_1
X_21410_ _06101_ net2046 _06219_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22390_ fetch.bht.bhtTable_tag\[14\]\[9\] fetch.bht.bhtTable_tag\[15\]\[9\] _06707_
+ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21341_ _06181_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24060_ net857 VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21272_ _09910_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold610 decode.regfile.registers_26\[9\] VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 fetch.bht.bhtTable_tag\[11\]\[13\] VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23011_ _07439_ fetch.bht.bhtTable_target_pc\[15\]\[7\] _07125_ VGND VGND VPWR VPWR
+ _07457_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_25_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold632 decode.regfile.registers_18\[18\] VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__dlygate4sd3_1
X_20223_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__clkbuf_4
Xhold643 decode.regfile.registers_16\[6\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 csr._mcycle_T_2\[13\] VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold665 decode.regfile.registers_20\[30\] VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold676 fetch.bht.bhtTable_tag\[4\]\[6\] VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold687 fetch.bht.bhtTable_target_pc\[9\]\[9\] VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 fetch.bht.bhtTable_target_pc\[2\]\[28\] VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd3_1
X_20154_ decode.id_ex_imm_reg\[19\] _05340_ _05345_ _05347_ VGND VGND VPWR VPWR _05359_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_111_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2000 fetch.bht.bhtTable_target_pc\[15\]\[11\] VGND VGND VPWR VPWR net2227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2011 fetch.bht.bhtTable_target_pc\[9\]\[8\] VGND VGND VPWR VPWR net2238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2022 fetch.bht.bhtTable_target_pc\[5\]\[30\] VGND VGND VPWR VPWR net2249 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2033 decode.regfile.registers_4\[24\] VGND VGND VPWR VPWR net2260 sky130_fd_sc_hd__dlygate4sd3_1
X_27750_ clknet_leaf_325_clock _00779_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20085_ _05297_ _05299_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__xor2_1
Xhold2044 execute.csr_write_address_out_reg\[10\] VGND VGND VPWR VPWR net2271 sky130_fd_sc_hd__dlygate4sd3_1
X_24962_ csr._mcycle_T_3\[56\] csr._mcycle_T_3\[55\] _08685_ _07148_ VGND VGND VPWR
+ VPWR _08688_ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1310 fetch.bht.bhtTable_target_pc\[15\]\[24\] VGND VGND VPWR VPWR net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2055 decode.regfile.registers_18\[21\] VGND VGND VPWR VPWR net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2066 decode.regfile.registers_2\[27\] VGND VGND VPWR VPWR net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1321 decode.regfile.registers_20\[13\] VGND VGND VPWR VPWR net1548 sky130_fd_sc_hd__dlygate4sd3_1
X_26701_ _09379_ _09710_ VGND VGND VPWR VPWR _09714_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1332 fetch.bht.bhtTable_tag\[3\]\[10\] VGND VGND VPWR VPWR net1559 sky130_fd_sc_hd__dlygate4sd3_1
X_23913_ _08126_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__clkbuf_1
Xhold2077 csr._mcycle_T_3\[44\] VGND VGND VPWR VPWR net2304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2088 fetch.bht.bhtTable_tag\[13\]\[19\] VGND VGND VPWR VPWR net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 _01224_ VGND VGND VPWR VPWR net1570 sky130_fd_sc_hd__dlygate4sd3_1
X_27681_ clknet_leaf_28_clock _00710_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_24893_ csr.mcycle\[10\] csr.mcycle\[9\] csr.mcycle\[12\] csr.mcycle\[13\] VGND VGND
+ VPWR VPWR _08642_ sky130_fd_sc_hd__and4_1
Xhold1354 decode.regfile.registers_24\[11\] VGND VGND VPWR VPWR net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2099 decode.regfile.registers_14\[19\] VGND VGND VPWR VPWR net2326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1365 fetch.bht.bhtTable_target_pc\[5\]\[16\] VGND VGND VPWR VPWR net1592 sky130_fd_sc_hd__dlygate4sd3_1
X_29420_ clknet_leaf_262_clock _02433_ VGND VGND VPWR VPWR decode.regfile.registers_5\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1376 fetch.bht.bhtTable_tag\[14\]\[10\] VGND VGND VPWR VPWR net1603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26632_ net1102 _09665_ _09673_ _09660_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__o211a_1
X_23844_ _08083_ net1044 _08079_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__mux2_1
Xhold1387 fetch.bht.bhtTable_target_pc\[0\]\[25\] VGND VGND VPWR VPWR net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1398 fetch.bht.bhtTable_tag\[1\]\[6\] VGND VGND VPWR VPWR net1625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29351_ clknet_leaf_228_clock _02364_ VGND VGND VPWR VPWR decode.regfile.registers_3\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_23775_ _08039_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26563_ _09392_ _09632_ VGND VGND VPWR VPWR _09634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20987_ _05976_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__clkbuf_1
X_28302_ clknet_leaf_164_clock _00004_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25514_ decode.regfile.registers_2\[26\] _09008_ _09015_ _09004_ VGND VGND VPWR VPWR
+ _02345_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29282_ clknet_leaf_242_clock _02295_ VGND VGND VPWR VPWR decode.regfile.registers_1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_22726_ _07255_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__buf_1
X_26494_ _09566_ VGND VGND VPWR VPWR _09595_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28233_ clknet_leaf_73_clock _01255_ VGND VGND VPWR VPWR csr._minstret_T_3\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22657_ net2746 _07208_ _07214_ _07164_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25445_ net2492 _08907_ _08974_ _08972_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_188_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21608_ csr._mcycle_T_2\[3\] _06325_ _06328_ csr.minstret\[2\] net2704 VGND VGND
+ VPWR VPWR _06334_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_36_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28164_ clknet_leaf_69_clock net736 VGND VGND VPWR VPWR csr._csr_read_data_T_9\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_213_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22588_ csr._minstret_T_3\[44\] csr._minstret_T_3\[43\] _07166_ _06422_ VGND VGND
+ VPWR VPWR _07169_ sky130_fd_sc_hd__a31o_1
X_25376_ _06578_ VGND VGND VPWR VPWR _08927_ sky130_fd_sc_hd__buf_2
XFILLER_0_192_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27115_ clknet_leaf_347_clock _00144_ VGND VGND VPWR VPWR decode.regfile.registers_25\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24327_ _08089_ net1484 _08334_ VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__mux2_1
X_21539_ _06289_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone76 _00000_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_6
X_28095_ clknet_leaf_70_clock net579 VGND VGND VPWR VPWR csr.minstret\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_181_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone87 _03977_ _03979_ _03982_ _03773_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__a31o_1
X_15060_ _11056_ VGND VGND VPWR VPWR _11057_ sky130_fd_sc_hd__buf_4
X_24258_ _08304_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__clkbuf_1
X_27046_ clknet_leaf_346_clock _00075_ VGND VGND VPWR VPWR decode.regfile.registers_23\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_226_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14011_ _10058_ _10255_ VGND VGND VPWR VPWR _10265_ sky130_fd_sc_hd__nand2_1
X_23209_ _07643_ _07110_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24189_ _08083_ net1592 _08266_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28997_ clknet_leaf_134_clock _02010_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18750_ _03890_ decode.id_ex_imm_reg\[5\] _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__a21oi_4
X_27948_ clknet_leaf_205_clock _00970_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15962_ _10961_ VGND VGND VPWR VPWR _11942_ sky130_fd_sc_hd__buf_2
XFILLER_0_41_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17701_ _02990_ _03068_ decode.regfile.registers_27\[22\] _13487_ VGND VGND VPWR
+ VPWR _03106_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14913_ _10943_ VGND VGND VPWR VPWR _10944_ sky130_fd_sc_hd__buf_2
XFILLER_0_222_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18681_ execute.csr_read_data_out_reg\[0\] _03657_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__or2_1
X_27879_ clknet_leaf_25_clock _00908_ VGND VGND VPWR VPWR csr._mcycle_T_2\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _11571_ net2776 _11722_ _11723_ _11724_ VGND VGND VPWR VPWR _11875_ sky130_fd_sc_hd__o2111a_1
X_17632_ decode.regfile.registers_3\[21\] _12836_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__nand2_1
X_29618_ clknet_leaf_280_clock _02631_ VGND VGND VPWR VPWR decode.regfile.registers_11\[24\]
+ sky130_fd_sc_hd__dfxtp_2
X_14844_ csr.io_mem_pc\[4\] _09891_ _09888_ csr.io_mem_pc\[5\] VGND VGND VPWR VPWR
+ _10887_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_177_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17563_ decode.regfile.registers_14\[19\] _12670_ _13494_ _02970_ VGND VGND VPWR
+ VPWR _02971_ sky130_fd_sc_hd__o22ai_1
X_29549_ clknet_leaf_273_clock _02562_ VGND VGND VPWR VPWR decode.regfile.registers_9\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_14775_ csr.io_mem_pc\[8\] _10816_ _10817_ VGND VGND VPWR VPWR _10818_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_67_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19302_ _03637_ _04056_ _04289_ net219 VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__and4_1
X_16514_ _11436_ decode.regfile.registers_26\[31\] _11349_ _10980_ _11347_ VGND VGND
+ VPWR VPWR _12480_ sky130_fd_sc_hd__o2111a_1
X_13726_ memory.csr_read_data_out_reg\[18\] _09986_ _10071_ _10072_ VGND VGND VPWR
+ VPWR _10073_ sky130_fd_sc_hd__a2bb2o_4
X_17494_ _12712_ decode.regfile.registers_24\[17\] _12997_ _12998_ _11025_ VGND VGND
+ VPWR VPWR _13442_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_50_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19233_ _04054_ _04056_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16445_ _11251_ _11259_ decode.regfile.registers_27\[29\] _12383_ _12412_ VGND VGND
+ VPWR VPWR _12413_ sky130_fd_sc_hd__o32a_1
XFILLER_0_67_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_1284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13657_ memory.csr_read_data_out_reg\[8\] _10010_ _10011_ _10013_ VGND VGND VPWR
+ VPWR _10014_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_112_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19164_ _04321_ _04274_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16376_ _12133_ net518 _12310_ _12345_ _12132_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__o221a_1
X_13588_ net66 VGND VGND VPWR VPWR _09953_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18115_ _03482_ _03480_ _03474_ net2129 VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15327_ _11059_ _11149_ _11127_ decode.regfile.registers_17\[1\] _11322_ VGND VGND
+ VPWR VPWR _11323_ sky130_fd_sc_hd__o221a_1
X_19095_ _04373_ _04255_ _04338_ _04231_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__o211a_2
XFILLER_0_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18046_ _12968_ _03439_ _03440_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15258_ _10962_ net2479 VGND VGND VPWR VPWR _11254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14209_ _09970_ _10377_ VGND VGND VPWR VPWR _10380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15189_ _11185_ VGND VGND VPWR VPWR _11186_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19997_ net788 decode.id_ex_pc_reg\[0\] VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_35_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18948_ _04246_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18879_ _04130_ _04142_ _04177_ _04168_ _04155_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_207_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20910_ _05925_ _05933_ net40 VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__and3_1
XFILLER_0_206_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21890_ csr.io_mret_vector\[16\] _10868_ _06515_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20841_ net107 _05891_ _05887_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23560_ net2773 _07917_ _07924_ _05805_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20772_ _03452_ _10668_ _10916_ _10018_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__and4b_1
XFILLER_0_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22511_ _07102_ _07104_ _07082_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23491_ net24 _07875_ _07884_ _07879_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25230_ _08844_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__clkbuf_1
X_22442_ _07036_ net85 VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__or2b_1
XFILLER_0_174_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25161_ _08808_ _09881_ _09884_ VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__or3b_2
X_22373_ _06966_ _06967_ _06631_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24112_ net1011 execute.io_target_pc\[11\] _08221_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21324_ _06172_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25092_ _06109_ net1390 _08596_ VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28920_ clknet_leaf_120_clock _01933_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24043_ _08193_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21255_ _06129_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__clkbuf_1
Xhold440 decode.regfile.registers_3\[11\] VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold451 decode.regfile.registers_30\[15\] VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 decode.regfile.registers_12\[0\] VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__dlygate4sd3_1
X_20206_ _00577_ _05227_ _05403_ _05267_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__a2bb2oi_2
Xhold473 decode.id_ex_rs1_data_reg\[8\] VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__dlygate4sd3_1
X_28851_ clknet_leaf_139_clock _01864_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold484 decode.regfile.registers_17\[12\] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_221_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21186_ _06088_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold495 decode.regfile.registers_30\[10\] VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27802_ clknet_leaf_327_clock _00831_ VGND VGND VPWR VPWR memory.io_wb_readdata\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20137_ _00567_ _05227_ _05344_ _05267_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__a2bb2oi_2
X_28782_ clknet_leaf_109_clock _01795_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_25994_ net2294 _09286_ _09293_ _09292_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27733_ clknet_leaf_69_clock _00762_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_20068_ decode.id_ex_imm_reg\[8\] decode.id_ex_pc_reg\[8\] decode.id_ex_pc_reg\[9\]
+ decode.id_ex_imm_reg\[9\] VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__a22oi_1
X_24945_ csr._mcycle_T_3\[50\] _08676_ _06318_ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__a21oi_1
Xhold1140 decode.regfile.registers_28\[20\] VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 fetch.bht.bhtTable_target_pc\[5\]\[0\] VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 fetch.bht.bhtTable_target_pc\[14\]\[1\] VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 fetch.bht.bhtTable_tag\[0\]\[6\] VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__dlygate4sd3_1
X_27664_ clknet_leaf_28_clock _00693_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24876_ csr.mcycle\[14\] csr.mcycle\[13\] csr.mcycle\[18\] csr.mcycle\[17\] VGND
+ VGND VPWR VPWR _08626_ sky130_fd_sc_hd__and4_1
Xhold1184 fetch.bht.bhtTable_target_pc\[3\]\[13\] VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1195 fetch.bht.bhtTable_target_pc\[15\]\[0\] VGND VGND VPWR VPWR net1422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29403_ clknet_leaf_247_clock _02416_ VGND VGND VPWR VPWR decode.regfile.registers_5\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_219_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26615_ _10149_ _10240_ _03672_ VGND VGND VPWR VPWR _09663_ sky130_fd_sc_hd__and3_1
X_23827_ execute.io_target_pc\[11\] VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_219_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27595_ clknet_leaf_147_clock _00624_ VGND VGND VPWR VPWR execute.io_target_pc\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_184_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29334_ clknet_leaf_226_clock _02347_ VGND VGND VPWR VPWR decode.regfile.registers_2\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_26546_ _09450_ _09623_ VGND VGND VPWR VPWR _09625_ sky130_fd_sc_hd__nand2_1
X_14560_ _10602_ VGND VGND VPWR VPWR _10603_ sky130_fd_sc_hd__buf_4
X_23758_ _06119_ net1688 _08030_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13511_ csr.io_mem_pc\[2\] VGND VGND VPWR VPWR _09891_ sky130_fd_sc_hd__buf_4
X_22709_ net2689 _07235_ _07243_ _07234_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__o211a_1
X_29265_ clknet_leaf_224_clock _02278_ VGND VGND VPWR VPWR decode.regfile.registers_0\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26477_ _09381_ _09579_ VGND VGND VPWR VPWR _09585_ sky130_fd_sc_hd__nand2_1
X_14491_ net463 _10533_ _10541_ _10535_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__o211a_1
X_23689_ net960 _10881_ _07992_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28216_ clknet_leaf_84_clock net1951 VGND VGND VPWR VPWR csr.mscratch\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16230_ _11435_ decode.regfile.registers_24\[24\] _11244_ _11080_ _11079_ VGND VGND
+ VPWR VPWR _12203_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25428_ _08962_ _08946_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_222_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29196_ clknet_leaf_245_clock _02209_ VGND VGND VPWR VPWR fetch.btb.btbTable\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28147_ clknet_leaf_195_clock _01169_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16161_ _10957_ decode.regfile.registers_22\[22\] _11450_ _10978_ _10990_ VGND VGND
+ VPWR VPWR _12136_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_3_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25359_ _08914_ _08907_ VGND VGND VPWR VPWR _08915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15112_ _11108_ VGND VGND VPWR VPWR _11109_ sky130_fd_sc_hd__clkbuf_4
X_28078_ clknet_leaf_216_clock _01100_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_131_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16092_ _11378_ _12067_ _12068_ VGND VGND VPWR VPWR _12069_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27029_ clknet_leaf_333_clock _00058_ VGND VGND VPWR VPWR decode.regfile.registers_23\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_15043_ _10994_ _10981_ _11039_ VGND VGND VPWR VPWR _11040_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19920_ _05161_ _05169_ _03854_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19851_ _03829_ net349 _03810_ _05098_ net188 VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__a32oi_4
X_18802_ _04098_ _03796_ _03706_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__a21oi_2
X_19782_ _04297_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__clkbuf_8
X_16994_ decode.regfile.registers_22\[5\] _12528_ _12953_ _12687_ VGND VGND VPWR VPWR
+ _12954_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_129_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18733_ net126 _03664_ _04031_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_30_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15945_ _11045_ decode.regfile.registers_12\[16\] _10649_ _11051_ _10631_ VGND VGND
+ VPWR VPWR _11926_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_218_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18664_ _03948_ _03960_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__o21ai_2
X_15876_ _11858_ decode.regfile.registers_17\[14\] _11356_ VGND VGND VPWR VPWR _11859_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _13081_ _13168_ decode.regfile.registers_23\[20\] _13041_ VGND VGND VPWR
+ VPWR _03022_ sky130_fd_sc_hd__or4_1
XFILLER_0_188_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14827_ _10765_ _10869_ VGND VGND VPWR VPWR _10870_ sky130_fd_sc_hd__or2_1
X_18595_ _03887_ _03893_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__and2_2
XFILLER_0_153_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17546_ _12486_ VGND VGND VPWR VPWR _13492_ sky130_fd_sc_hd__clkbuf_4
X_14758_ _10800_ net282 VGND VGND VPWR VPWR _10801_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13709_ _10058_ _10016_ VGND VGND VPWR VPWR _10059_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17477_ _12729_ _13423_ _13424_ VGND VGND VPWR VPWR _13425_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_28_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14689_ decode.id_ex_pc_reg\[23\] VGND VGND VPWR VPWR _10732_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19216_ _04509_ _04511_ _04475_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__o21a_1
X_16428_ _12385_ _12395_ _11184_ decode.regfile.registers_10\[29\] VGND VGND VPWR
+ VPWR _12396_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_60_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19147_ _04394_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__clkbuf_4
X_16359_ _12327_ _12328_ VGND VGND VPWR VPWR _12329_ sky130_fd_sc_hd__nand2_2
XFILLER_0_27_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19078_ decode.id_ex_rs1_data_reg\[9\] _03689_ _04133_ _03701_ _04136_ VGND VGND
+ VPWR VPWR _04376_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_112_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18029_ _12499_ _12490_ _12512_ decode.regfile.registers_12\[31\] _12745_ VGND VGND
+ VPWR VPWR _03425_ sky130_fd_sc_hd__o32a_1
XFILLER_0_61_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21040_ _06005_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout227 net95 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_4
XFILLER_0_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22991_ _07076_ _07433_ _07435_ _07437_ VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__o22a_1
X_24730_ _08549_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21942_ _06568_ _06493_ _06566_ _06569_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24661_ net911 execute.io_target_pc\[19\] _08508_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__mux2_1
X_21873_ net2708 _06521_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26400_ net1545 _09534_ _09539_ _09540_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23612_ _07940_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_167_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20824_ net130 _05879_ _05887_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27380_ clknet_leaf_15_clock _00409_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[21\]
+ sky130_fd_sc_hd__dfxtp_2
X_24592_ net1853 VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26331_ net549 _09491_ _09500_ _09499_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23543_ net79 _07903_ _07914_ _07907_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__o211a_1
X_20755_ _05846_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29050_ clknet_leaf_129_clock _02063_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23474_ net16 _07861_ _07874_ _07865_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__o211a_2
XFILLER_0_18_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26262_ _09392_ _09459_ VGND VGND VPWR VPWR _09461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_210_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20686_ _03728_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_210_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_210_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28001_ clknet_leaf_204_clock _01023_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25213_ _08835_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__clkbuf_1
X_22425_ fetch.bht.bhtTable_tag\[4\]\[12\] fetch.bht.bhtTable_tag\[5\]\[12\] _06878_
+ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26193_ net2571 _09395_ _09414_ _09394_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22356_ _06948_ _06672_ _06950_ _06640_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25144_ net92 _07348_ _07399_ _03580_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__a211o_2
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21307_ _06163_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25075_ _08764_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__clkbuf_1
X_22287_ fetch.bht.bhtTable_tag\[8\]\[11\] fetch.bht.bhtTable_tag\[9\]\[11\] fetch.bht.bhtTable_tag\[10\]\[11\]
+ fetch.bht.bhtTable_tag\[11\]\[11\] _06754_ _06675_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__mux4_1
X_24026_ _08184_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__clkbuf_1
X_28903_ clknet_leaf_112_clock _01916_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_208_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21238_ net943 _06117_ _09912_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__mux2_1
Xhold270 decode.regfile.registers_26\[8\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
X_29883_ clknet_leaf_305_clock _02896_ VGND VGND VPWR VPWR decode.regfile.registers_20\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_208_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold281 decode.regfile.registers_31\[6\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_208_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold292 decode.regfile.registers_17\[15\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28834_ clknet_leaf_135_clock _01847_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21169_ _06074_ _06070_ net548 VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_161_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28765_ clknet_leaf_179_clock _01778_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_13991_ net1366 _10243_ _10253_ _10249_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__o211a_1
X_25977_ net2345 _09243_ _09282_ _09277_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15730_ _11074_ _11687_ _11715_ _11716_ VGND VGND VPWR VPWR _11717_ sky130_fd_sc_hd__a22o_1
X_27716_ clknet_leaf_20_clock _00745_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24928_ net2304 _08665_ _06318_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__a21oi_1
X_28696_ clknet_leaf_121_clock _01709_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27647_ clknet_leaf_45_clock _00676_ VGND VGND VPWR VPWR execute.io_reg_pc\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15661_ _11094_ _11119_ _11093_ _11101_ decode.regfile.registers_20\[9\] VGND VGND
+ VPWR VPWR _11649_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24859_ _08617_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_110 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_132 _10662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17400_ _12611_ _13348_ _13349_ VGND VGND VPWR VPWR _13350_ sky130_fd_sc_hd__o21ai_1
X_14612_ _10654_ VGND VGND VPWR VPWR _10655_ sky130_fd_sc_hd__buf_6
XANTENNA_143 decode.id_ex_rs2_data_reg\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18380_ _03676_ _03677_ _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__nand3_1
X_27578_ clknet_leaf_160_clock _00607_ VGND VGND VPWR VPWR csr.io_mem_pc\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _11143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15592_ decode.regfile.registers_4\[7\] _11375_ _11577_ _11581_ VGND VGND VPWR VPWR
+ _11582_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_120_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29317_ clknet_leaf_228_clock _02330_ VGND VGND VPWR VPWR decode.regfile.registers_2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_17331_ _12874_ _13280_ _13281_ _13282_ VGND VGND VPWR VPWR _13283_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14543_ _10580_ _10583_ decode.control.io_opcode\[3\] _10585_ VGND VGND VPWR VPWR
+ _10586_ sky130_fd_sc_hd__o2bb2a_1
X_26529_ _09434_ _09602_ VGND VGND VPWR VPWR _09614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29248_ clknet_leaf_235_clock _02261_ VGND VGND VPWR VPWR decode.regfile.registers_0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_17262_ _13215_ decode.regfile.registers_28\[11\] _13093_ VGND VGND VPWR VPWR _13216_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14474_ _10081_ _10530_ VGND VGND VPWR VPWR _10532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19001_ _04299_ decode.id_ex_aluop_reg\[1\] decode.id_ex_aluop_reg\[3\] decode.id_ex_aluop_reg\[2\]
+ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__or4b_1
XFILLER_0_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16213_ _11194_ decode.regfile.registers_12\[23\] decode.regfile.registers_13\[23\]
+ _11196_ _11198_ VGND VGND VPWR VPWR _12187_ sky130_fd_sc_hd__o221a_1
XFILLER_0_181_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29179_ clknet_leaf_167_clock _02192_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_141_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17193_ _13141_ _13147_ _12726_ VGND VGND VPWR VPWR _13148_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16144_ _10988_ _11113_ _11119_ _12119_ VGND VGND VPWR VPWR _12120_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16075_ _11646_ _11834_ _11944_ decode.regfile.registers_29\[19\] _12052_ VGND VGND
+ VPWR VPWR _12053_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_90_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15026_ _10657_ _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__a31o_1
X_19903_ _04317_ _05171_ _04985_ _04537_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_220_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19834_ _03811_ _03829_ _05079_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_127_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1909 execute.csr_write_data_out_reg\[21\] VGND VGND VPWR VPWR net2136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19765_ _04508_ _04415_ _04654_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__and3_1
X_16977_ decode.regfile.registers_2\[5\] _10615_ _12729_ VGND VGND VPWR VPWR _12937_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 net380 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15928_ _11761_ net438 _11875_ _11909_ _11760_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__o221a_1
X_18716_ _03796_ _04012_ decode.id_ex_immsrc_reg VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__a21oi_4
X_19696_ _04189_ _03894_ _04972_ _04957_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18647_ decode.id_ex_rs2_data_reg\[21\] net199 _03940_ net258 VGND VGND VPWR VPWR
+ _03946_ sky130_fd_sc_hd__o22a_1
X_15859_ decode.regfile.registers_0\[14\] VGND VGND VPWR VPWR _11842_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18578_ _03710_ _09931_ _03875_ _03876_ _03735_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17529_ decode.regfile.registers_19\[18\] _10599_ _10589_ _12518_ _12543_ VGND VGND
+ VPWR VPWR _13476_ sky130_fd_sc_hd__o41a_1
XFILLER_0_15_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20540_ csr.mscratch\[14\] _05591_ _05554_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20471_ csr.minstret\[5\] _05574_ _05586_ csr.mcycle\[5\] VGND VGND VPWR VPWR _05626_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22210_ _06804_ _06642_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23190_ _07622_ _07623_ _07624_ _07625_ _07080_ _06637_ VGND VGND VPWR VPWR _07626_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22141_ _06620_ _06735_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_320_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_320_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22072_ fetch.bht.bhtTable_tag\[14\]\[18\] fetch.bht.bhtTable_tag\[15\]\[18\] _06618_
+ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25900_ _08973_ _09198_ VGND VGND VPWR VPWR _09238_ sky130_fd_sc_hd__nand2_1
X_21023_ execute.csr_read_data_out_reg\[2\] _05989_ _05985_ VGND VGND VPWR VPWR _05996_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_199_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26880_ net705 _09809_ _09816_ _09812_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_335_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_335_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25831_ _09198_ VGND VGND VPWR VPWR _09199_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_203_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28550_ clknet_leaf_168_clock _01563_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_25762_ _08910_ _09157_ VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__nand2_1
X_22974_ fetch.bht.bhtTable_target_pc\[8\]\[5\] fetch.bht.bhtTable_target_pc\[9\]\[5\]
+ fetch.bht.bhtTable_target_pc\[10\]\[5\] fetch.bht.bhtTable_target_pc\[11\]\[5\]
+ _07068_ _07110_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__mux4_1
XFILLER_0_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27501_ clknet_leaf_34_clock _00530_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dfxtp_2
X_24713_ _08540_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_195_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21925_ csr._mcycle_T_2\[26\] _06545_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__or2_1
X_28481_ clknet_leaf_221_clock _01494_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_195_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25693_ net2373 _09111_ _09119_ _09115_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27432_ clknet_leaf_51_clock _00461_ VGND VGND VPWR VPWR decode.id_ex_isbranch_reg
+ sky130_fd_sc_hd__dfxtp_1
X_24644_ net1074 execute.io_target_pc\[11\] _08497_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21856_ csr.io_mret_vector\[6\] _10820_ _06040_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_218_Right_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20807_ _05878_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__clkbuf_1
X_27363_ clknet_leaf_30_clock _00392_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_24575_ _08469_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__clkbuf_1
X_21787_ csr.io_csr_write_address\[0\] VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29102_ clknet_leaf_17_clock _02115_ VGND VGND VPWR VPWR csr._mcycle_T_3\[50\] sky130_fd_sc_hd__dfxtp_1
X_26314_ _09489_ VGND VGND VPWR VPWR _09490_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23526_ net226 _07903_ _07905_ _07893_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27294_ clknet_leaf_5_clock _00323_ VGND VGND VPWR VPWR decode.regfile.registers_31\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20738_ _05818_ decode.id_ex_rs1_data_reg\[26\] _03585_ VGND VGND VPWR VPWR _05840_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29033_ clknet_leaf_100_clock _02046_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26245_ net562 _09447_ _09451_ _09440_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__o211a_1
X_23457_ net7 _07861_ _07864_ _07865_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__o211a_2
X_20669_ decode.id_ex_rs1_data_reg\[1\] decode.id_ex_ex_rs1_reg\[1\] _05056_ VGND
+ VGND VPWR VPWR _05796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22408_ _07002_ _06678_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14190_ net1208 _10359_ _10367_ _10357_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26176_ _09402_ _09390_ VGND VGND VPWR VPWR _09403_ sky130_fd_sc_hd__nand2_1
X_23388_ execute.io_target_pc\[29\] _10757_ _10970_ _06037_ VGND VGND VPWR VPWR _07812_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25127_ _06145_ net1110 _08562_ VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22339_ fetch.bht.bhtTable_tag\[0\]\[10\] fetch.bht.bhtTable_tag\[1\]\[10\] _06643_
+ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25058_ _03580_ _08752_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_163_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29935_ clknet_leaf_340_clock _02948_ VGND VGND VPWR VPWR decode.regfile.registers_21\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16900_ _12546_ VGND VGND VPWR VPWR _12862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24009_ net989 execute.io_target_pc\[25\] _07960_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__mux2_1
X_29866_ clknet_leaf_298_clock _02879_ VGND VGND VPWR VPWR decode.regfile.registers_19\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17880_ _12541_ _12722_ _03279_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_228_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16831_ _10598_ _10588_ _12549_ _12776_ VGND VGND VPWR VPWR _12794_ sky130_fd_sc_hd__and4_4
X_28817_ clknet_leaf_104_clock _01830_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_29797_ clknet_leaf_292_clock _02810_ VGND VGND VPWR VPWR decode.regfile.registers_17\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19550_ _04829_ _04831_ _04211_ _04526_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a31o_1
X_28748_ clknet_leaf_109_clock _01761_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16762_ _12725_ VGND VGND VPWR VPWR _12726_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13974_ _10242_ VGND VGND VPWR VPWR _10243_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18501_ _03709_ decode.id_ex_imm_reg\[28\] _03798_ _03799_ VGND VGND VPWR VPWR _03800_
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_219_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15713_ decode.regfile.registers_7\[10\] _11378_ _11170_ decode.regfile.registers_6\[10\]
+ _11166_ VGND VGND VPWR VPWR _11700_ sky130_fd_sc_hd__a221o_1
X_19481_ _04761_ _04764_ _04766_ _04104_ _04425_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__a32o_2
XFILLER_0_198_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28679_ clknet_leaf_115_clock _01692_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16693_ _12657_ VGND VGND VPWR VPWR _12658_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18432_ decode.io_wb_rd\[0\] csr.io_csr_address\[0\] VGND VGND VPWR VPWR _03731_
+ sky130_fd_sc_hd__or2b_1
X_15644_ _11124_ _11631_ _11632_ VGND VGND VPWR VPWR _11633_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18363_ _03660_ _03661_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__nand2_4
XFILLER_0_200_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _11236_ _11562_ _11563_ _11565_ VGND VGND VPWR VPWR _11566_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17314_ decode.regfile.registers_11\[13\] _12878_ VGND VGND VPWR VPWR _13266_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14526_ net410 _10570_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18294_ decode.id_ex_rs2_data_reg\[13\] _03605_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17245_ _13190_ _13198_ _12599_ decode.regfile.registers_10\[11\] VGND VGND VPWR
+ VPWR _13199_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_154_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14457_ _10036_ _10517_ VGND VGND VPWR VPWR _10523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_226_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17176_ _13087_ decode.regfile.registers_26\[9\] _12814_ _13047_ _13088_ VGND VGND
+ VPWR VPWR _13132_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_49_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14388_ _10053_ _10474_ VGND VGND VPWR VPWR _10483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16127_ decode.regfile.registers_2\[21\] _11369_ _11142_ _11110_ VGND VGND VPWR VPWR
+ _12103_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_109_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16058_ decode.regfile.registers_13\[19\] _11276_ _12034_ _12035_ VGND VGND VPWR
+ VPWR _12036_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15009_ _11018_ VGND VGND VPWR VPWR _11019_ sky130_fd_sc_hd__clkbuf_4
Xhold2407 decode.regfile.registers_19\[25\] VGND VGND VPWR VPWR net2634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2418 csr._mcycle_T_2\[3\] VGND VGND VPWR VPWR net2645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2429 decode.id_ex_rs1_data_reg\[25\] VGND VGND VPWR VPWR net2656 sky130_fd_sc_hd__dlygate4sd3_1
X_19817_ _04471_ _04439_ _04509_ _04949_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__a31o_1
Xhold1706 decode.regfile.registers_4\[12\] VGND VGND VPWR VPWR net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1717 fetch.bht.bhtTable_tag\[15\]\[12\] VGND VGND VPWR VPWR net1944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1728 decode.io_id_pc\[13\] VGND VGND VPWR VPWR net1955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 decode.regfile.registers_3\[13\] VGND VGND VPWR VPWR net1966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19748_ _03912_ _04863_ _04935_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19679_ _04932_ _04192_ _04191_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_32_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21710_ csr.minstret\[20\] csr.minstret\[21\] csr.minstret\[22\] VGND VGND VPWR VPWR
+ _06411_ sky130_fd_sc_hd__and3_1
X_22690_ net2692 _07222_ _07232_ _07221_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21641_ csr.minstret\[12\] _06338_ _06355_ _06329_ csr._mcycle_T_2\[13\] VGND VGND
+ VPWR VPWR _06357_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_190_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24360_ net2098 execute.io_target_pc\[3\] _08356_ VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__mux2_1
X_21572_ _06143_ net1191 _06306_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_10 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_21 _05621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_32 _09954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23311_ net221 net222 net223 _07716_ VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__and4_1
XANTENNA_43 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20523_ net924 _05671_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__nor2_1
X_24291_ _08053_ net1759 _06210_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_915 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_54 _10598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _11012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_76 _11100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26030_ _08952_ _09310_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__nand2_1
XANTENNA_87 decode.id_ex_rs1_data_reg\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23242_ net224 _07536_ _07537_ _07675_ _07535_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__o311a_1
X_20454_ csr.mcycle\[3\] _05537_ _05601_ _05610_ _03595_ VGND VGND VPWR VPWR _00690_
+ sky130_fd_sc_hd__o221a_1
XANTENNA_98 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_41_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23173_ _07406_ _07605_ _07097_ _07609_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20385_ _05531_ _05546_ net2764 VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22124_ net225 _06698_ _06717_ _06718_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27981_ clknet_leaf_195_clock _01003_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput150 net150 VGND VGND VPWR VPWR io_memory_write_data[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput161 net161 VGND VGND VPWR VPWR io_memory_write_data[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29720_ clknet_leaf_311_clock _02733_ VGND VGND VPWR VPWR decode.regfile.registers_14\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_274_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_274_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22055_ _06649_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__buf_4
X_26932_ net1209 _09839_ _09846_ _09836_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_1 _00550_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21006_ net2724 _05977_ _05985_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_197_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29651_ clknet_leaf_279_clock _02664_ VGND VGND VPWR VPWR decode.regfile.registers_12\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_26863_ _09389_ _09806_ VGND VGND VPWR VPWR _09807_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_197_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28602_ clknet_leaf_129_clock _01615_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_25814_ _08962_ _09179_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29582_ clknet_leaf_275_clock _02595_ VGND VGND VPWR VPWR decode.regfile.registers_10\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26794_ net503 _09766_ _09767_ _09758_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_289_clock clknet_5_18__leaf_clock VGND VGND VPWR VPWR clknet_leaf_289_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_3_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28533_ clknet_leaf_216_clock _01546_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25745_ _08968_ _09110_ VGND VGND VPWR VPWR _09149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22957_ _07371_ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__buf_4
XFILLER_0_211_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28464_ clknet_leaf_138_clock _01477_ VGND VGND VPWR VPWR decode.io_id_pc\[22\] sky130_fd_sc_hd__dfxtp_1
X_21908_ _06542_ _06543_ _06544_ _06546_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__o211a_1
X_13690_ _10042_ _10016_ VGND VGND VPWR VPWR _10043_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_3_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_3_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25676_ net1863 _09069_ _09108_ _09100_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__o211a_1
X_22888_ net1813 _10777_ _07335_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_212_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_212_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27415_ clknet_leaf_15_clock _00444_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[24\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_194_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24627_ net1244 execute.io_target_pc\[3\] _07308_ VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__mux2_1
X_28395_ clknet_leaf_142_clock _01408_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_4
X_21839_ net559 _06497_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15360_ _10650_ _11111_ _11117_ VGND VGND VPWR VPWR _11355_ sky130_fd_sc_hd__and3_1
X_27346_ clknet_leaf_43_clock _00375_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[19\]
+ sky130_fd_sc_hd__dfxtp_2
X_24558_ _08460_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14311_ net535 _10434_ _10438_ _10427_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23509_ net94 _07889_ _07895_ _07893_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27277_ clknet_leaf_9_clock _00306_ VGND VGND VPWR VPWR decode.regfile.registers_30\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_15291_ _11286_ VGND VGND VPWR VPWR _11287_ sky130_fd_sc_hd__buf_2
X_24489_ _08049_ net1942 _07276_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_227_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_227_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29016_ clknet_leaf_122_clock _02029_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_17030_ decode.regfile.registers_17\[6\] _12580_ _12826_ _12988_ VGND VGND VPWR VPWR
+ _12989_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14242_ net2078 _10390_ _10397_ _10398_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__o211a_1
X_26228_ _09438_ _09372_ VGND VGND VPWR VPWR _09439_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14173_ net1088 _10346_ _10358_ _10357_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__o211a_1
X_26159_ _09389_ _09390_ VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_186_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18981_ _04279_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ _03329_ _12695_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__a21o_1
X_29918_ clknet_leaf_334_clock _02931_ VGND VGND VPWR VPWR decode.regfile.registers_21\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17863_ _13451_ net2788 _13492_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__o21a_1
X_29849_ clknet_leaf_310_clock _02862_ VGND VGND VPWR VPWR decode.regfile.registers_18\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19602_ _04805_ _04370_ _04729_ _04883_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__a31o_1
XFILLER_0_191_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16814_ decode.regfile.registers_8\[2\] _12776_ _12550_ _12604_ _12607_ VGND VGND
+ VPWR VPWR _12777_ sky130_fd_sc_hd__a41o_1
XFILLER_0_191_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17794_ _12498_ _12540_ _12977_ decode.regfile.registers_7\[25\] _12645_ VGND VGND
+ VPWR VPWR _03196_ sky130_fd_sc_hd__o32a_1
XFILLER_0_156_1343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19533_ _04626_ _04816_ _04349_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__mux2_1
X_16745_ _12708_ VGND VGND VPWR VPWR _12709_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13957_ _10112_ _10223_ VGND VGND VPWR VPWR _10233_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19464_ _04332_ _04284_ _04317_ _04287_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__o211a_1
X_16676_ _12632_ _12634_ _12640_ VGND VGND VPWR VPWR _12641_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_200 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13888_ net568 _10180_ _10191_ _10188_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_211 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_222 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15627_ decode.regfile.registers_1\[8\] _11117_ _11057_ _11109_ VGND VGND VPWR VPWR
+ _11616_ sky130_fd_sc_hd__and4_1
X_18415_ _03711_ _03712_ _09921_ _03713_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__o211ai_4
XINSDIODE1_233 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19395_ _04165_ _04167_ _04663_ _04683_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_185_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_244 net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_255 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_266 _06422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18346_ execute.io_mem_rd\[2\] decode.id_ex_ex_rs1_reg\[2\] VGND VGND VPWR VPWR _03645_
+ sky130_fd_sc_hd__or2b_4
XINSDIODE1_277 _11012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15558_ _11535_ _11545_ _11548_ VGND VGND VPWR VPWR _11549_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_173_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_288 _12504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_299 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14509_ _09879_ _09882_ _10551_ _10553_ VGND VGND VPWR VPWR _10554_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18277_ decode.id_ex_rs2_data_reg\[5\] _03596_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__and2_1
X_15489_ decode.regfile.registers_23\[4\] _11088_ _11451_ _11481_ VGND VGND VPWR VPWR
+ _11482_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17228_ _12492_ VGND VGND VPWR VPWR _13182_ sky130_fd_sc_hd__clkbuf_4
Xinput30 net737 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput41 io_memory_read_data[16] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput52 io_memory_read_data[26] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
XFILLER_0_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput63 io_memory_read_data[7] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
XFILLER_0_130_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold803 decode.regfile.registers_23\[6\] VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold814 decode.regfile.registers_18\[8\] VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ decode.regfile.registers_11\[9\] _12724_ _12722_ _12540_ VGND VGND VPWR VPWR
+ _13115_ sky130_fd_sc_hd__o2bb2a_1
Xhold825 fetch.bht.bhtTable_tag\[8\]\[18\] VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 fetch.bht.bhtTable_target_pc\[12\]\[0\] VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold847 fetch.bht.bhtTable_target_pc\[12\]\[11\] VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 fetch.bht.bhtTable_tag\[5\]\[15\] VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__dlygate4sd3_1
X_20170_ _05370_ _05372_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__xnor2_1
Xhold869 fetch.bht.bhtTable_tag\[12\]\[4\] VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2204 decode.regfile.registers_9\[14\] VGND VGND VPWR VPWR net2431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2215 fetch.btb.btbTable\[2\]\[1\] VGND VGND VPWR VPWR net2442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2226 decode.regfile.registers_24\[31\] VGND VGND VPWR VPWR net2453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2237 decode.regfile.registers_25\[29\] VGND VGND VPWR VPWR net2464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1503 decode.regfile.registers_25\[25\] VGND VGND VPWR VPWR net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2248 decode.regfile.registers_22\[4\] VGND VGND VPWR VPWR net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_7__f_clock clknet_2_0_0_clock VGND VGND VPWR VPWR clknet_5_7__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
Xhold1514 fetch.bht.bhtTable_tag\[15\]\[8\] VGND VGND VPWR VPWR net1741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2259 decode.regfile.registers_20\[27\] VGND VGND VPWR VPWR net2486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1525 decode.regfile.registers_10\[31\] VGND VGND VPWR VPWR net1752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1536 fetch.bht.bhtTable_target_pc\[5\]\[22\] VGND VGND VPWR VPWR net1763 sky130_fd_sc_hd__dlygate4sd3_1
X_23860_ _08094_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__clkbuf_1
Xhold1547 decode.regfile.registers_10\[14\] VGND VGND VPWR VPWR net1774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1558 execute.csr_write_data_out_reg\[5\] VGND VGND VPWR VPWR net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1569 decode.regfile.registers_26\[16\] VGND VGND VPWR VPWR net1796 sky130_fd_sc_hd__dlygate4sd3_1
X_22811_ net781 _10800_ _07297_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23791_ _06153_ net1145 _08041_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_192_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25530_ _09023_ VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__buf_2
X_22742_ _07263_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25461_ net2398 _08979_ _08985_ _08972_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22673_ csr._mcycle_T_2\[12\] _07223_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27200_ clknet_leaf_361_clock _00229_ VGND VGND VPWR VPWR decode.regfile.registers_28\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_24412_ _08383_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28180_ clknet_leaf_60_clock _01202_ VGND VGND VPWR VPWR csr.io_mret_vector\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_21624_ net2483 _06317_ csr.minstret\[7\] _05856_ _06345_ VGND VGND VPWR VPWR _01124_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_47_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25392_ _08937_ _08923_ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27131_ clknet_leaf_359_clock _00160_ VGND VGND VPWR VPWR decode.regfile.registers_26\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24343_ _08105_ net1175 _06187_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__mux2_1
X_21555_ _06126_ net1754 _06295_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27062_ clknet_leaf_330_clock _00091_ VGND VGND VPWR VPWR decode.regfile.registers_24\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20506_ _05439_ _05656_ _03449_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__and3b_1
X_24274_ _08312_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__clkbuf_1
X_21486_ _06115_ net2132 _06252_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26013_ _08935_ _09297_ VGND VGND VPWR VPWR _09304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23225_ _07655_ _07657_ _07111_ _07658_ _07075_ VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__o221a_1
X_20437_ _05534_ _05526_ _05536_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__and3_2
XFILLER_0_120_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23156_ fetch.bht.bhtTable_target_pc\[12\]\[15\] fetch.bht.bhtTable_target_pc\[13\]\[15\]
+ fetch.bht.bhtTable_target_pc\[14\]\[15\] fetch.bht.bhtTable_target_pc\[15\]\[15\]
+ _07107_ _07114_ VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__mux4_1
X_20368_ _05518_ _05522_ _05530_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_149_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22107_ fetch.bht.bhtTable_tag\[0\]\[3\] fetch.bht.bhtTable_tag\[1\]\[3\] _06680_
+ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23087_ _07085_ _07524_ _07526_ _07528_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__a2bb2o_2
X_27964_ clknet_leaf_223_clock _00986_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_224_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20299_ _05475_ _05219_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_224_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22038_ _06632_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__buf_4
X_29703_ clknet_leaf_284_clock _02716_ VGND VGND VPWR VPWR decode.regfile.registers_14\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26915_ _09956_ VGND VGND VPWR VPWR _09836_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_8_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27895_ clknet_leaf_22_clock _00924_ VGND VGND VPWR VPWR csr._mcycle_T_2\[16\] sky130_fd_sc_hd__dfxtp_2
X_14860_ decode.id_ex_pc_reg\[22\] _10863_ _10866_ _10867_ _10902_ VGND VGND VPWR
+ VPWR _10903_ sky130_fd_sc_hd__o221ai_1
X_29634_ clknet_leaf_287_clock _02647_ VGND VGND VPWR VPWR decode.regfile.registers_12\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_26846_ net2008 _09795_ _09797_ _09784_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__o211a_1
X_13811_ _10060_ memory.io_wb_aluresult\[31\] _10004_ memory.io_wb_readdata\[31\]
+ _10005_ VGND VGND VPWR VPWR _10145_ sky130_fd_sc_hd__a221o_1
X_29565_ clknet_leaf_251_clock _02578_ VGND VGND VPWR VPWR decode.regfile.registers_10\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14791_ decode.id_ex_pc_reg\[2\] VGND VGND VPWR VPWR _10834_ sky130_fd_sc_hd__clkbuf_4
X_26777_ _09701_ VGND VGND VPWR VPWR _09758_ sky130_fd_sc_hd__clkbuf_4
X_23989_ net1188 execute.io_target_pc\[15\] _08164_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28516_ clknet_leaf_197_clock _01529_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_16530_ _11010_ _12494_ _12491_ _10939_ VGND VGND VPWR VPWR _12495_ sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_151_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_151_clock
+ sky130_fd_sc_hd__clkbuf_8
X_13742_ _10086_ VGND VGND VPWR VPWR _10087_ sky130_fd_sc_hd__buf_6
X_25728_ _08952_ _09136_ VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29496_ clknet_leaf_249_clock _02509_ VGND VGND VPWR VPWR decode.regfile.registers_7\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28447_ clknet_leaf_144_clock _01460_ VGND VGND VPWR VPWR decode.io_id_pc\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16461_ _12421_ _12427_ _11289_ VGND VGND VPWR VPWR _12428_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25659_ _08990_ VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__buf_4
X_13673_ _09946_ _09947_ memory.io_wb_reg_pc\[10\] VGND VGND VPWR VPWR _10028_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_175_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18200_ decode.control.io_funct7\[5\] _03523_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_175_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15412_ _11354_ VGND VGND VPWR VPWR _11406_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_182_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19180_ _04349_ _04471_ _04475_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__o21ai_2
X_28378_ clknet_leaf_190_clock _01391_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16392_ _11134_ _12359_ _12360_ VGND VGND VPWR VPWR _12361_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_117_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_166_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_166_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18131_ _03482_ _03493_ _03487_ net2236 VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_108_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27329_ clknet_leaf_55_clock _00358_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15343_ _10958_ decode.regfile.registers_26\[1\] _11261_ _11338_ _10992_ VGND VGND
+ VPWR VPWR _11339_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_54_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18062_ _10965_ _10964_ _10951_ _10582_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_0_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15274_ _10651_ _10633_ _10640_ _11111_ VGND VGND VPWR VPWR _11270_ sky130_fd_sc_hd__and4_1
XFILLER_0_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17013_ decode.regfile.registers_4\[6\] _12549_ _12532_ decode.regfile.registers_5\[6\]
+ _12615_ VGND VGND VPWR VPWR _12972_ sky130_fd_sc_hd__a221oi_2
X_14225_ _10025_ _10387_ VGND VGND VPWR VPWR _10389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14156_ _10042_ _10342_ VGND VGND VPWR VPWR _10349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14087_ _10058_ _10299_ VGND VGND VPWR VPWR _10309_ sky130_fd_sc_hd__nand2_1
X_18964_ _04262_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_104_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_37_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _03311_ _03312_ _03313_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_143_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18895_ _03872_ _03881_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__nor2_1
XFILLER_0_193_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17846_ _10595_ _10599_ _10588_ _12542_ _03246_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_33_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14989_ _11005_ VGND VGND VPWR VPWR _11006_ sky130_fd_sc_hd__clkbuf_4
X_17777_ _12968_ _03177_ _03178_ _03179_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_119_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_119_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_221_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19516_ _04602_ _04291_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16728_ _12500_ _12507_ _12517_ _12692_ VGND VGND VPWR VPWR _12693_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_88_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19447_ _04733_ _04690_ _04248_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16659_ decode.regfile.registers_4\[0\] _12618_ _12620_ decode.regfile.registers_5\[0\]
+ _12623_ VGND VGND VPWR VPWR _12624_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19378_ _04503_ _04137_ _04667_ _04143_ _04142_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18329_ _03630_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21340_ net854 _10759_ _06179_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21271_ _10773_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold600 fetch.bht.bhtTable_target_pc\[1\]\[5\] VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold611 decode.regfile.registers_22\[13\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_1286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold622 decode.regfile.registers_4\[9\] VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 fetch.bht.bhtTable_target_pc\[3\]\[26\] VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__dlygate4sd3_1
X_23010_ _07454_ _07455_ _07076_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20222_ _05415_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__buf_2
Xhold644 fetch.bht.bhtTable_target_pc\[11\]\[29\] VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold655 _01233_ VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold666 decode.regfile.registers_29\[26\] VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 decode.regfile.registers_24\[10\] VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 fetch.bht.bhtTable_target_pc\[11\]\[2\] VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__dlygate4sd3_1
X_20153_ _05350_ _05356_ _05357_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold699 decode.regfile.registers_2\[12\] VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2001 decode.regfile.registers_29\[8\] VGND VGND VPWR VPWR net2228 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2012 decode.regfile.registers_6\[30\] VGND VGND VPWR VPWR net2239 sky130_fd_sc_hd__dlygate4sd3_1
X_20084_ _05283_ _05292_ _05298_ _05289_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_5_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2023 decode.regfile.registers_21\[0\] VGND VGND VPWR VPWR net2250 sky130_fd_sc_hd__dlygate4sd3_1
X_24961_ csr._mcycle_T_3\[55\] csr._mcycle_T_3\[54\] csr._mcycle_T_3\[53\] _08682_
+ VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__and4_1
Xhold2034 decode.regfile.registers_9\[2\] VGND VGND VPWR VPWR net2261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1300 fetch.bht.bhtTable_target_pc\[9\]\[3\] VGND VGND VPWR VPWR net1527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2045 decode.regfile.registers_30\[18\] VGND VGND VPWR VPWR net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 fetch.bht.bhtTable_tag\[15\]\[15\] VGND VGND VPWR VPWR net1538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2056 decode.regfile.registers_26\[27\] VGND VGND VPWR VPWR net2283 sky130_fd_sc_hd__dlygate4sd3_1
X_26700_ net1638 _09709_ _09713_ _09702_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__o211a_1
X_23912_ net1082 _08070_ _08119_ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__mux2_1
Xhold1322 decode.regfile.registers_25\[20\] VGND VGND VPWR VPWR net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2067 decode.regfile.registers_9\[4\] VGND VGND VPWR VPWR net2294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27680_ clknet_leaf_27_clock _00709_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1333 fetch.bht.bhtTable_target_pc\[15\]\[27\] VGND VGND VPWR VPWR net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2078 decode.io_id_pc\[17\] VGND VGND VPWR VPWR net2305 sky130_fd_sc_hd__dlygate4sd3_1
X_24892_ csr.mcycle\[21\] csr.mcycle\[24\] _08640_ VGND VGND VPWR VPWR _08641_ sky130_fd_sc_hd__and3_1
Xhold2089 decode.regfile.registers_26\[21\] VGND VGND VPWR VPWR net2316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1344 decode.regfile.registers_30\[30\] VGND VGND VPWR VPWR net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1355 decode.regfile.registers_23\[20\] VGND VGND VPWR VPWR net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 decode.regfile.registers_12\[28\] VGND VGND VPWR VPWR net1593 sky130_fd_sc_hd__dlygate4sd3_1
X_26631_ _09385_ _09666_ VGND VGND VPWR VPWR _09673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_224_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23843_ execute.io_target_pc\[16\] VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__buf_2
Xhold1377 fetch.bht.bhtTable_tag\[10\]\[3\] VGND VGND VPWR VPWR net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1388 fetch.bht.bhtTable_tag\[11\]\[8\] VGND VGND VPWR VPWR net1615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1399 fetch.bht.bhtTable_target_pc\[5\]\[13\] VGND VGND VPWR VPWR net1626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29350_ clknet_leaf_257_clock _02363_ VGND VGND VPWR VPWR decode.regfile.registers_3\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26562_ net613 _09622_ _09633_ _09619_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__o211a_1
X_23774_ _06136_ net916 _08030_ VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20986_ execute.io_reg_pc\[18\] _05965_ _05973_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__and3_1
X_28301_ clknet_leaf_164_clock _00011_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25513_ _08964_ _09005_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29281_ clknet_leaf_241_clock _02294_ VGND VGND VPWR VPWR decode.regfile.registers_1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_22725_ _10913_ _07248_ _07254_ _10916_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_149_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26493_ _09398_ _09589_ VGND VGND VPWR VPWR _09594_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_83_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_83_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_217_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28232_ clknet_leaf_73_clock _01254_ VGND VGND VPWR VPWR csr._minstret_T_3\[32\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_48_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25444_ _08973_ _08905_ VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22656_ net1370 _07210_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21607_ _06332_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__buf_2
X_28163_ clknet_leaf_69_clock net513 VGND VGND VPWR VPWR csr._csr_read_data_T_9\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25375_ _08925_ _08923_ VGND VGND VPWR VPWR _08926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22587_ csr._minstret_T_3\[43\] csr._minstret_T_3\[42\] csr._minstret_T_3\[41\] _07160_
+ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_170_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27114_ clknet_leaf_347_clock _00143_ VGND VGND VPWR VPWR decode.regfile.registers_25\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xclone44 net274 _04104_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__nand2_1
X_24326_ _08339_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28094_ clknet_leaf_184_clock _01116_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21538_ _06109_ net2164 _06284_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_98_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_98_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_211_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27045_ clknet_leaf_342_clock _00074_ VGND VGND VPWR VPWR decode.regfile.registers_23\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_24257_ _08085_ net1828 _08300_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__mux2_1
X_21469_ _10557_ _09900_ _09916_ _10556_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_50_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_226_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14010_ net1471 _10258_ _10264_ _10262_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__o211a_1
X_23208_ fetch.bht.bhtTable_target_pc\[10\]\[18\] fetch.bht.bhtTable_target_pc\[11\]\[18\]
+ _07067_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24188_ _08268_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_21_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23139_ _07577_ _07082_ VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__and2_1
XFILLER_0_222_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28996_ clknet_leaf_128_clock _02009_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15961_ _11761_ net399 _11910_ _11941_ _11760_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__o221a_1
X_27947_ clknet_leaf_204_clock _00969_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14912_ decode.control.io_funct3\[1\] VGND VGND VPWR VPWR _10943_ sky130_fd_sc_hd__buf_2
X_17700_ _12968_ _03102_ _03103_ _03104_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__a31o_1
X_27878_ clknet_leaf_65_clock _00907_ VGND VGND VPWR VPWR csr.io_ecause\[1\] sky130_fd_sc_hd__dfxtp_1
X_15892_ _11761_ net431 _11833_ _11874_ _11760_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18680_ net229 net233 _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_106_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_36_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_106_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14843_ _10721_ _10813_ _10882_ VGND VGND VPWR VPWR _10886_ sky130_fd_sc_hd__and3_1
X_17631_ decode.regfile.registers_2\[21\] _12634_ _12629_ _03036_ VGND VGND VPWR VPWR
+ _03037_ sky130_fd_sc_hd__o211ai_4
X_29617_ clknet_leaf_279_clock _02630_ VGND VGND VPWR VPWR decode.regfile.registers_11\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_26829_ _09432_ _09776_ VGND VGND VPWR VPWR _09787_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_177_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17562_ decode.regfile.registers_12\[19\] _12542_ _12723_ _12659_ _02969_ VGND VGND
+ VPWR VPWR _02970_ sky130_fd_sc_hd__o311a_1
XFILLER_0_59_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14774_ csr.io_mem_pc\[9\] VGND VGND VPWR VPWR _10817_ sky130_fd_sc_hd__buf_4
X_29548_ clknet_leaf_274_clock _02561_ VGND VGND VPWR VPWR decode.regfile.registers_9\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19301_ _04280_ _04282_ _04592_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__o31a_1
X_16513_ _11050_ _11090_ decode.regfile.registers_25\[31\] _12452_ _12478_ VGND VGND
+ VPWR VPWR _12479_ sky130_fd_sc_hd__o32a_1
XFILLER_0_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13725_ _10003_ memory.io_wb_aluresult\[18\] _10004_ memory.io_wb_readdata\[18\]
+ _10005_ VGND VGND VPWR VPWR _10072_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17493_ decode.regfile.registers_23\[17\] _12714_ _13416_ _13440_ _12515_ VGND VGND
+ VPWR VPWR _13441_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29479_ clknet_leaf_269_clock _02492_ VGND VGND VPWR VPWR decode.regfile.registers_7\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19232_ _04034_ _04055_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__or2_1
X_16444_ _11075_ _12410_ _12411_ _11486_ VGND VGND VPWR VPWR _12412_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13656_ _10012_ memory.io_wb_aluresult\[8\] _09981_ memory.io_wb_readdata\[8\] _09995_
+ VGND VGND VPWR VPWR _10013_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19163_ _04423_ _04441_ _04458_ _04459_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__o31a_2
XFILLER_0_183_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16375_ _10961_ _11834_ _11944_ decode.regfile.registers_29\[27\] _12344_ VGND VGND
+ VPWR VPWR _12345_ sky130_fd_sc_hd__o221a_1
XFILLER_0_183_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13587_ _09950_ _09951_ VGND VGND VPWR VPWR _09952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18114_ _03484_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15326_ _11124_ _11320_ _11321_ VGND VGND VPWR VPWR _11322_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19094_ _03637_ _04056_ _04391_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__and3_2
XFILLER_0_87_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18045_ _12494_ decode.regfile.registers_26\[31\] _13002_ _11010_ _11026_ VGND VGND
+ VPWR VPWR _03441_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_53_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15257_ _11252_ VGND VGND VPWR VPWR _11253_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_197_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14208_ net601 _10376_ _10379_ _10369_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15188_ _10660_ _10655_ _11143_ VGND VGND VPWR VPWR _11185_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14139_ _09993_ _10333_ VGND VGND VPWR VPWR _10339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19996_ net788 decode.id_ex_pc_reg\[0\] VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_25__f_clock clknet_2_3_0_clock VGND VGND VPWR VPWR clknet_5_25__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_226_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18947_ _03990_ _03991_ _03996_ _03706_ decode.id_ex_imm_reg\[1\] VGND VGND VPWR
+ VPWR _04246_ sky130_fd_sc_hd__a32o_2
XFILLER_0_207_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18878_ _04137_ _04141_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_206_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17829_ decode.regfile.registers_8\[26\] _12889_ _12607_ VGND VGND VPWR VPWR _03230_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20840_ _05896_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20771_ _05854_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22510_ fetch.bht.bhtTable_target_pc\[8\]\[1\] fetch.bht.bhtTable_target_pc\[9\]\[1\]
+ fetch.bht.bhtTable_target_pc\[10\]\[1\] fetch.bht.bhtTable_target_pc\[11\]\[1\]
+ _07099_ _07103_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23490_ decode.control.io_funct7\[5\] _07876_ _07873_ VGND VGND VPWR VPWR _07884_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22441_ _06641_ _06811_ _06815_ _06819_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_91_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25160_ _10568_ _09894_ VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__nand2_1
X_22372_ fetch.bht.bhtTable_tag\[4\]\[16\] fetch.bht.bhtTable_tag\[5\]\[16\] fetch.bht.bhtTable_tag\[6\]\[16\]
+ fetch.bht.bhtTable_tag\[7\]\[16\] _06878_ _06621_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__mux4_1
XFILLER_0_206_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24111_ _08228_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21323_ net1177 _10800_ _06168_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25091_ _08773_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21254_ net1623 _06128_ _06120_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__mux2_1
X_24042_ net1457 execute.io_target_pc\[9\] _08187_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold430 decode.regfile.registers_12\[4\] VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 decode.regfile.registers_30\[21\] VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold452 decode.regfile.registers_21\[6\] VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold463 decode.regfile.registers_1\[3\] VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20205_ _05401_ _05402_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap182 net183 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
X_28850_ clknet_leaf_119_clock _01863_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_21185_ _06086_ _06082_ net1269 VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__and3_1
Xhold474 decode.regfile.registers_10\[29\] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold485 decode.regfile.registers_13\[9\] VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap193 _10096_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_221_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold496 csr._mcycle_T_2\[23\] VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__buf_1
XFILLER_0_141_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20136_ _05342_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__xor2_1
X_27801_ clknet_leaf_331_clock _00830_ VGND VGND VPWR VPWR memory.io_wb_readdata\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_28781_ clknet_leaf_99_clock _01794_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25993_ _08914_ _09287_ VGND VGND VPWR VPWR _09293_ sky130_fd_sc_hd__nand2_1
X_27732_ clknet_leaf_70_clock _00761_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20067_ _05282_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__and2b_1
X_24944_ csr._mcycle_T_3\[49\] csr._mcycle_T_3\[48\] _08672_ VGND VGND VPWR VPWR _08676_
+ sky130_fd_sc_hd__and3_1
Xhold1130 fetch.bht.bhtTable_tag\[9\]\[6\] VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 fetch.bht.bhtTable_target_pc\[15\]\[31\] VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1152 fetch.bht.bhtTable_target_pc\[4\]\[14\] VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__dlygate4sd3_1
X_27663_ clknet_leaf_28_clock _00692_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_24875_ _08625_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__clkbuf_1
Xhold1163 fetch.bht.bhtTable_tag\[14\]\[4\] VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1174 fetch.bht.bhtTable_tag\[6\]\[3\] VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 _08197_ VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1196 fetch.bht.bhtTable_target_pc\[2\]\[7\] VGND VGND VPWR VPWR net1423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26614_ net2259 _09623_ _09662_ _09660_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__o211a_1
X_29402_ clknet_leaf_248_clock _02415_ VGND VGND VPWR VPWR decode.regfile.registers_5\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_219_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23826_ _08071_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_219_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27594_ clknet_leaf_147_clock _00623_ VGND VGND VPWR VPWR execute.io_target_pc\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_68_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29333_ clknet_leaf_226_clock _02346_ VGND VGND VPWR VPWR decode.regfile.registers_2\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_26545_ net1729 _09622_ _09624_ _09619_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__o211a_1
X_23757_ _09905_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__clkbuf_8
X_20969_ execute.io_reg_pc\[10\] _05965_ _05961_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _09881_ _09884_ _09885_ _09890_ net395 VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__a41o_1
X_22708_ csr._mcycle_T_2\[28\] _07236_ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_172_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29264_ clknet_leaf_223_clock _02277_ VGND VGND VPWR VPWR decode.regfile.registers_0\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26476_ net2438 _09578_ _09584_ _09582_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__o211a_1
X_14490_ _10117_ _10530_ VGND VGND VPWR VPWR _10541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23688_ _07994_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28215_ clknet_leaf_84_clock net1418 VGND VGND VPWR VPWR csr.mscratch\[17\] sky130_fd_sc_hd__dfxtp_1
X_25427_ net192 VGND VGND VPWR VPWR _08962_ sky130_fd_sc_hd__buf_4
XFILLER_0_180_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22639_ csr._minstret_T_3\[61\] _07202_ _07179_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__a21oi_1
X_29195_ clknet_leaf_163_clock _02208_ VGND VGND VPWR VPWR fetch.btb.btbTable\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28146_ clknet_leaf_198_clock _01168_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_16160_ _10959_ decode.regfile.registers_26\[22\] _11447_ _11348_ _10993_ VGND VGND
+ VPWR VPWR _12135_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_183_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25358_ _09983_ VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15111_ _11107_ VGND VGND VPWR VPWR _11108_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24309_ _08330_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28077_ clknet_leaf_206_clock _01099_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_131_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16091_ decode.regfile.registers_7\[20\] _11378_ _11134_ VGND VGND VPWR VPWR _12068_
+ sky130_fd_sc_hd__a21oi_1
X_25289_ _08869_ decode.regfile.registers_0\[6\] VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27028_ clknet_leaf_333_clock _00057_ VGND VGND VPWR VPWR decode.regfile.registers_23\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_15042_ _11038_ VGND VGND VPWR VPWR _11039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19850_ _03639_ net189 _03803_ _04667_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18801_ _04096_ net355 _03687_ decode.id_ex_rs1_data_reg\[13\] _04099_ VGND VGND
+ VPWR VPWR _04100_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_222_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19781_ _04225_ _04667_ _05050_ _05053_ _05054_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__o221ai_2
X_28979_ clknet_leaf_134_clock _01992_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_16993_ decode.regfile.registers_21\[5\] _12822_ _12924_ _12952_ _12806_ VGND VGND
+ VPWR VPWR _12953_ sky130_fd_sc_hd__o221a_1
XFILLER_0_207_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18732_ execute.csr_read_data_out_reg\[4\] _03658_ execute.io_reg_pc\[4\] _03662_
+ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__o22a_1
XFILLER_0_207_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ _11922_ _11923_ _11924_ VGND VGND VPWR VPWR _11925_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_30_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15875_ decode.regfile.registers_16\[14\] _11123_ _11838_ _11857_ VGND VGND VPWR
+ VPWR _11858_ sky130_fd_sc_hd__o22a_1
X_18663_ _10091_ _03772_ _03961_ _03947_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_125_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _10868_ _10803_ _10764_ csr.io_mem_pc\[18\] VGND VGND VPWR VPWR _10869_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_153_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17614_ decode.regfile.registers_22\[20\] _13100_ _03020_ _13289_ VGND VGND VPWR
+ VPWR _03021_ sky130_fd_sc_hd__a211o_1
X_18594_ _03708_ decode.id_ex_imm_reg\[22\] _03891_ _03892_ VGND VGND VPWR VPWR _03893_
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_114_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14757_ csr.io_mem_pc\[19\] VGND VGND VPWR VPWR _10800_ sky130_fd_sc_hd__clkbuf_8
X_17545_ net469 _12872_ _13452_ _13491_ _13219_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_138_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13708_ _10057_ VGND VGND VPWR VPWR _10058_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17476_ decode.regfile.registers_2\[17\] _12834_ _12639_ decode.regfile.registers_3\[17\]
+ _12837_ VGND VGND VPWR VPWR _13424_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14688_ _10730_ VGND VGND VPWR VPWR _10731_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19215_ _04470_ _04510_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13639_ memory.csr_read_data_out_reg\[6\] _09989_ _09997_ VGND VGND VPWR VPWR _09998_
+ sky130_fd_sc_hd__o21ai_4
X_16427_ decode.regfile.registers_7\[29\] _11378_ _12393_ _12394_ _11134_ VGND VGND
+ VPWR VPWR _12395_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_171_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16358_ _11194_ decode.regfile.registers_12\[27\] decode.regfile.registers_13\[27\]
+ _11196_ _11198_ VGND VGND VPWR VPWR _12328_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19146_ _04442_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15309_ _11043_ decode.regfile.registers_4\[1\] _11190_ _10628_ _11083_ VGND VGND
+ VPWR VPWR _11305_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16289_ decode.regfile.registers_19\[25\] _11354_ _11218_ _12260_ VGND VGND VPWR
+ VPWR _12261_ sky130_fd_sc_hd__o211a_1
X_19077_ _04334_ _04117_ _04233_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18028_ _12595_ _03422_ _03423_ _12591_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_2_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19979_ net432 _05217_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22990_ _07112_ _07436_ _07082_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21941_ net2800 _06496_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__or2_1
XFILLER_0_222_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24660_ net1107 VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__clkbuf_1
X_21872_ _06496_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_132_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23611_ _07951_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20823_ _03582_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24591_ net1852 execute.io_target_pc\[17\] _08473_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26330_ _09385_ _09492_ VGND VGND VPWR VPWR _09500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_212_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23542_ net2210 _07904_ _07901_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__or3b_1
XFILLER_0_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20754_ csr.io_csr_address\[4\] _05214_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_214_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26261_ net597 _09447_ _09460_ _09458_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__o211a_1
X_23473_ _10662_ _07862_ _07873_ VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20685_ _03728_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__buf_2
X_28000_ clknet_leaf_204_clock _01022_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25212_ _08051_ net1574 _08041_ VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22424_ fetch.bht.bhtTable_tag\[0\]\[12\] fetch.bht.bhtTable_tag\[1\]\[12\] fetch.bht.bhtTable_tag\[2\]\[12\]
+ fetch.bht.bhtTable_tag\[3\]\[12\] _06644_ _06650_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__mux4_1
XFILLER_0_165_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26192_ _09412_ _09413_ VGND VGND VPWR VPWR _09414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25143_ net89 _06248_ _10916_ _07383_ _05856_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__o311a_2
X_22355_ _06949_ _06677_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21306_ net1327 _10812_ _06157_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25074_ _10019_ _08762_ _08763_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__and3_1
X_22286_ _06879_ _06880_ _06627_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24025_ net1470 execute.io_target_pc\[1\] _08014_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__mux2_1
X_28902_ clknet_leaf_97_clock _01915_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_21237_ _10872_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__buf_2
Xhold260 decode.regfile.registers_27\[30\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_208_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29882_ clknet_leaf_305_clock _02895_ VGND VGND VPWR VPWR decode.regfile.registers_20\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold271 decode.regfile.registers_30\[31\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_208_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold282 decode.regfile.registers_31\[25\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_1
XFILLER_0_218_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_208_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 decode.regfile.registers_19\[11\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
X_28833_ clknet_leaf_183_clock _01846_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_21168_ _06078_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20119_ _05327_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__and2_1
X_28764_ clknet_leaf_181_clock _01777_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21099_ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__clkbuf_4
X_13990_ _09999_ _10244_ VGND VGND VPWR VPWR _10253_ sky130_fd_sc_hd__nand2_1
X_25976_ _08973_ _09241_ VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_1007 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24927_ csr._mcycle_T_3\[43\] csr._mcycle_T_3\[42\] _08661_ VGND VGND VPWR VPWR _08665_
+ sky130_fd_sc_hd__and3_1
X_27715_ clknet_leaf_19_clock _00744_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_28695_ clknet_leaf_117_clock _01708_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15660_ _11059_ _10976_ _11048_ _11085_ VGND VGND VPWR VPWR _11648_ sky130_fd_sc_hd__or4_4
XFILLER_0_77_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_100 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24858_ _06136_ net2224 _08607_ VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__mux2_1
X_27646_ clknet_leaf_45_clock _00675_ VGND VGND VPWR VPWR execute.io_reg_pc\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_111 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ decode.immGen._imm_T_24\[2\] VGND VGND VPWR VPWR _10654_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23809_ execute.io_target_pc\[5\] VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__buf_2
XANTENNA_133 _10662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27577_ clknet_leaf_159_clock _00606_ VGND VGND VPWR VPWR csr.io_mem_pc\[18\] sky130_fd_sc_hd__dfxtp_4
X_15591_ decode.regfile.registers_2\[7\] _11129_ _11147_ _11151_ _11580_ VGND VGND
+ VPWR VPWR _11581_ sky130_fd_sc_hd__o311a_1
XANTENNA_144 execute.io_reg_pc\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24789_ _08083_ net1146 _08574_ VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _12500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17330_ decode.regfile.registers_15\[13\] _12555_ _10923_ _12876_ _13031_ VGND VGND
+ VPWR VPWR _13282_ sky130_fd_sc_hd__a41o_1
XFILLER_0_28_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29316_ clknet_leaf_225_clock _02329_ VGND VGND VPWR VPWR decode.regfile.registers_2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14542_ _10583_ _10584_ VGND VGND VPWR VPWR _10585_ sky130_fd_sc_hd__nand2_1
X_26528_ net2343 _09605_ _09613_ _09608_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17261_ _10928_ VGND VGND VPWR VPWR _13215_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_78_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29247_ clknet_leaf_233_clock _02260_ VGND VGND VPWR VPWR decode.regfile.registers_0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_26459_ net2428 _09561_ _09573_ _09567_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__o211a_1
X_14473_ net469 _10520_ _10531_ _10522_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19000_ decode.id_ex_aluop_reg\[0\] VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16212_ _11072_ _11205_ _12185_ VGND VGND VPWR VPWR _12186_ sky130_fd_sc_hd__a21oi_1
X_29178_ clknet_leaf_164_clock _02191_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17192_ _13142_ _13144_ _13146_ VGND VGND VPWR VPWR _13147_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28129_ clknet_leaf_217_clock _01151_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16143_ decode.regfile.registers_16\[21\] _11124_ _12101_ _12118_ VGND VGND VPWR
+ VPWR _12119_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_12_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16074_ _11403_ _12049_ _12050_ _12051_ VGND VGND VPWR VPWR _12052_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15025_ _11032_ _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__a31o_1
X_19902_ _05170_ _05115_ _04248_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19833_ _03811_ _05079_ _03829_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_87_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19764_ _04508_ _04301_ _04650_ _05033_ _05038_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__o311a_1
XFILLER_0_78_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16976_ decode.regfile.registers_1\[5\] _12932_ _12933_ _10615_ _12935_ VGND VGND
+ VPWR VPWR _12936_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_78_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18715_ _04010_ _03699_ net246 decode.id_ex_rs1_data_reg\[2\] _04013_ VGND VGND VPWR
+ VPWR _04014_ sky130_fd_sc_hd__o221a_2
Xinput6 net384 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
X_15927_ _11445_ _11907_ _11908_ VGND VGND VPWR VPWR _11909_ sky130_fd_sc_hd__o21a_1
XFILLER_0_223_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19695_ _04191_ _03956_ _03959_ _03947_ _03944_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__a32o_1
XFILLER_0_204_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18646_ _03797_ _03942_ _03889_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15858_ decode.regfile.registers_5\[14\] _10636_ _11138_ VGND VGND VPWR VPWR _11841_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_176_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14809_ _10786_ _10789_ _10793_ _10794_ _10851_ VGND VGND VPWR VPWR _10852_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_176_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18577_ decode.io_wb_rd\[2\] csr.io_csr_address\[2\] VGND VGND VPWR VPWR _03876_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_59_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15789_ decode.regfile.registers_8\[12\] _11046_ _11175_ VGND VGND VPWR VPWR _11774_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17528_ _12572_ _13473_ _13474_ VGND VGND VPWR VPWR _13475_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17459_ _13407_ decode.regfile.registers_25\[16\] _13045_ _13294_ VGND VGND VPWR
+ VPWR _13408_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20470_ _05611_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19129_ _04321_ _04234_ _04277_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22140_ fetch.bht.bhtTable_tag\[0\]\[4\] fetch.bht.bhtTable_tag\[1\]\[4\] net303
+ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22071_ fetch.bht.bhtTable_tag\[12\]\[18\] fetch.bht.bhtTable_tag\[13\]\[18\] _06619_
+ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21022_ _05995_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25830_ _09197_ VGND VGND VPWR VPWR _09198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25761_ net1344 _09156_ _09159_ _09153_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__o211a_1
X_22973_ _07419_ _07420_ _06633_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24712_ _08074_ net1732 _08531_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__mux2_1
X_27500_ clknet_leaf_30_clock _00529_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_195_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21924_ csr.io_mret_vector\[26\] _10760_ _06539_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__mux2_1
X_28480_ clknet_leaf_165_clock _01493_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25692_ _08916_ _09112_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_195_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27431_ clknet_leaf_49_clock _00460_ VGND VGND VPWR VPWR decode.id_ex_memread_reg
+ sky130_fd_sc_hd__dfxtp_4
X_24643_ _08504_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_182_Right_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21855_ _06507_ _06494_ _06495_ _06508_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27362_ clknet_leaf_33_clock _00391_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_20806_ net100 _05867_ _05875_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__and3_1
XFILLER_0_195_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24574_ net1084 execute.io_target_pc\[9\] _08462_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21786_ _06456_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29101_ clknet_leaf_17_clock _02114_ VGND VGND VPWR VPWR csr._mcycle_T_3\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26313_ _10373_ _10195_ _10240_ _08903_ VGND VGND VPWR VPWR _09489_ sky130_fd_sc_hd__and4_1
X_23525_ net2200 _07904_ _07901_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__or3b_1
XFILLER_0_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27293_ clknet_leaf_5_clock _00322_ VGND VGND VPWR VPWR decode.regfile.registers_31\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_20737_ _05804_ _03596_ _05839_ net183 net2656 VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29032_ clknet_leaf_99_clock _02045_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_154_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26244_ _09450_ _09448_ VGND VGND VPWR VPWR _09451_ sky130_fd_sc_hd__nand2_1
X_23456_ _04459_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20668_ _05576_ _05579_ _05584_ _03594_ decode.id_ex_funct3_reg\[1\] VGND VGND VPWR
+ VPWR _05795_ sky130_fd_sc_hd__o311a_1
XFILLER_0_18_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22407_ fetch.bht.bhtTable_tag\[6\]\[21\] fetch.bht.bhtTable_tag\[7\]\[21\] _06707_
+ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__mux2_1
X_26175_ _10047_ VGND VGND VPWR VPWR _09402_ sky130_fd_sc_hd__buf_4
X_23387_ _07807_ _07810_ _07084_ VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20599_ _05541_ csr.io_mret_vector\[22\] _05602_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_167_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25126_ _08791_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__clkbuf_1
X_22338_ fetch.bht.bhtTable_tag\[2\]\[10\] fetch.bht.bhtTable_tag\[3\]\[10\] _06644_
+ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25057_ csr._mcycle_T_2\[23\] _08704_ _08750_ _08751_ VGND VGND VPWR VPWR _08752_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_163_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29934_ clknet_leaf_341_clock _02947_ VGND VGND VPWR VPWR decode.regfile.registers_21\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_22269_ _06834_ _06849_ _06863_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_163_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24008_ _08175_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29865_ clknet_leaf_302_clock _02878_ VGND VGND VPWR VPWR decode.regfile.registers_19\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28816_ clknet_leaf_121_clock _01829_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_16830_ decode.regfile.registers_10\[2\] _12790_ _12792_ VGND VGND VPWR VPWR _12793_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_228_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29796_ clknet_leaf_292_clock _02809_ VGND VGND VPWR VPWR decode.regfile.registers_17\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28747_ clknet_leaf_95_clock _01760_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13973_ _10241_ VGND VGND VPWR VPWR _10242_ sky130_fd_sc_hd__clkbuf_4
X_16761_ _11016_ _10608_ _12508_ _12502_ VGND VGND VPWR VPWR _12725_ sky130_fd_sc_hd__or4_4
XFILLER_0_219_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25959_ _08956_ _09267_ VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_122_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18500_ _03759_ _03793_ decode.id_ex_rs2_data_reg\[28\] _03747_ _03728_ VGND VGND
+ VPWR VPWR _03799_ sky130_fd_sc_hd__o221a_1
X_15712_ _11698_ decode.regfile.registers_5\[10\] _11291_ VGND VGND VPWR VPWR _11699_
+ sky130_fd_sc_hd__mux2_1
X_16692_ _12497_ _10606_ _10935_ _12510_ VGND VGND VPWR VPWR _12657_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19480_ _04504_ _04225_ net271 _04465_ _04765_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__o311a_1
X_28678_ clknet_leaf_95_clock _01691_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_87_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18431_ decode.io_wb_rd\[4\] csr.io_csr_address\[4\] VGND VGND VPWR VPWR _03730_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_200_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27629_ clknet_leaf_154_clock _00658_ VGND VGND VPWR VPWR execute.io_reg_pc\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_15643_ _11094_ _11114_ _11119_ _11203_ decode.regfile.registers_16\[8\] VGND VGND
+ VPWR VPWR _11632_ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_1210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15574_ _11436_ decode.regfile.registers_26\[6\] _11349_ _10980_ _11564_ VGND VGND
+ VPWR VPWR _11565_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_83_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ execute.io_mem_memtoreg\[0\] VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14525_ _10569_ _09881_ _09884_ VGND VGND VPWR VPWR _10570_ sky130_fd_sc_hd__or3b_2
X_17313_ decode.regfile.registers_17\[13\] _11022_ _12567_ _12586_ VGND VGND VPWR
+ VPWR _13265_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18293_ _03611_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14456_ net514 _10520_ _10521_ _10522_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__o211a_1
X_17244_ decode.regfile.registers_8\[11\] _12889_ _12606_ _13197_ VGND VGND VPWR VPWR
+ _13198_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17175_ _12915_ decode.regfile.registers_25\[9\] _13045_ _12812_ VGND VGND VPWR VPWR
+ _13131_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_42_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14387_ net430 _10477_ _10482_ _10481_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16126_ decode.regfile.registers_11\[21\] _11071_ _11204_ _11407_ VGND VGND VPWR
+ VPWR _12102_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16057_ decode.regfile.registers_12\[19\] _11047_ _11690_ VGND VGND VPWR VPWR _12035_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_55_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15008_ _11017_ VGND VGND VPWR VPWR _11018_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2408 fetch.btb.btbTable\[13\]\[1\] VGND VGND VPWR VPWR net2635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2419 _01287_ VGND VGND VPWR VPWR net2646 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19816_ _04949_ _05085_ _05086_ _05088_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__o31a_1
Xhold1707 fetch.bht.bhtTable_target_pc\[6\]\[13\] VGND VGND VPWR VPWR net1934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1718 decode.regfile.registers_12\[15\] VGND VGND VPWR VPWR net1945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1729 execute.csr_write_data_out_reg\[29\] VGND VGND VPWR VPWR net1956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19747_ _03924_ _03937_ _03903_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_194_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16959_ _12701_ decode.regfile.registers_28\[4\] _12698_ VGND VGND VPWR VPWR _12920_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_205_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19678_ _04191_ _03960_ _04938_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__nand3_1
XFILLER_0_79_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18629_ _03817_ _03927_ _03774_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_177_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21640_ net2749 _06338_ _06355_ _06356_ _06336_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__a311oi_1
XTAP_TAPCELL_ROW_190_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21571_ _06282_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_16_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 _01447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_22 _05857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23310_ execute.io_target_pc\[24\] _07090_ _06041_ _06037_ VGND VGND VPWR VPWR _07739_
+ sky130_fd_sc_hd__a211o_1
X_20522_ _03588_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_33 _10019_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24290_ _08320_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_44 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 _10604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_66 _11027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23241_ _07619_ _07573_ _07620_ _07674_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__a31o_1
XANTENNA_77 _11143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20453_ csr.msip _05539_ _05522_ _05606_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__o32a_1
XANTENNA_88 decode.id_ex_rs1_data_reg\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23172_ _07606_ _07112_ _07076_ _07608_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20384_ net2802 _05531_ _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22123_ net98 VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__buf_4
XFILLER_0_112_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27980_ clknet_leaf_198_clock _01002_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput140 net140 VGND VGND VPWR VPWR io_memory_write_data[13] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput151 net151 VGND VGND VPWR VPWR io_memory_write_data[23] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput162 net162 VGND VGND VPWR VPWR io_memory_write_data[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22054_ _00001_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__buf_4
X_26931_ _09992_ _09840_ VGND VGND VPWR VPWR _09846_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_2 _00551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21005_ _05986_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__clkbuf_1
X_29650_ clknet_leaf_280_clock _02663_ VGND VGND VPWR VPWR decode.regfile.registers_12\[24\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_197_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26862_ _09794_ VGND VGND VPWR VPWR _09806_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_197_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28601_ clknet_leaf_127_clock _01614_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25813_ net2466 _09183_ _09188_ _09182_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26793_ _09396_ _09763_ VGND VGND VPWR VPWR _09767_ sky130_fd_sc_hd__nand2_1
X_29581_ clknet_leaf_273_clock _02594_ VGND VGND VPWR VPWR decode.regfile.registers_10\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_28532_ clknet_leaf_237_clock _01545_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25744_ net2452 _09139_ _09148_ _09142_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__o211a_1
X_22956_ _07076_ _07404_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21907_ net2754 _06545_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28463_ clknet_leaf_138_clock _01476_ VGND VGND VPWR VPWR decode.io_id_pc\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25675_ _08975_ _09067_ VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22887_ _07340_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24626_ _08495_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_156_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27414_ clknet_leaf_10_clock _00443_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[23\]
+ sky130_fd_sc_hd__dfxtp_4
X_28394_ clknet_leaf_142_clock _01407_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_2
X_21838_ _06496_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27345_ clknet_leaf_44_clock _00374_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[18\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_14_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24557_ net1117 execute.io_target_pc\[1\] _07335_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21769_ _06447_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14310_ _10048_ _10431_ VGND VGND VPWR VPWR _10438_ sky130_fd_sc_hd__nand2_1
X_23508_ net2195 _07890_ _07887_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27276_ clknet_leaf_11_clock _00305_ VGND VGND VPWR VPWR decode.regfile.registers_30\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15290_ _11129_ _10627_ _11042_ _11069_ VGND VGND VPWR VPWR _11286_ sky130_fd_sc_hd__or4b_1
X_24488_ _08424_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__clkbuf_1
Xwire212 net350 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29015_ clknet_leaf_125_clock _02028_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_26227_ _10135_ VGND VGND VPWR VPWR _09438_ sky130_fd_sc_hd__buf_4
XFILLER_0_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14241_ _10290_ VGND VGND VPWR VPWR _10398_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23439_ net31 _07846_ _07854_ _07851_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_115_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14172_ _10081_ _10355_ VGND VGND VPWR VPWR _10358_ sky130_fd_sc_hd__nand2_1
X_26158_ _09372_ VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_186_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25109_ _06126_ net1902 _08778_ VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26089_ _08935_ _09340_ VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18980_ decode.id_ex_rs2_data_reg\[2\] net199 _04010_ _04046_ _04015_ VGND VGND VPWR
+ VPWR _04279_ sky130_fd_sc_hd__o221a_4
X_17931_ _10928_ decode.regfile.registers_26\[28\] _12814_ _11011_ _11027_ VGND VGND
+ VPWR VPWR _03330_ sky130_fd_sc_hd__o2111a_1
X_29917_ clknet_leaf_335_clock _02930_ VGND VGND VPWR VPWR decode.regfile.registers_21\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29848_ clknet_leaf_307_clock _02861_ VGND VGND VPWR VPWR decode.regfile.registers_18\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17862_ net463 _12872_ _03225_ _03262_ _03073_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19601_ _04442_ _04294_ _04362_ _04806_ _04728_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__o311a_4
XFILLER_0_219_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16813_ _10593_ VGND VGND VPWR VPWR _12776_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_145_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29779_ clknet_leaf_294_clock _02792_ VGND VGND VPWR VPWR decode.regfile.registers_16\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_17793_ decode.regfile.registers_6\[25\] _10603_ _12615_ _12623_ _03194_ VGND VGND
+ VPWR VPWR _03195_ sky130_fd_sc_hd__o32a_1
XFILLER_0_191_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19532_ _04281_ _04283_ _04814_ _04815_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_85_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16744_ _12707_ VGND VGND VPWR VPWR _12708_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_220_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13956_ net2566 _10226_ _10231_ _10232_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19463_ _04112_ _04118_ _04425_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__a31o_2
X_16675_ decode.regfile.registers_2\[0\] _10608_ _12636_ _12639_ VGND VGND VPWR VPWR
+ _12640_ sky130_fd_sc_hd__a31o_1
X_13887_ _10136_ _10152_ VGND VGND VPWR VPWR _10191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_201 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_212 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18414_ _03640_ csr.io_csr_address\[3\] VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15626_ decode.regfile.registers_0\[8\] _11154_ _11503_ _11148_ VGND VGND VPWR VPWR
+ _11615_ sky130_fd_sc_hd__o2bb2ai_1
XINSDIODE1_223 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_234 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19394_ _04664_ _04142_ _04177_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_245 net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_256 clknet_0_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_267 _06691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18345_ _09921_ _03641_ _03643_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_278 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ decode.regfile.registers_8\[6\] _11166_ _11547_ decode.regfile.registers_9\[6\]
+ _11183_ VGND VGND VPWR VPWR _11548_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_84_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_289 _12504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14508_ _09879_ _10552_ _09882_ VGND VGND VPWR VPWR _10553_ sky130_fd_sc_hd__and3b_1
Xclkbuf_leaf_334_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_334_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15488_ decode.regfile.registers_21\[4\] _11062_ _11100_ _11229_ _11480_ VGND VGND
+ VPWR VPWR _11481_ sky130_fd_sc_hd__o311a_1
X_18276_ _03602_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput20 net377 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17227_ _13055_ net2791 _13097_ VGND VGND VPWR VPWR _13181_ sky130_fd_sc_hd__o21a_1
Xinput31 net530 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
X_14439_ net918 _10506_ _10512_ _10509_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 io_memory_read_data[17] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_163_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput53 io_memory_read_data[27] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput64 io_memory_read_data[8] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_1
Xhold804 fetch.bht.bhtTable_target_pc\[3\]\[21\] VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__dlygate4sd3_1
X_17158_ _12654_ _13111_ _13112_ _13113_ VGND VGND VPWR VPWR _13114_ sky130_fd_sc_hd__a31o_1
XFILLER_0_204_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold815 decode.regfile.registers_25\[10\] VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 fetch.bht.bhtTable_tag\[1\]\[1\] VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold837 csr.minstret\[0\] VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold848 fetch.bht.bhtTable_tag\[15\]\[22\] VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ _10958_ decode.regfile.registers_24\[20\] _11074_ VGND VGND VPWR VPWR _12086_
+ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_349_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_349_clock
+ sky130_fd_sc_hd__clkbuf_8
X_17089_ _11010_ VGND VGND VPWR VPWR _13047_ sky130_fd_sc_hd__clkbuf_4
Xhold859 decode.regfile.registers_17\[8\] VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2205 decode.regfile.registers_5\[22\] VGND VGND VPWR VPWR net2432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2216 decode.regfile.registers_23\[22\] VGND VGND VPWR VPWR net2443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2227 decode.regfile.registers_4\[26\] VGND VGND VPWR VPWR net2454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2238 decode.regfile.registers_17\[24\] VGND VGND VPWR VPWR net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 fetch.bht.bhtTable_tag\[13\]\[18\] VGND VGND VPWR VPWR net2476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1504 decode.regfile.registers_19\[1\] VGND VGND VPWR VPWR net1731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1515 fetch.bht.bhtTable_target_pc\[7\]\[31\] VGND VGND VPWR VPWR net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 fetch.bht.bhtTable_tag\[2\]\[12\] VGND VGND VPWR VPWR net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1537 csr._minstret_T_3\[57\] VGND VGND VPWR VPWR net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1548 fetch.bht.bhtTable_target_pc\[2\]\[10\] VGND VGND VPWR VPWR net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 fetch.bht.bhtTable_tag\[9\]\[1\] VGND VGND VPWR VPWR net1786 sky130_fd_sc_hd__dlygate4sd3_1
X_22810_ _07300_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23790_ _08047_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22741_ _06115_ net1364 _09903_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25460_ _08912_ _08980_ VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22672_ _07209_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_220_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24411_ net1080 execute.io_target_pc\[28\] _09911_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__mux2_1
X_21623_ _06343_ _06344_ _06317_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25391_ _10052_ VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__buf_6
XFILLER_0_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27130_ clknet_leaf_357_clock _00159_ VGND VGND VPWR VPWR decode.regfile.registers_26\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24342_ _08347_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_151_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21554_ _06297_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20505_ csr._csr_read_data_T_8\[9\] _05622_ _05651_ _05653_ _05655_ VGND VGND VPWR
+ VPWR _05656_ sky130_fd_sc_hd__a221o_2
XFILLER_0_132_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27061_ clknet_leaf_331_clock _00090_ VGND VGND VPWR VPWR decode.regfile.registers_24\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24273_ _08101_ net1391 _06218_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__mux2_1
X_21485_ _06259_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26012_ net2297 _09300_ _09303_ _09292_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23224_ fetch.bht.bhtTable_target_pc\[12\]\[19\] fetch.bht.bhtTable_target_pc\[13\]\[19\]
+ _07119_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20436_ _05559_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23155_ fetch.bht.bhtTable_target_pc\[0\]\[15\] fetch.bht.bhtTable_target_pc\[1\]\[15\]
+ fetch.bht.bhtTable_target_pc\[2\]\[15\] fetch.bht.bhtTable_target_pc\[3\]\[15\]
+ _07107_ _07114_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__mux4_1
X_20367_ csr.io_csr_address\[11\] _05523_ _05520_ _05524_ _05529_ VGND VGND VPWR VPWR
+ _05530_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_149_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22106_ fetch.bht.bhtTable_tag\[2\]\[3\] fetch.bht.bhtTable_tag\[3\]\[3\] _06700_
+ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23086_ _07076_ _07527_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__nand2_1
X_27963_ clknet_leaf_218_clock _00985_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_224_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20298_ _05418_ _05338_ _05473_ _05474_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_41_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_224_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29702_ clknet_leaf_286_clock _02715_ VGND VGND VPWR VPWR decode.regfile.registers_14\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22037_ _06631_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26914_ _09443_ _09794_ VGND VGND VPWR VPWR _09835_ sky130_fd_sc_hd__nand2_1
X_27894_ clknet_leaf_18_clock _00923_ VGND VGND VPWR VPWR csr._mcycle_T_2\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_76_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29633_ clknet_leaf_287_clock _02646_ VGND VGND VPWR VPWR decode.regfile.registers_12\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26845_ _10245_ _09796_ VGND VGND VPWR VPWR _09797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13810_ memory.io_wb_reg_pc\[31\] _10001_ VGND VGND VPWR VPWR _10144_ sky130_fd_sc_hd__and2_1
X_14790_ decode.id_ex_pc_reg\[1\] csr.io_mem_pc\[1\] VGND VGND VPWR VPWR _10833_ sky130_fd_sc_hd__and2_1
X_29564_ clknet_leaf_251_clock _02577_ VGND VGND VPWR VPWR decode.regfile.registers_10\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_23988_ _08165_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26776_ _09379_ _09753_ VGND VGND VPWR VPWR _09757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28515_ clknet_leaf_193_clock _01528_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13741_ memory.csr_read_data_out_reg\[20\] _10010_ _10085_ VGND VGND VPWR VPWR _10086_
+ sky130_fd_sc_hd__o21ai_4
X_22939_ fetch.bht.bhtTable_target_pc\[0\]\[3\] fetch.bht.bhtTable_target_pc\[1\]\[3\]
+ fetch.bht.bhtTable_target_pc\[2\]\[3\] fetch.bht.bhtTable_target_pc\[3\]\[3\] _07384_
+ _07113_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__mux4_1
X_25727_ _09110_ VGND VGND VPWR VPWR _09139_ sky130_fd_sc_hd__clkbuf_4
X_29495_ clknet_leaf_264_clock _02508_ VGND VGND VPWR VPWR decode.regfile.registers_7\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28446_ clknet_leaf_145_clock _01459_ VGND VGND VPWR VPWR decode.io_id_pc\[4\] sky130_fd_sc_hd__dfxtp_1
X_16460_ _12422_ _12425_ _12426_ VGND VGND VPWR VPWR _12427_ sky130_fd_sc_hd__o21ai_1
X_13672_ _09937_ VGND VGND VPWR VPWR _10027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_211_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25658_ _08958_ _09092_ VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_175_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15411_ _10957_ decode.regfile.registers_22\[3\] _11404_ _10978_ _10990_ VGND VGND
+ VPWR VPWR _11405_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_66_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24609_ net950 execute.io_target_pc\[26\] _09897_ VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16391_ decode.regfile.registers_8\[28\] _11285_ _11365_ decode.regfile.registers_9\[28\]
+ _11381_ VGND VGND VPWR VPWR _12360_ sky130_fd_sc_hd__o221a_1
X_28377_ clknet_leaf_192_clock _01390_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25589_ net2349 _09052_ _09058_ _09059_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18130_ _10909_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__clkbuf_2
X_15342_ _10978_ VGND VGND VPWR VPWR _11338_ sky130_fd_sc_hd__clkbuf_4
X_27328_ clknet_leaf_41_clock _00357_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18061_ _10910_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__buf_2
X_15273_ _11268_ VGND VGND VPWR VPWR _11269_ sky130_fd_sc_hd__buf_2
XFILLER_0_151_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27259_ clknet_leaf_5_clock _00288_ VGND VGND VPWR VPWR decode.regfile.registers_30\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17012_ decode.regfile.registers_1\[6\] _12778_ _12830_ _12970_ VGND VGND VPWR VPWR
+ _12971_ sky130_fd_sc_hd__o211ai_2
X_14224_ net706 _10376_ _10388_ _10385_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14155_ net660 _10346_ _10348_ _10344_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14086_ net2532 _10302_ _10308_ _10304_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__o211a_1
X_18963_ _03990_ _03991_ _03996_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17914_ decode.regfile.registers_7\[28\] _10615_ _13020_ _12621_ decode.regfile.registers_6\[28\]
+ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18894_ _04191_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_219_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17845_ decode.regfile.registers_15\[26\] _12585_ _03244_ _03245_ VGND VGND VPWR
+ VPWR _03246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_201_Left_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17776_ _02986_ decode.regfile.registers_26\[24\] _13002_ _13484_ _02987_ VGND VGND
+ VPWR VPWR _03179_ sky130_fd_sc_hd__o2111a_1
X_14988_ decode.control.io_opcode\[3\] _10583_ _10584_ _10968_ VGND VGND VPWR VPWR
+ _11005_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19515_ _04514_ _04798_ _04633_ _04799_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_18_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16727_ _12521_ _12689_ _12691_ VGND VGND VPWR VPWR _12692_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13939_ net2104 _10213_ _10222_ _10219_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19446_ _04112_ _04149_ _04234_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16658_ _12622_ VGND VGND VPWR VPWR _12623_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_102_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15609_ decode.regfile.registers_20\[7\] _11103_ _11222_ _11598_ VGND VGND VPWR VPWR
+ _11599_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_273_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_273_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19377_ _04311_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16589_ _12523_ VGND VGND VPWR VPWR _12554_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18328_ decode.id_ex_rs2_data_reg\[29\] _03627_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_210_Left_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18259_ csr.io_trapped csr.io_mret VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__nor2_4
XFILLER_0_114_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_288_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_288_clock
+ sky130_fd_sc_hd__clkbuf_8
X_21270_ _06139_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold601 fetch.bht.bhtTable_target_pc\[11\]\[15\] VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold612 fetch.bht.bhtTable_target_pc\[1\]\[31\] VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold623 fetch.bht.bhtTable_target_pc\[4\]\[28\] VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__dlygate4sd3_1
X_20221_ decode.id_ex_rdsel_reg VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__inv_2
Xhold634 fetch.bht.bhtTable_tag\[2\]\[25\] VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold645 decode.regfile.registers_11\[31\] VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 fetch.bht.bhtTable_target_pc\[8\]\[19\] VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold667 decode.regfile.registers_19\[13\] VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_2_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20152_ decode.id_ex_imm_reg\[22\] _10864_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold678 decode.regfile.registers_21\[31\] VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 fetch.bht.bhtTable_tag\[9\]\[17\] VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_211_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_211_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2002 execute.csr_write_data_out_reg\[14\] VGND VGND VPWR VPWR net2229 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2013 decode.regfile.registers_8\[17\] VGND VGND VPWR VPWR net2240 sky130_fd_sc_hd__dlygate4sd3_1
X_24960_ net2354 _08685_ _08686_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__o21ba_1
Xhold2024 fetch.bht.bhtTable_tag\[2\]\[21\] VGND VGND VPWR VPWR net2251 sky130_fd_sc_hd__dlygate4sd3_1
X_20083_ decode.id_ex_imm_reg\[11\] decode.id_ex_pc_reg\[11\] VGND VGND VPWR VPWR
+ _05298_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2035 fetch.bht.bhtTable_tag\[5\]\[11\] VGND VGND VPWR VPWR net2262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1301 decode.regfile.registers_28\[19\] VGND VGND VPWR VPWR net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2046 decode.regfile.registers_28\[22\] VGND VGND VPWR VPWR net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23911_ _08125_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__clkbuf_1
Xhold1312 fetch.bht.bhtTable_tag\[14\]\[1\] VGND VGND VPWR VPWR net1539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2057 decode.regfile.registers_8\[22\] VGND VGND VPWR VPWR net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 fetch.bht.bhtTable_tag\[13\]\[0\] VGND VGND VPWR VPWR net1550 sky130_fd_sc_hd__dlygate4sd3_1
X_24891_ _03555_ csr.mcycle\[23\] csr.mcycle\[26\] csr.mcycle\[25\] VGND VGND VPWR
+ VPWR _08640_ sky130_fd_sc_hd__and4_1
Xhold2068 decode.regfile.registers_18\[3\] VGND VGND VPWR VPWR net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2079 csr._csr_read_data_T_8\[8\] VGND VGND VPWR VPWR net2306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 execute.csr_write_data_out_reg\[9\] VGND VGND VPWR VPWR net1561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 decode.regfile.registers_22\[5\] VGND VGND VPWR VPWR net1572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23842_ _08082_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1356 fetch.bht.bhtTable_tag\[9\]\[5\] VGND VGND VPWR VPWR net1583 sky130_fd_sc_hd__dlygate4sd3_1
X_26630_ net888 _09665_ _09672_ _09660_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1367 fetch.bht.bhtTable_tag\[6\]\[10\] VGND VGND VPWR VPWR net1594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_226_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_226_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1378 fetch.bht.bhtTable_tag\[10\]\[9\] VGND VGND VPWR VPWR net1605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1389 fetch.bht.bhtTable_target_pc\[5\]\[5\] VGND VGND VPWR VPWR net1616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23773_ _08038_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__clkbuf_1
X_26561_ _09389_ _09632_ VGND VGND VPWR VPWR _09633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20985_ _05975_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28300_ clknet_leaf_164_clock _00012_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25512_ net2507 _09008_ _09014_ _09004_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__o211a_1
X_22724_ _10941_ _03458_ _03541_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__and3_1
X_29280_ clknet_leaf_243_clock _02293_ VGND VGND VPWR VPWR decode.regfile.registers_1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_26492_ net1197 _09592_ _09593_ _09582_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28231_ clknet_leaf_55_clock _01253_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfxtp_2
X_25443_ _10141_ VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_217_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22655_ net2654 _07208_ _07213_ _07164_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21606_ csr.minstret\[0\] csr.minstret\[1\] csr.minstret\[2\] csr.minstret\[3\] VGND
+ VGND VPWR VPWR _06332_ sky130_fd_sc_hd__and4_1
XFILLER_0_165_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28162_ clknet_leaf_67_clock net560 VGND VGND VPWR VPWR csr._csr_read_data_T_9\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_25374_ _10024_ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__buf_4
X_22586_ net2501 _07166_ _07167_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24325_ _08087_ net1383 _08334_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27113_ clknet_leaf_348_clock _00142_ VGND VGND VPWR VPWR decode.regfile.registers_25\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28093_ clknet_leaf_168_clock _01115_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_21537_ _06288_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__clkbuf_1
Xclone45 net354 net228 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__nand2_2
XFILLER_0_133_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27044_ clknet_leaf_345_clock _00073_ VGND VGND VPWR VPWR decode.regfile.registers_23\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_24256_ _08303_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__clkbuf_1
X_21468_ net27 _10972_ _06249_ _10546_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_226_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_226_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23207_ _07110_ _07641_ _07080_ VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20419_ _05555_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24187_ _08081_ net1095 _08266_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21399_ _06147_ net1972 _06210_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23138_ fetch.bht.bhtTable_target_pc\[8\]\[14\] fetch.bht.bhtTable_target_pc\[9\]\[14\]
+ fetch.bht.bhtTable_target_pc\[10\]\[14\] fetch.bht.bhtTable_target_pc\[11\]\[14\]
+ _07123_ _07111_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__mux4_1
X_28995_ clknet_leaf_130_clock _02008_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23069_ _07439_ fetch.bht.bhtTable_target_pc\[14\]\[10\] _07125_ _07511_ VGND VGND
+ VPWR VPWR _07512_ sky130_fd_sc_hd__o211a_1
X_27946_ clknet_leaf_202_clock _00968_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_15960_ _11445_ _11939_ _11940_ _11246_ VGND VGND VPWR VPWR _11941_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14911_ _10942_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__clkbuf_1
X_27877_ clknet_leaf_65_clock _00906_ VGND VGND VPWR VPWR csr.io_ecause\[0\] sky130_fd_sc_hd__dfxtp_1
X_15891_ _11646_ _11834_ _11064_ decode.regfile.registers_29\[14\] _11873_ VGND VGND
+ VPWR VPWR _11874_ sky130_fd_sc_hd__o221a_1
XFILLER_0_216_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ decode.regfile.registers_1\[21\] _12636_ _13145_ _03035_ VGND VGND VPWR VPWR
+ _03036_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_106_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29616_ clknet_leaf_280_clock _02629_ VGND VGND VPWR VPWR decode.regfile.registers_11\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14842_ _10820_ _10821_ _10815_ csr.io_mem_pc\[8\] VGND VGND VPWR VPWR _10885_ sky130_fd_sc_hd__a31o_1
X_26828_ net2634 _09779_ _09786_ _09784_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1890 decode.regfile.registers_17\[0\] VGND VGND VPWR VPWR net2117 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_177_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17561_ decode.regfile.registers_11\[19\] _12595_ _12588_ _12551_ _02968_ VGND VGND
+ VPWR VPWR _02969_ sky130_fd_sc_hd__a221o_1
X_29547_ clknet_leaf_266_clock _02560_ VGND VGND VPWR VPWR decode.regfile.registers_9\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14773_ csr.io_mem_pc\[6\] csr.io_mem_pc\[7\] _10815_ VGND VGND VPWR VPWR _10816_
+ sky130_fd_sc_hd__and3_1
X_26759_ net2095 _09736_ _09746_ _09743_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19300_ _04279_ _04019_ _04427_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16512_ decode.regfile.registers_23\[31\] _11262_ _12453_ _12477_ _11335_ VGND VGND
+ VPWR VPWR _12478_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_67_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13724_ _10005_ _10001_ memory.io_wb_reg_pc\[18\] VGND VGND VPWR VPWR _10071_ sky130_fd_sc_hd__o21ai_1
X_17492_ decode.regfile.registers_21\[17\] _12716_ _13417_ _13439_ _12909_ VGND VGND
+ VPWR VPWR _13440_ sky130_fd_sc_hd__o221a_1
X_29478_ clknet_leaf_263_clock _02491_ VGND VGND VPWR VPWR decode.regfile.registers_7\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19231_ _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16443_ decode.regfile.registers_25\[29\] _11483_ _11484_ decode.regfile.registers_24\[29\]
+ VGND VGND VPWR VPWR _12411_ sky130_fd_sc_hd__o22a_1
X_28429_ clknet_leaf_247_clock _01442_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[19\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_112_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13655_ _09943_ VGND VGND VPWR VPWR _10012_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19162_ _03594_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16374_ _11396_ _12341_ _12342_ _12343_ VGND VGND VPWR VPWR _12344_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13586_ _09937_ VGND VGND VPWR VPWR _09951_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_136_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18113_ _03482_ _03480_ _03474_ net1955 VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__and4bb_1
X_15325_ _10651_ _11111_ _11118_ _11202_ decode.regfile.registers_16\[1\] VGND VGND
+ VPWR VPWR _11321_ sky130_fd_sc_hd__a32o_1
XFILLER_0_164_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19093_ decode.id_ex_aluop_reg\[1\] decode.id_ex_aluop_reg\[3\] decode.id_ex_aluop_reg\[2\]
+ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_42_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18044_ _10938_ decode.regfile.registers_25\[31\] _12505_ _12811_ VGND VGND VPWR
+ VPWR _03440_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15256_ _11062_ _11066_ _11054_ VGND VGND VPWR VPWR _11252_ sky130_fd_sc_hd__or3_2
XFILLER_0_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14207_ _09964_ _10377_ VGND VGND VPWR VPWR _10379_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15187_ _11183_ VGND VGND VPWR VPWR _11184_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14138_ net542 _10332_ _10338_ _10328_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__o211a_1
X_19995_ decode.id_ex_pcsel_reg VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18946_ _04244_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__clkbuf_4
X_14069_ net744 _10287_ _10298_ _10291_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18877_ _04166_ _04164_ _04154_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17828_ decode.regfile.registers_11\[26\] _12724_ _12587_ _12551_ VGND VGND VPWR
+ VPWR _03229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17759_ _03160_ _12603_ _12600_ _03161_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20770_ _03452_ _05425_ decode.csr_write_reg VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__and3b_1
XFILLER_0_193_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19429_ _04715_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22440_ net76 _07034_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22371_ fetch.bht.bhtTable_tag\[0\]\[16\] fetch.bht.bhtTable_tag\[1\]\[16\] fetch.bht.bhtTable_tag\[2\]\[16\]
+ fetch.bht.bhtTable_tag\[3\]\[16\] _06878_ _06621_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_212_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24110_ net1249 execute.io_target_pc\[10\] _08221_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21322_ _06171_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__clkbuf_1
X_25090_ _06107_ net2054 _08596_ VGND VGND VPWR VPWR _08773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24041_ _08192_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21253_ _10800_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__buf_2
Xhold420 decode.regfile.registers_23\[12\] VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold431 io_fetch_data[5] VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_150_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_150_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold442 decode.regfile.registers_16\[12\] VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20204_ _05385_ _05392_ _05395_ _05393_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_25_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold453 decode.regfile.registers_12\[27\] VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold464 decode.regfile.registers_8\[10\] VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__dlygate4sd3_1
X_21184_ _06087_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__clkbuf_1
Xhold475 decode.regfile.registers_22\[29\] VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 csr._minstret_T_3\[37\] VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap194 _10135_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_221_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold497 _01243_ VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27800_ clknet_leaf_317_clock _00829_ VGND VGND VPWR VPWR memory.io_wb_readdata\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20135_ _05332_ _05337_ _05333_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__o21ai_1
X_28780_ clknet_leaf_87_clock _01793_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_25992_ net2555 _09286_ _09291_ _09292_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27731_ clknet_leaf_70_clock _00760_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_165_clock clknet_5_25__leaf_clock VGND VGND VPWR VPWR clknet_leaf_165_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20066_ decode.id_ex_imm_reg\[10\] decode.id_ex_pc_reg\[10\] VGND VGND VPWR VPWR
+ _05283_ sky130_fd_sc_hd__nand2_1
X_24943_ net759 _08674_ _08675_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__o21ba_1
Xhold1120 fetch.bht.bhtTable_tag\[4\]\[22\] VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1131 fetch.bht.bhtTable_tag\[6\]\[1\] VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 fetch.bht.bhtTable_target_pc\[10\]\[19\] VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 _08233_ VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__dlygate4sd3_1
X_27662_ clknet_leaf_46_clock _00691_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_24874_ _06153_ net1504 _08388_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__mux2_1
Xhold1164 fetch.bht.bhtTable_target_pc\[6\]\[25\] VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 fetch.bht.bhtTable_tag\[3\]\[23\] VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_116_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29401_ clknet_leaf_247_clock _02414_ VGND VGND VPWR VPWR decode.regfile.registers_4\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1186 fetch.bht.bhtTable_tag\[11\]\[4\] VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__dlygate4sd3_1
X_26613_ _09443_ _09621_ VGND VGND VPWR VPWR _09662_ sky130_fd_sc_hd__nand2_1
XFILLER_0_224_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23825_ _08070_ net1091 _08058_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__mux2_1
Xhold1197 fetch.bht.bhtTable_target_pc\[9\]\[19\] VGND VGND VPWR VPWR net1424 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_219_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27593_ clknet_leaf_146_clock _00622_ VGND VGND VPWR VPWR execute.io_target_pc\[2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_135_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_219_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29332_ clknet_leaf_225_clock _02345_ VGND VGND VPWR VPWR decode.regfile.registers_2\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_23756_ _08029_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26544_ _10245_ _09623_ VGND VGND VPWR VPWR _09624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20968_ _05966_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_172_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22707_ net2575 _07235_ _07242_ _07234_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_172_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29263_ clknet_leaf_224_clock _02276_ VGND VGND VPWR VPWR decode.regfile.registers_0\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23687_ net821 _10821_ _07992_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__mux2_1
X_26475_ _09379_ _09579_ VGND VGND VPWR VPWR _09584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20899_ _05925_ _05921_ net35 VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28214_ clknet_leaf_84_clock net1610 VGND VGND VPWR VPWR csr.mscratch\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22638_ _07199_ _07200_ _07202_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__nor3_1
X_25426_ net507 _08951_ _08961_ _08950_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_103_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_103_clock
+ sky130_fd_sc_hd__clkbuf_8
X_29194_ clknet_leaf_245_clock _02207_ VGND VGND VPWR VPWR fetch.btb.btbTable\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28145_ clknet_leaf_200_clock _01167_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_25357_ net690 _08906_ _08913_ _07247_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__o211a_1
X_22569_ csr._minstret_T_3\[40\] _07153_ _06336_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15110_ decode.immGen._imm_T_24\[3\] decode.immGen._imm_T_24\[2\] VGND VGND VPWR
+ VPWR _11107_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_75_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24308_ _08070_ net1579 _08323_ VGND VGND VPWR VPWR _08330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16090_ decode.regfile.registers_6\[20\] _11170_ _12064_ _12066_ VGND VGND VPWR VPWR
+ _12067_ sky130_fd_sc_hd__a22oi_1
X_28076_ clknet_leaf_221_clock _01098_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25288_ _08874_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_131_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15041_ _11037_ VGND VGND VPWR VPWR _11038_ sky130_fd_sc_hd__clkbuf_4
X_24239_ _08294_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__clkbuf_1
X_27027_ clknet_leaf_331_clock _00056_ VGND VGND VPWR VPWR decode.regfile.registers_23\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_118_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_118_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18800_ _04098_ _03816_ net353 VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__a21oi_2
X_19780_ _05045_ net212 _05019_ _05031_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__or4_1
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28978_ clknet_leaf_108_clock _01991_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_16992_ decode.regfile.registers_19\[5\] _12679_ _12925_ _12951_ _12545_ VGND VGND
+ VPWR VPWR _12952_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_196_Right_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18731_ _09982_ _09979_ _10010_ memory.csr_read_data_out_reg\[4\] VGND VGND VPWR
+ VPWR _04030_ sky130_fd_sc_hd__o2bb2a_1
X_27929_ clknet_leaf_162_clock _00010_ VGND VGND VPWR VPWR fetch.bht.bhtTable_valid\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15943_ decode.regfile.registers_11\[16\] _11180_ _11183_ decode.regfile.registers_10\[16\]
+ _11278_ VGND VGND VPWR VPWR _11924_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_129_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_Left_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18662_ decode.id_ex_rs1_data_reg\[21\] _03688_ _03943_ VGND VGND VPWR VPWR _03961_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15874_ _11196_ _11855_ _11856_ VGND VGND VPWR VPWR _11857_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17613_ _12822_ decode.regfile.registers_21\[20\] _13164_ _03019_ VGND VGND VPWR
+ VPWR _03020_ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14825_ csr.io_mem_pc\[16\] VGND VGND VPWR VPWR _10868_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18593_ decode.id_ex_rs2_data_reg\[22\] _03746_ _03764_ _03883_ VGND VGND VPWR VPWR
+ _03892_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17544_ _13099_ _13262_ _13182_ decode.regfile.registers_29\[18\] _13490_ VGND VGND
+ VPWR VPWR _13491_ sky130_fd_sc_hd__o221a_1
X_14756_ _10767_ _10797_ _10798_ VGND VGND VPWR VPWR _10799_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13707_ memory.csr_read_data_out_reg\[15\] _09989_ _10055_ _10056_ VGND VGND VPWR
+ VPWR _10057_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_168_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17475_ decode.regfile.registers_0\[17\] _12778_ _13422_ VGND VGND VPWR VPWR _13423_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_28_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14687_ decode.id_ex_pc_reg\[7\] VGND VGND VPWR VPWR _10730_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_28_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19214_ _04281_ _04283_ _03704_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16426_ _11044_ decode.regfile.registers_6\[29\] _11085_ _11318_ VGND VGND VPWR VPWR
+ _12394_ sky130_fd_sc_hd__a211o_1
XFILLER_0_172_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13638_ memory.io_wb_reg_pc\[6\] _09978_ _09995_ _09996_ VGND VGND VPWR VPWR _09997_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_143_Left_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19145_ _04359_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_99_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16357_ decode.regfile.registers_11\[27\] _11181_ _12325_ _12326_ _11187_ VGND VGND
+ VPWR VPWR _12327_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13569_ decode.io_wb_rd\[3\] VGND VGND VPWR VPWR _09934_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15308_ _11294_ _11303_ VGND VGND VPWR VPWR _11304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19076_ _04054_ _03971_ _04321_ _04373_ _04307_ _04338_ VGND VGND VPWR VPWR _04374_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16288_ _11105_ _12258_ _12259_ VGND VGND VPWR VPWR _12260_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18027_ _11019_ _12504_ _12649_ decode.regfile.registers_11\[31\] VGND VGND VPWR
+ VPWR _03423_ sky130_fd_sc_hd__or4b_1
X_15239_ _11235_ VGND VGND VPWR VPWR _11236_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_1314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_82_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19978_ net1792 _05217_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_152_Left_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18929_ _03997_ _03998_ _03999_ _04002_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_197_1082 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21940_ csr.io_mret_vector\[31\] csr.io_mem_pc\[31\] _06481_ VGND VGND VPWR VPWR
+ _06568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_97_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_97_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_173_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21871_ _03449_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23610_ _06140_ net1885 _07941_ VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__mux2_1
X_20822_ _05886_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24590_ _08477_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23541_ net224 _07903_ _07913_ _07907_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20753_ _03755_ _05671_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_20_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_20_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_161_Left_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26260_ _09389_ _09459_ VGND VGND VPWR VPWR _09460_ sky130_fd_sc_hd__nand2_1
X_23472_ decode.id_ex_memread_reg VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__buf_2
XFILLER_0_175_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20684_ _05804_ _05805_ _05807_ _05806_ _05801_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__a32o_1
XFILLER_0_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_210_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25211_ _08834_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_210_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22423_ net96 _07017_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__xor2_1
XFILLER_0_169_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26191_ _09372_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__buf_2
XFILLER_0_169_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25142_ _10949_ _08800_ _10999_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_35_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22354_ fetch.bht.bhtTable_tag\[6\]\[14\] fetch.bht.bhtTable_tag\[7\]\[14\] _06706_
+ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21305_ _06162_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25073_ csr.mcycle\[28\] _08761_ VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22285_ fetch.bht.bhtTable_tag\[0\]\[11\] fetch.bht.bhtTable_tag\[1\]\[11\] fetch.bht.bhtTable_tag\[2\]\[11\]
+ fetch.bht.bhtTable_tag\[3\]\[11\] _06878_ _06621_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__mux4_1
X_24024_ _08183_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__clkbuf_1
X_28901_ clknet_leaf_141_clock _01914_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21236_ _06116_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__clkbuf_1
Xhold250 _10713_ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29881_ clknet_leaf_305_clock _02894_ VGND VGND VPWR VPWR decode.regfile.registers_19\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold261 decode.regfile.registers_7\[13\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_208_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold272 decode.regfile.registers_17\[13\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_208_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold283 decode.regfile.registers_29\[5\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
X_28832_ clknet_leaf_172_clock _01845_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold294 fetch.bht.bhtTable_tag\[15\]\[0\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21167_ _06074_ _06070_ net2290 VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__and3_1
X_20118_ decode.id_ex_imm_reg\[17\] _10806_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__or2_1
X_28763_ clknet_leaf_172_clock _01776_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21098_ _06038_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__buf_2
X_25975_ net2404 _09270_ _09281_ _09277_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27714_ clknet_leaf_20_clock _00743_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20049_ decode.id_ex_imm_reg\[7\] _10730_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__nor2_1
X_24926_ net790 _08662_ _08664_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__o21a_1
XFILLER_0_217_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28694_ clknet_leaf_124_clock _01707_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27645_ clknet_leaf_46_clock _00674_ VGND VGND VPWR VPWR execute.io_reg_pc\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_24857_ _08616_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_101 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 clknet_0_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14610_ _10652_ decode.id_ex_ex_rd_reg\[4\] VGND VGND VPWR VPWR _10653_ sky130_fd_sc_hd__xor2_1
X_23808_ _08059_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_134 _10662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27576_ clknet_leaf_159_clock _00605_ VGND VGND VPWR VPWR csr.io_mem_pc\[17\] sky130_fd_sc_hd__dfxtp_1
X_15590_ _11147_ _10645_ _11578_ _11579_ VGND VGND VPWR VPWR _11580_ sky130_fd_sc_hd__o211ai_1
X_24788_ _08580_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_120_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 execute.io_reg_pc\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _12500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29315_ clknet_leaf_230_clock _02328_ VGND VGND VPWR VPWR decode.regfile.registers_2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14541_ decode.control.io_opcode\[2\] decode.control.io_opcode\[1\] decode.control.io_opcode\[0\]
+ VGND VGND VPWR VPWR _10584_ sky130_fd_sc_hd__and3_1
X_26527_ _09432_ _09602_ VGND VGND VPWR VPWR _09613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23739_ _06101_ net2045 _09907_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29246_ clknet_leaf_234_clock _02259_ VGND VGND VPWR VPWR decode.regfile.registers_0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_17260_ _13091_ _13176_ decode.regfile.registers_27\[11\] _13050_ VGND VGND VPWR
+ VPWR _13214_ sky130_fd_sc_hd__or4_1
X_26458_ _09438_ _09533_ VGND VGND VPWR VPWR _09573_ sky130_fd_sc_hd__nand2_1
X_14472_ _10074_ _10530_ VGND VGND VPWR VPWR _10531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16211_ decode.regfile.registers_10\[23\] _11184_ _12183_ _12184_ VGND VGND VPWR
+ VPWR _12185_ sky130_fd_sc_hd__a22oi_1
X_25409_ _06578_ VGND VGND VPWR VPWR _08950_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29177_ clknet_leaf_238_clock _02190_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__dfxtp_1
X_17191_ decode.regfile.registers_4\[10\] _12548_ _13145_ decode.regfile.registers_5\[10\]
+ _12614_ VGND VGND VPWR VPWR _13146_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26389_ _09532_ VGND VGND VPWR VPWR _09533_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28128_ clknet_leaf_214_clock _01150_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16142_ _12116_ _12117_ _11054_ _11318_ VGND VGND VPWR VPWR _12118_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_49_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28059_ clknet_leaf_198_clock _01081_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16073_ _11756_ decode.regfile.registers_28\[19\] _11871_ _11681_ _11440_ VGND VGND
+ VPWR VPWR _12051_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19901_ _03863_ _03781_ _04254_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__mux2_1
X_15024_ _10981_ VGND VGND VPWR VPWR _11032_ sky130_fd_sc_hd__buf_4
X_19832_ _03829_ _05078_ _05069_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_159_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19763_ _04330_ _04945_ _05037_ _04303_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_53_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16975_ _12934_ _12616_ _12557_ decode.regfile.registers_0\[5\] VGND VGND VPWR VPWR
+ _12935_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_53_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18714_ _03815_ _04012_ net353 VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__a21oi_1
X_15926_ _11489_ decode.regfile.registers_28\[15\] decode.regfile.registers_29\[15\]
+ _11255_ _11246_ VGND VGND VPWR VPWR _11908_ sky130_fd_sc_hd__o221a_1
X_19694_ _04953_ _04970_ _04971_ _04883_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 io_fetch_data[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
X_18645_ decode.id_ex_rs1_data_reg\[21\] _03687_ _03940_ _03914_ _03943_ VGND VGND
+ VPWR VPWR _03944_ sky130_fd_sc_hd__o221a_4
X_15857_ decode.regfile.registers_9\[14\] _11280_ _11134_ _11183_ VGND VGND VPWR VPWR
+ _11840_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_1309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14808_ _10786_ _10789_ _10799_ _10850_ VGND VGND VPWR VPWR _10851_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_204_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18576_ _09929_ csr.io_csr_address\[2\] VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__nor2_1
X_15788_ _11289_ _11771_ _11772_ VGND VGND VPWR VPWR _11773_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17527_ decode.regfile.registers_18\[18\] _12571_ _12561_ VGND VGND VPWR VPWR _13474_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14739_ _10759_ _10769_ csr.io_mem_pc\[28\] VGND VGND VPWR VPWR _10782_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17458_ _10595_ VGND VGND VPWR VPWR _13407_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_129_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16409_ _11076_ decode.regfile.registers_27\[28\] _11869_ VGND VGND VPWR VPWR _12378_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_43_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17389_ _12515_ VGND VGND VPWR VPWR _13339_ sky130_fd_sc_hd__buf_2
XFILLER_0_132_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19128_ _03638_ _04424_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__nor2_2
XFILLER_0_160_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_1310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19059_ _04353_ _04356_ _04272_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22070_ _06664_ _06629_ _06637_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21021_ net2739 _05989_ _05985_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22972_ fetch.bht.bhtTable_target_pc\[4\]\[5\] fetch.bht.bhtTable_target_pc\[5\]\[5\]
+ fetch.bht.bhtTable_target_pc\[6\]\[5\] fetch.bht.bhtTable_target_pc\[7\]\[5\] _07098_
+ _07100_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__mux4_1
X_25760_ _08982_ _09157_ VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24711_ _08539_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__clkbuf_1
X_21923_ _06555_ _06543_ _06544_ _06556_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_195_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25691_ net1467 _09111_ _09118_ _09115_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_195_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_195_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27430_ clknet_leaf_52_clock _00459_ VGND VGND VPWR VPWR decode.id_ex_memwrite_reg
+ sky130_fd_sc_hd__dfxtp_1
X_24642_ net951 execute.io_target_pc\[10\] _08497_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__mux2_1
X_21854_ net2790 _06497_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20805_ _05877_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__clkbuf_1
X_27361_ clknet_leaf_34_clock _00390_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_24573_ _08468_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__clkbuf_1
X_21785_ net1183 csr.io_mem_pc\[31\] _06450_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29100_ clknet_leaf_71_clock _02113_ VGND VGND VPWR VPWR csr._mcycle_T_3\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26312_ net1490 _09448_ _09488_ _09484_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23524_ _10670_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20736_ _05818_ decode.id_ex_rs1_data_reg\[25\] _05759_ VGND VGND VPWR VPWR _05839_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27292_ clknet_leaf_12_clock _00321_ VGND VGND VPWR VPWR decode.regfile.registers_31\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29031_ clknet_leaf_111_clock _02044_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_154_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26243_ net211 VGND VGND VPWR VPWR _09450_ sky130_fd_sc_hd__buf_4
X_23455_ _12765_ _07862_ _07859_ VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__or3b_1
XFILLER_0_163_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20667_ _05794_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22406_ _06650_ _07000_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23386_ _07808_ _07809_ _07081_ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__mux2_1
X_26174_ net1666 _09395_ _09401_ _09394_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20598_ csr.minstret\[22\] _05572_ _05582_ _03555_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22337_ _06685_ _06929_ _06627_ _06931_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__a211oi_1
X_25125_ _06143_ net1744 _08562_ VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25056_ _03555_ csr.mcycle\[23\] _08747_ VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__and3_1
X_29933_ clknet_leaf_341_clock _02946_ VGND VGND VPWR VPWR decode.regfile.registers_21\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_22268_ net222 _06862_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_163_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24007_ net961 execute.io_target_pc\[24\] _07960_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__mux2_1
X_21219_ _10881_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__buf_2
X_29864_ clknet_leaf_298_clock _02877_ VGND VGND VPWR VPWR decode.regfile.registers_19\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_22199_ _06637_ _06788_ _06793_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_40_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28815_ clknet_leaf_110_clock _01828_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_29795_ clknet_leaf_309_clock _02808_ VGND VGND VPWR VPWR decode.regfile.registers_17\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28746_ clknet_leaf_98_clock _01759_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_16760_ _12594_ VGND VGND VPWR VPWR _12724_ sky130_fd_sc_hd__clkbuf_4
X_13972_ _09930_ _10194_ _09933_ _10240_ VGND VGND VPWR VPWR _10241_ sky130_fd_sc_hd__and4b_1
X_25958_ net2508 _09270_ _09272_ _09264_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_122_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15711_ decode.regfile.registers_4\[10\] _11192_ _11410_ _11694_ _11697_ VGND VGND
+ VPWR VPWR _11698_ sky130_fd_sc_hd__o32a_1
XFILLER_0_214_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24909_ net776 _08652_ _08653_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__o21a_1
X_28677_ clknet_leaf_136_clock _01690_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16691_ _12600_ _12648_ _12655_ VGND VGND VPWR VPWR _12656_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25889_ _08962_ _09223_ VGND VGND VPWR VPWR _09232_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18430_ _03715_ _03725_ _03668_ _03728_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__o31a_1
XFILLER_0_154_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27628_ clknet_leaf_154_clock _00657_ VGND VGND VPWR VPWR execute.io_reg_pc\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_15642_ decode.regfile.registers_14\[8\] _11208_ _11629_ _11199_ _11630_ VGND VGND
+ VPWR VPWR _11631_ sky130_fd_sc_hd__a221o_1
XFILLER_0_201_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ execute.io_mem_memtoreg\[1\] VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27559_ clknet_leaf_54_clock _00588_ VGND VGND VPWR VPWR csr.io_mem_pc\[0\] sky130_fd_sc_hd__dfxtp_1
X_15573_ _11079_ VGND VGND VPWR VPWR _11564_ sky130_fd_sc_hd__buf_2
XFILLER_0_51_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17312_ decode.regfile.registers_18\[13\] _12571_ _12561_ VGND VGND VPWR VPWR _13264_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14524_ _10568_ _09890_ VGND VGND VPWR VPWR _10569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18292_ decode.id_ex_rs2_data_reg\[12\] _03605_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_891 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29229_ clknet_leaf_114_clock _02242_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17243_ _13195_ _13196_ _12888_ VGND VGND VPWR VPWR _13197_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_96_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14455_ _10426_ VGND VGND VPWR VPWR _10522_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17174_ _13127_ _13128_ _13129_ VGND VGND VPWR VPWR _13130_ sky130_fd_sc_hd__a21o_1
XFILLER_0_226_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14386_ _10048_ _10474_ VGND VGND VPWR VPWR _10482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16125_ decode.regfile.registers_14\[21\] _11208_ _11274_ decode.regfile.registers_15\[21\]
+ _11202_ VGND VGND VPWR VPWR _12101_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16056_ _12032_ _11364_ _12033_ VGND VGND VPWR VPWR _12034_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_55_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15007_ _11016_ VGND VGND VPWR VPWR _11017_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2409 decode.regfile.registers_1\[5\] VGND VGND VPWR VPWR net2636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19815_ _04805_ _05087_ _04729_ _05041_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__a31o_1
Xhold1708 decode.regfile.registers_21\[4\] VGND VGND VPWR VPWR net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 decode.regfile.registers_22\[19\] VGND VGND VPWR VPWR net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16958_ _10940_ _12706_ decode.regfile.registers_27\[4\] _12507_ VGND VGND VPWR VPWR
+ _12919_ sky130_fd_sc_hd__or4_1
X_19746_ _03894_ _03882_ _04194_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_223_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15909_ decode.regfile.registers_9\[15\] _11280_ _11281_ _11183_ VGND VGND VPWR VPWR
+ _11891_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19677_ _03960_ _04938_ _04191_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__a21o_1
X_16889_ decode.regfile.registers_12\[3\] _12541_ _12722_ _12658_ _12850_ VGND VGND
+ VPWR VPWR _12851_ sky130_fd_sc_hd__o311a_1
XFILLER_0_220_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_205_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18628_ net107 _03665_ _03926_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18559_ _03656_ _03856_ _03701_ _03857_ _03670_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_190_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_190_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21570_ _06305_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_12 _01447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20521_ net923 _05622_ _05667_ _05669_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__a211oi_4
XANTENNA_23 _05857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 _10019_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_45 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_56 _10633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23240_ csr._csr_read_data_T_8\[19\] _06480_ csr.io_mret_vector\[19\] _07621_ _07673_
+ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__o221a_1
XANTENNA_67 _11027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20452_ csr._csr_read_data_T_8\[3\] _05592_ _05516_ _05528_ _05608_ VGND VGND VPWR
+ VPWR _05609_ sky130_fd_sc_hd__a41o_1
XFILLER_0_133_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_78 _11143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 decode.id_ex_rs2_data_reg\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23171_ _07115_ _07607_ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__and2b_1
XFILLER_0_179_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20383_ _05537_ _05538_ _05545_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__and3_1
X_22122_ _06699_ _06704_ _06710_ _06716_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__o31a_2
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput130 net130 VGND VGND VPWR VPWR io_memory_address[8] sky130_fd_sc_hd__clkbuf_4
Xoutput141 net141 VGND VGND VPWR VPWR io_memory_write_data[14] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput152 net152 VGND VGND VPWR VPWR io_memory_write_data[24] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22053_ fetch.bht.bhtTable_tag\[6\]\[22\] fetch.bht.bhtTable_tag\[7\]\[22\] _06645_
+ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__mux2_1
X_26930_ net1935 _09839_ _09845_ _09836_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__o211a_1
Xoutput163 net163 VGND VGND VPWR VPWR io_memory_write_data[5] sky130_fd_sc_hd__clkbuf_4
X_21004_ net2334 _05977_ _05985_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__and3_1
XFILLER_0_227_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_3 _00569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26861_ net1359 _09795_ _09805_ _09799_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_197_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28600_ clknet_leaf_122_clock _01613_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_197_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25812_ _08960_ _09179_ VGND VGND VPWR VPWR _09188_ sky130_fd_sc_hd__nand2_1
X_29580_ clknet_leaf_275_clock _02593_ VGND VGND VPWR VPWR decode.regfile.registers_10\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_26792_ _09751_ VGND VGND VPWR VPWR _09766_ sky130_fd_sc_hd__clkbuf_4
X_28531_ clknet_leaf_239_clock _01544_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25743_ _08966_ _09136_ VGND VGND VPWR VPWR _09148_ sky130_fd_sc_hd__nand2_1
X_22955_ fetch.bht.bhtTable_target_pc\[0\]\[4\] fetch.bht.bhtTable_target_pc\[1\]\[4\]
+ fetch.bht.bhtTable_target_pc\[2\]\[4\] fetch.bht.bhtTable_target_pc\[3\]\[4\] _07108_
+ _07115_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_1147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28462_ clknet_leaf_137_clock _01475_ VGND VGND VPWR VPWR decode.io_id_pc\[20\] sky130_fd_sc_hd__dfxtp_1
X_21906_ _06496_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_168_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25674_ net1580 _09069_ _09107_ _09100_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__o211a_1
X_22886_ net1103 csr.io_mem_pc\[29\] _07335_ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27413_ clknet_leaf_10_clock _00442_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[22\]
+ sky130_fd_sc_hd__dfxtp_2
X_24625_ net1254 execute.io_target_pc\[2\] _07308_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28393_ clknet_leaf_142_clock _01406_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_156_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21837_ _06315_ csr.io_csr_write_address\[1\] csr.io_csr_write_address\[0\] _06472_
+ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27344_ clknet_leaf_44_clock _00373_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[17\]
+ sky130_fd_sc_hd__dfxtp_4
X_21768_ net1861 csr.io_mem_pc\[23\] _06439_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__mux2_1
X_24556_ _08459_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23507_ net93 _07889_ _07894_ _07893_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__o211a_1
X_20719_ _05056_ _05828_ csr.mcycle\[18\] _05537_ _05716_ VGND VGND VPWR VPWR _05829_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27275_ clknet_leaf_11_clock _00304_ VGND VGND VPWR VPWR decode.regfile.registers_30\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24487_ _08113_ net2435 _08422_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__mux2_1
X_21699_ csr.minstret\[16\] csr.minstret\[19\] csr.minstret\[20\] csr.minstret\[21\]
+ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire213 net351 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
X_29014_ clknet_leaf_126_clock _02027_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14240_ _10064_ _10387_ VGND VGND VPWR VPWR _10397_ sky130_fd_sc_hd__nand2_1
X_26226_ net2696 _09419_ _09437_ _09418_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23438_ decode.immGen._imm_T_10\[1\] _07847_ _05206_ VGND VGND VPWR VPWR _07854_
+ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_115_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14171_ net2134 _10346_ _10356_ _10357_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__o211a_1
X_23369_ _07099_ fetch.bht.bhtTable_target_pc\[12\]\[28\] _07071_ VGND VGND VPWR VPWR
+ _07794_ sky130_fd_sc_hd__o21ba_1
X_26157_ _10014_ VGND VGND VPWR VPWR _09389_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_186_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25108_ _08782_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_186_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26088_ net2275 _09343_ _09347_ _09346_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__o211a_1
X_17930_ _12513_ decode.regfile.registers_25\[28\] _03302_ _03328_ VGND VGND VPWR
+ VPWR _03329_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25039_ net2487 _08738_ _08739_ _06419_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_30_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29916_ clknet_leaf_335_clock _02929_ VGND VGND VPWR VPWR decode.regfile.registers_21\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29847_ clknet_leaf_296_clock _02860_ VGND VGND VPWR VPWR decode.regfile.registers_18\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17861_ _02997_ _12767_ _12965_ decode.regfile.registers_29\[26\] _03261_ VGND VGND
+ VPWR VPWR _03262_ sky130_fd_sc_hd__o221a_1
XFILLER_0_218_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19600_ _04509_ _04428_ _04877_ _04881_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__a31o_1
X_16812_ _12774_ VGND VGND VPWR VPWR _12775_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_145_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17792_ _12732_ _03189_ _03190_ _03193_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__a2bb2oi_1
X_29778_ clknet_leaf_295_clock _02791_ VGND VGND VPWR VPWR decode.regfile.registers_16\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19531_ _04281_ _04283_ _04705_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__o21ai_1
X_28729_ clknet_leaf_127_clock _01742_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16743_ _10940_ _10606_ _10937_ _12706_ VGND VGND VPWR VPWR _12707_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_85_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13955_ _10131_ VGND VGND VPWR VPWR _10232_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_85_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19462_ _04747_ _04505_ _04748_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16674_ net209 VGND VGND VPWR VPWR _12639_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13886_ net534 _10180_ _10190_ _10188_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_202 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18413_ execute.io_mem_rd\[1\] _03710_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15625_ _11292_ VGND VGND VPWR VPWR _11614_ sky130_fd_sc_hd__buf_2
XINSDIODE1_213 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19393_ _04359_ _04160_ _04444_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_224 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_235 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_246 net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_257 clknet_0_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18344_ _03642_ decode.id_ex_ex_rs1_reg\[0\] VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_268 _06691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15556_ _11546_ VGND VGND VPWR VPWR _11547_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_44_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_279 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ fetch.btb.btbTable\[8\]\[1\] fetch.btb.btbTable\[9\]\[1\] fetch.btb.btbTable\[10\]\[1\]
+ fetch.btb.btbTable\[11\]\[1\] _09891_ _09888_ VGND VGND VPWR VPWR _10552_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18275_ decode.id_ex_rs2_data_reg\[4\] _03596_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__and2_1
X_15487_ decode.regfile.registers_20\[4\] _11452_ _11223_ _11479_ VGND VGND VPWR VPWR
+ _11480_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_100_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17226_ net514 _12709_ _13138_ _13180_ _12705_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__o221a_1
X_14438_ _09975_ _10507_ VGND VGND VPWR VPWR _10512_ sky130_fd_sc_hd__nand2_1
Xclkbuf_5_19__f_clock clknet_2_2_0_clock VGND VGND VPWR VPWR clknet_5_19__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
Xinput10 io_fetch_data[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 net379 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput32 net444 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_226_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput43 io_memory_read_data[18] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput54 io_memory_read_data[28] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17157_ decode.regfile.registers_10\[9\] _12790_ _12792_ VGND VGND VPWR VPWR _13113_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold805 fetch.bht.bhtTable_target_pc\[9\]\[11\] VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__dlygate4sd3_1
Xinput65 io_memory_read_data[9] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlymetal6s2s_1
X_14369_ _09999_ _10464_ VGND VGND VPWR VPWR _10472_ sky130_fd_sc_hd__nand2_1
Xhold816 fetch.bht.bhtTable_tag\[8\]\[11\] VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__dlygate4sd3_1
X_16108_ decode.regfile.registers_22\[20\] _11096_ _12083_ _12084_ _11232_ VGND VGND
+ VPWR VPWR _12085_ sky130_fd_sc_hd__a221oi_2
Xhold827 decode.regfile.registers_14\[30\] VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 _01118_ VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 fetch.bht.bhtTable_tag\[4\]\[7\] VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17088_ _12915_ decode.regfile.registers_25\[7\] _13045_ _12812_ VGND VGND VPWR VPWR
+ _13046_ sky130_fd_sc_hd__or4_1
XFILLER_0_161_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16039_ decode.regfile.registers_14\[19\] _11360_ _11274_ decode.regfile.registers_15\[19\]
+ _11202_ VGND VGND VPWR VPWR _12017_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2206 decode.regfile.registers_10\[0\] VGND VGND VPWR VPWR net2433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2217 csr.minstret\[13\] VGND VGND VPWR VPWR net2444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2228 decode.regfile.registers_16\[29\] VGND VGND VPWR VPWR net2455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2239 decode.regfile.registers_6\[24\] VGND VGND VPWR VPWR net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_200_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1505 fetch.bht.bhtTable_target_pc\[13\]\[12\] VGND VGND VPWR VPWR net1732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1516 decode.regfile.registers_20\[16\] VGND VGND VPWR VPWR net1743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 fetch.bht.bhtTable_tag\[13\]\[12\] VGND VGND VPWR VPWR net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 decode.regfile.registers_18\[22\] VGND VGND VPWR VPWR net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1549 fetch.bht.bhtTable_target_pc\[8\]\[21\] VGND VGND VPWR VPWR net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19729_ _04295_ _04362_ _04629_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_0_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_192_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22740_ _07262_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22671_ _07207_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__buf_2
XFILLER_0_220_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24410_ _08382_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__clkbuf_1
X_21622_ csr.minstret\[6\] csr.minstret\[7\] _06342_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25390_ net876 _08928_ _08936_ _08927_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24341_ _08103_ net2031 _06187_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__mux2_1
X_21553_ _06124_ net1716 _06295_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20504_ csr._minstret_T_3\[41\] _05577_ _05578_ _05654_ VGND VGND VPWR VPWR _05655_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24272_ _08311_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27060_ clknet_leaf_331_clock _00089_ VGND VGND VPWR VPWR decode.regfile.registers_24\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21484_ _06113_ net1746 _06252_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23223_ _07555_ fetch.bht.bhtTable_target_pc\[15\]\[19\] _07656_ VGND VGND VPWR VPWR
+ _07657_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26011_ _08933_ _09297_ VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20435_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23154_ fetch.bht.bhtTable_target_pc\[4\]\[15\] fetch.bht.bhtTable_target_pc\[5\]\[15\]
+ fetch.bht.bhtTable_target_pc\[6\]\[15\] fetch.bht.bhtTable_target_pc\[7\]\[15\]
+ _07555_ _07114_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_228_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20366_ csr.io_csr_address\[11\] _05526_ _05523_ _05520_ _05528_ VGND VGND VPWR VPWR
+ _05529_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_228_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22105_ _06691_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_149_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23085_ fetch.bht.bhtTable_target_pc\[4\]\[11\] fetch.bht.bhtTable_target_pc\[5\]\[11\]
+ fetch.bht.bhtTable_target_pc\[6\]\[11\] fetch.bht.bhtTable_target_pc\[7\]\[11\]
+ _07108_ _07125_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__mux4_1
X_27962_ clknet_leaf_214_clock _00984_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20297_ decode.id_ex_pc_reg\[18\] _05470_ _05416_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_224_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29701_ clknet_leaf_286_clock _02714_ VGND VGND VPWR VPWR decode.regfile.registers_14\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_224_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22036_ _00002_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26913_ net892 _09796_ _09834_ _09825_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_8_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27893_ clknet_leaf_19_clock _00922_ VGND VGND VPWR VPWR csr._mcycle_T_2\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29632_ clknet_5_20__leaf_clock _02645_ VGND VGND VPWR VPWR decode.regfile.registers_12\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26844_ _09794_ VGND VGND VPWR VPWR _09796_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29563_ clknet_leaf_251_clock _02576_ VGND VGND VPWR VPWR decode.regfile.registers_10\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26775_ net2220 _09752_ _09756_ _09743_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__o211a_1
X_23987_ net865 execute.io_target_pc\[14\] _08164_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__mux2_1
X_28514_ clknet_leaf_211_clock _01527_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13740_ memory.io_wb_reg_pc\[20\] _09946_ _09947_ _10084_ VGND VGND VPWR VPWR _10085_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25726_ net1148 _09125_ _09138_ _09129_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22938_ fetch.bht.bhtTable_target_pc\[4\]\[3\] fetch.bht.bhtTable_target_pc\[5\]\[3\]
+ fetch.bht.bhtTable_target_pc\[6\]\[3\] fetch.bht.bhtTable_target_pc\[7\]\[3\] _07106_
+ _07386_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__mux4_1
X_29494_ clknet_leaf_263_clock _02507_ VGND VGND VPWR VPWR decode.regfile.registers_7\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_179_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28445_ clknet_leaf_145_clock _01458_ VGND VGND VPWR VPWR decode.io_id_pc\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25657_ net2494 _09095_ _09098_ _09087_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__o211a_1
X_13671_ net588 _09938_ _10026_ _10020_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_80_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22869_ net944 csr.io_mem_pc\[21\] _07324_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15410_ _11093_ VGND VGND VPWR VPWR _11404_ sky130_fd_sc_hd__buf_2
X_24608_ _08486_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_175_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28376_ clknet_leaf_187_clock _01389_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_175_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16390_ _12358_ decode.regfile.registers_7\[28\] _11378_ VGND VGND VPWR VPWR _12359_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25588_ _08990_ VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_117_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27327_ clknet_5_6__leaf_clock _00356_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_15341_ decode.regfile.registers_25\[1\] _11333_ _11336_ decode.regfile.registers_24\[1\]
+ VGND VGND VPWR VPWR _11337_ sky130_fd_sc_hd__o22a_1
X_24539_ _08099_ net2114 _09902_ VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18060_ _03451_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__clkbuf_1
X_15272_ _11047_ _11111_ _10651_ _10633_ VGND VGND VPWR VPWR _11268_ sky130_fd_sc_hd__and4_2
X_27258_ clknet_leaf_8_clock _00287_ VGND VGND VPWR VPWR decode.regfile.registers_30\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17011_ _12532_ _10593_ _12559_ decode.regfile.registers_0\[6\] VGND VGND VPWR VPWR
+ _12970_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_78_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26209_ net200 VGND VGND VPWR VPWR _09426_ sky130_fd_sc_hd__buf_4
X_14223_ _10015_ _10387_ VGND VGND VPWR VPWR _10388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27189_ clknet_leaf_6_clock _00218_ VGND VGND VPWR VPWR decode.regfile.registers_28\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14154_ _10036_ _10342_ VGND VGND VPWR VPWR _10348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18962_ decode.id_ex_imm_reg\[1\] VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__buf_4
X_14085_ _10053_ _10299_ VGND VGND VPWR VPWR _10308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ decode.regfile.registers_4\[28\] _12547_ _12531_ decode.regfile.registers_5\[28\]
+ _12625_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18893_ _03957_ _03960_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_37_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17844_ _11021_ _12491_ _12666_ decode.regfile.registers_14\[26\] _12670_ VGND VGND
+ VPWR VPWR _03245_ sky130_fd_sc_hd__o32a_1
XFILLER_0_191_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17775_ _13407_ decode.regfile.registers_25\[24\] _13482_ _12811_ VGND VGND VPWR
+ VPWR _03178_ sky130_fd_sc_hd__or4_1
X_14987_ _10998_ VGND VGND VPWR VPWR _11004_ sky130_fd_sc_hd__buf_2
XFILLER_0_221_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19514_ _04290_ _04273_ _04410_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__and3_1
X_16726_ _11025_ _12690_ _10604_ VGND VGND VPWR VPWR _12691_ sky130_fd_sc_hd__and3_1
X_13938_ _10069_ _10210_ VGND VGND VPWR VPWR _10222_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19445_ _04732_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__buf_1
XFILLER_0_88_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16657_ _12621_ VGND VGND VPWR VPWR _12622_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_102_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13869_ net1582 _10180_ _10181_ _10175_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15608_ decode.regfile.registers_19\[7\] _11406_ _11325_ _11597_ VGND VGND VPWR VPWR
+ _11598_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19376_ _04131_ _04662_ _04663_ _04665_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__o211a_1
X_16588_ _12552_ VGND VGND VPWR VPWR _12553_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18327_ _03629_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15539_ _10956_ decode.regfile.registers_22\[6\] _11093_ _11264_ _11265_ VGND VGND
+ VPWR VPWR _11530_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_63_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18258_ _03589_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17209_ _12755_ VGND VGND VPWR VPWR _13164_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18189_ _03522_ _03525_ _03526_ _10582_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__o31a_1
XFILLER_0_142_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold602 fetch.bht.bhtTable_target_pc\[4\]\[6\] VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold613 fetch.bht.bhtTable_tag\[3\]\[6\] VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__dlygate4sd3_1
X_20220_ decode.id_ex_pc_reg\[0\] _05412_ _05413_ _05414_ VGND VGND VPWR VPWR _00652_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold624 decode.regfile.registers_29\[14\] VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold635 fetch.bht.bhtTable_target_pc\[1\]\[23\] VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold646 fetch.bht.bhtTable_tag\[4\]\[3\] VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold657 csr.mscratch\[9\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 fetch.bht.bhtTable_target_pc\[1\]\[14\] VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd3_1
X_20151_ decode.id_ex_imm_reg\[20\] _10867_ _10798_ decode.id_ex_imm_reg\[21\] _05353_
+ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold679 fetch.bht.bhtTable_tag\[2\]\[3\] VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2003 fetch.bht.bhtTable_tag\[7\]\[7\] VGND VGND VPWR VPWR net2230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20082_ _05295_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__and2b_1
XFILLER_0_176_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2014 decode.regfile.registers_21\[28\] VGND VGND VPWR VPWR net2241 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2025 decode.regfile.registers_7\[19\] VGND VGND VPWR VPWR net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2036 decode.regfile.registers_1\[25\] VGND VGND VPWR VPWR net2263 sky130_fd_sc_hd__dlygate4sd3_1
X_23910_ net890 _08068_ _08119_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__mux2_1
Xhold1302 decode.regfile.registers_15\[19\] VGND VGND VPWR VPWR net1529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2047 decode.regfile.registers_15\[21\] VGND VGND VPWR VPWR net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1313 fetch.bht.bhtTable_target_pc\[10\]\[18\] VGND VGND VPWR VPWR net1540 sky130_fd_sc_hd__dlygate4sd3_1
X_24890_ csr.mcycle\[28\] csr.mcycle\[27\] csr.mcycle\[30\] csr.mcycle\[29\] VGND
+ VGND VPWR VPWR _08639_ sky130_fd_sc_hd__and4_1
Xhold2058 decode.regfile.registers_14\[21\] VGND VGND VPWR VPWR net2285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1003 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1324 fetch.bht.bhtTable_target_pc\[13\]\[8\] VGND VGND VPWR VPWR net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2069 fetch.bht.bhtTable_target_pc\[7\]\[1\] VGND VGND VPWR VPWR net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 fetch.bht.bhtTable_target_pc\[13\]\[25\] VGND VGND VPWR VPWR net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 fetch.bht.bhtTable_tag\[9\]\[21\] VGND VGND VPWR VPWR net1573 sky130_fd_sc_hd__dlygate4sd3_1
X_23841_ _08081_ net2288 _08079_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__mux2_1
Xhold1357 fetch.bht.bhtTable_target_pc\[0\]\[5\] VGND VGND VPWR VPWR net1584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1368 fetch.bht.bhtTable_tag\[6\]\[9\] VGND VGND VPWR VPWR net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1379 fetch.bht.bhtTable_tag\[14\]\[9\] VGND VGND VPWR VPWR net1606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26560_ _09621_ VGND VGND VPWR VPWR _09632_ sky130_fd_sc_hd__clkbuf_4
X_23772_ _06134_ net1232 _08030_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__mux2_1
X_20984_ execute.io_reg_pc\[17\] _05965_ _05973_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__and3_1
XFILLER_0_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25511_ _08962_ _09005_ VGND VGND VPWR VPWR _09014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22723_ _03546_ _07248_ _07253_ _03551_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__nor4_1
XFILLER_0_211_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26491_ _09396_ _09589_ VGND VGND VPWR VPWR _09593_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28230_ clknet_leaf_56_clock _01252_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_2
X_25442_ net515 _08951_ _08971_ _08972_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__o211a_1
X_22654_ csr._mcycle_T_2\[4\] _07210_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_217_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21605_ net2608 _06328_ _06330_ _06331_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__a211oi_1
X_28161_ clknet_leaf_67_clock net1159 VGND VGND VPWR VPWR csr._csr_read_data_T_9\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22585_ csr._minstret_T_3\[43\] csr._minstret_T_3\[42\] csr._minstret_T_3\[41\] _07162_
+ _07148_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__a41o_1
X_25373_ net763 _08906_ _08924_ _07247_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27112_ clknet_leaf_358_clock _00141_ VGND VGND VPWR VPWR decode.regfile.registers_25\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24324_ _08338_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28092_ clknet_leaf_188_clock _01114_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_170_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21536_ _06107_ net2002 _06284_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27043_ clknet_leaf_346_clock _00072_ VGND VGND VPWR VPWR decode.regfile.registers_23\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24255_ _08083_ net1783 _08300_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__mux2_1
X_21467_ _10964_ _06248_ _10915_ _10908_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_177_Right_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_226_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23206_ fetch.bht.bhtTable_target_pc\[8\]\[18\] fetch.bht.bhtTable_target_pc\[9\]\[18\]
+ _07067_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_189_Left_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20418_ _05534_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__clkbuf_4
X_24186_ _08267_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__clkbuf_1
X_21398_ _06212_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23137_ _07574_ _07575_ _07122_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__mux2_1
X_20349_ _10684_ decode.id_ex_pc_reg\[31\] _05508_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__or3_1
X_28994_ clknet_leaf_134_clock _02007_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23068_ fetch.bht.bhtTable_target_pc\[15\]\[10\] _07407_ VGND VGND VPWR VPWR _07511_
+ sky130_fd_sc_hd__or2b_1
X_27945_ clknet_leaf_211_clock _00967_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22019_ net1158 _06571_ _06614_ _06605_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__o211a_1
X_14910_ _10912_ _10913_ _10921_ _10941_ VGND VGND VPWR VPWR _10942_ sky130_fd_sc_hd__and4bb_1
X_27876_ clknet_leaf_56_clock _00905_ VGND VGND VPWR VPWR csr.io_trapped sky130_fd_sc_hd__dfxtp_1
X_15890_ _11403_ _11868_ _11870_ _11872_ VGND VGND VPWR VPWR _11873_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_333_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_333_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold2570 csr._mcycle_T_2\[31\] VGND VGND VPWR VPWR net2797 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _10881_ _10816_ VGND VGND VPWR VPWR _10884_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_106_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29615_ clknet_leaf_279_clock _02628_ VGND VGND VPWR VPWR decode.regfile.registers_11\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_26827_ _09430_ _09776_ VGND VGND VPWR VPWR _09786_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_198_Left_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1880 fetch.bht.bhtTable_target_pc\[9\]\[30\] VGND VGND VPWR VPWR net2107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17560_ decode.regfile.registers_10\[19\] _12790_ _13495_ _02967_ _12878_ VGND VGND
+ VPWR VPWR _02968_ sky130_fd_sc_hd__o221a_1
X_29546_ clknet_leaf_266_clock _02559_ VGND VGND VPWR VPWR decode.regfile.registers_9\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1891 fetch.bht.bhtTable_tag\[7\]\[25\] VGND VGND VPWR VPWR net2118 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_177_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ csr.io_mem_pc\[4\] csr.io_mem_pc\[5\] _09894_ VGND VGND VPWR VPWR _10815_
+ sky130_fd_sc_hd__and3_1
X_26758_ _09436_ _09708_ VGND VGND VPWR VPWR _09746_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_177_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16511_ decode.regfile.registers_21\[31\] _11267_ _11098_ _11227_ _12476_ VGND VGND
+ VPWR VPWR _12477_ sky130_fd_sc_hd__o311a_1
X_25709_ net2327 _09125_ _09127_ _09129_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__o211a_1
X_13723_ net1719 _10027_ _10070_ _10020_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_67_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17491_ decode.regfile.registers_19\[17\] _12678_ _13418_ _13438_ _12906_ VGND VGND
+ VPWR VPWR _13439_ sky130_fd_sc_hd__o221a_1
X_29477_ clknet_leaf_263_clock _02490_ VGND VGND VPWR VPWR decode.regfile.registers_7\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_348_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_348_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26689_ _09443_ _09664_ VGND VGND VPWR VPWR _09706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19230_ _03637_ decode.id_ex_aluop_reg\[1\] decode.id_ex_aluop_reg\[3\] decode.id_ex_aluop_reg\[2\]
+ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__or4_4
X_28428_ clknet_leaf_246_clock _01441_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_16442_ decode.regfile.registers_23\[29\] _11088_ _12384_ _12409_ VGND VGND VPWR
+ VPWR _12410_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13654_ _09995_ _09978_ memory.io_wb_reg_pc\[8\] VGND VGND VPWR VPWR _10011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19161_ _04024_ _04447_ _04446_ _04457_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28359_ clknet_leaf_223_clock _01372_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16373_ _11756_ decode.regfile.registers_28\[27\] _11871_ _11037_ _11448_ VGND VGND
+ VPWR VPWR _12343_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_6_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13585_ _09949_ VGND VGND VPWR VPWR _09950_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18112_ _03483_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15324_ decode.regfile.registers_14\[1\] _11208_ _11274_ decode.regfile.registers_15\[1\]
+ _11319_ VGND VGND VPWR VPWR _11320_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19092_ _04325_ _04388_ _04308_ _04389_ _04306_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_186_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18043_ _12515_ _03436_ _03437_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__a31o_1
X_15255_ _11250_ VGND VGND VPWR VPWR _11251_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14206_ net573 _10376_ _10378_ _10369_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_39_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15186_ _11182_ VGND VGND VPWR VPWR _11183_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14137_ _09984_ _10333_ VGND VGND VPWR VPWR _10338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_1316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19994_ net2711 _05219_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18945_ _04243_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__clkbuf_4
X_14068_ _10008_ _10288_ VGND VGND VPWR VPWR _10298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_219_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18876_ _04053_ _04057_ _04076_ _04170_ _04174_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__a311o_1
XFILLER_0_158_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17827_ _12524_ _12568_ _12535_ _12674_ decode.regfile.registers_16\[26\] VGND VGND
+ VPWR VPWR _03228_ sky130_fd_sc_hd__a32o_1
XFILLER_0_221_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17758_ decode.regfile.registers_9\[24\] _12604_ _12532_ _12776_ VGND VGND VPWR VPWR
+ _03161_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16709_ _12673_ VGND VGND VPWR VPWR _12674_ sky130_fd_sc_hd__clkbuf_4
X_17689_ decode.regfile.registers_16\[22\] _12575_ _03077_ _03093_ _12578_ VGND VGND
+ VPWR VPWR _03094_ sky130_fd_sc_hd__o221a_1
XFILLER_0_175_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19428_ _04166_ _04164_ _04684_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19359_ _04296_ _04646_ _04649_ _04349_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22370_ _06956_ _06964_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_212_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_212_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21321_ net1227 csr.io_mem_pc\[18\] _06168_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24040_ net1481 execute.io_target_pc\[8\] _08187_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__mux2_1
X_21252_ _06127_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold410 decode.regfile.registers_3\[0\] VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold421 execute.csr_write_data_out_reg\[4\] VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold432 decode.regfile.registers_21\[10\] VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__dlygate4sd3_1
X_20203_ _05399_ _05400_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__nor2_1
Xhold443 decode.regfile.registers_22\[3\] VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold454 decode.regfile.registers_7\[10\] VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__dlygate4sd3_1
X_21183_ _06086_ _06082_ net638 VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__and3_1
Xhold465 fetch.bht.bhtTable_tag\[12\]\[17\] VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold476 decode.regfile.registers_29\[9\] VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _01259_ VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap195 _10121_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_221_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20134_ _05339_ _05341_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__nand2_1
Xhold498 decode.regfile.registers_21\[2\] VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25991_ _09263_ VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__clkbuf_4
X_27730_ clknet_leaf_69_clock _00759_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20065_ decode.id_ex_imm_reg\[10\] decode.id_ex_pc_reg\[10\] VGND VGND VPWR VPWR
+ _05282_ sky130_fd_sc_hd__nor2_1
X_24942_ csr._mcycle_T_3\[49\] csr._mcycle_T_3\[48\] _08672_ _07148_ VGND VGND VPWR
+ VPWR _08675_ sky130_fd_sc_hd__a31o_1
Xhold1110 decode.regfile.registers_7\[7\] VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1121 decode.regfile.registers_21\[3\] VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 decode.regfile.registers_20\[7\] VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27661_ clknet_leaf_26_clock _00690_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24873_ _08624_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__clkbuf_1
Xhold1143 csr._mcycle_T_2\[5\] VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__clkbuf_2
Xhold1154 fetch.bht.bhtTable_target_pc\[8\]\[5\] VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1165 csr._minstret_T_3\[60\] VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__dlygate4sd3_1
X_29400_ clknet_leaf_246_clock _02413_ VGND VGND VPWR VPWR decode.regfile.registers_4\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1176 fetch.bht.bhtTable_tag\[6\]\[25\] VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26612_ net2484 _09623_ _09661_ _09660_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1187 fetch.bht.bhtTable_target_pc\[0\]\[16\] VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__dlygate4sd3_1
X_23824_ execute.io_target_pc\[10\] VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__buf_2
X_27592_ clknet_leaf_147_clock _00621_ VGND VGND VPWR VPWR execute.io_target_pc\[1\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_219_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 fetch.bht.bhtTable_tag\[8\]\[25\] VGND VGND VPWR VPWR net1425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_219_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29331_ clknet_leaf_225_clock _02344_ VGND VGND VPWR VPWR decode.regfile.registers_2\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_26543_ _09621_ VGND VGND VPWR VPWR _09623_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23755_ _06117_ net1331 _09907_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20967_ execute.io_reg_pc\[9\] _05965_ _05961_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22706_ net1957 _07236_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_172_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29262_ clknet_leaf_223_clock _02275_ VGND VGND VPWR VPWR decode.regfile.registers_0\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26474_ net1802 _09578_ _09583_ _09582_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_172_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23686_ _07993_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20898_ _05928_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28213_ clknet_leaf_83_clock net1835 VGND VGND VPWR VPWR csr.mscratch\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25425_ _08960_ _08946_ VGND VGND VPWR VPWR _08961_ sky130_fd_sc_hd__nand2_1
X_22637_ _07201_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__clkbuf_2
X_29193_ clknet_leaf_238_clock _02206_ VGND VGND VPWR VPWR fetch.btb.btbTable\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28144_ clknet_leaf_197_clock _01166_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25356_ _08912_ _08907_ VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22568_ _06377_ _07150_ _07153_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__nor3_1
XFILLER_0_106_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24307_ _08329_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21519_ _06277_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__clkbuf_1
X_28075_ clknet_leaf_238_clock _01097_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25287_ _08869_ decode.regfile.registers_0\[5\] VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22499_ csr.io_mret_vector\[0\] VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15040_ _11036_ VGND VGND VPWR VPWR _11037_ sky130_fd_sc_hd__clkbuf_8
X_27026_ clknet_leaf_331_clock _00055_ VGND VGND VPWR VPWR decode.regfile.registers_23\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_24238_ _08066_ net2100 _08289_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24169_ _08258_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16991_ decode.regfile.registers_17\[5\] _12580_ _12826_ _12950_ VGND VGND VPWR VPWR
+ _12951_ sky130_fd_sc_hd__o211a_1
X_28977_ clknet_leaf_103_clock _01990_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18730_ _04027_ _04028_ _04022_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__o21a_1
X_15942_ decode.regfile.registers_8\[16\] _11284_ _11287_ decode.regfile.registers_9\[16\]
+ _11131_ VGND VGND VPWR VPWR _11923_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_129_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27928_ clknet_leaf_36_clock _00957_ VGND VGND VPWR VPWR execute.io_mem_rd\[4\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_129_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _10086_ _03772_ _03774_ _03955_ _03959_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_204_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15873_ decode.regfile.registers_13\[14\] _11196_ _11198_ VGND VGND VPWR VPWR _11856_
+ sky130_fd_sc_hd__o21ai_1
X_27859_ clknet_leaf_317_clock _00888_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14824_ decode.id_ex_pc_reg\[20\] VGND VGND VPWR VPWR _10867_ sky130_fd_sc_hd__buf_4
X_17612_ decode.regfile.registers_20\[20\] _12771_ _03018_ _12537_ VGND VGND VPWR
+ VPWR _03019_ sky130_fd_sc_hd__a211o_1
XFILLER_0_192_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18592_ _03797_ _03885_ _03890_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_203_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_287_clock clknet_5_20__leaf_clock VGND VGND VPWR VPWR clknet_leaf_287_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17543_ _13221_ _13486_ _13488_ _13489_ VGND VGND VPWR VPWR _13490_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_1231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14755_ decode.id_ex_pc_reg\[21\] VGND VGND VPWR VPWR _10798_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29529_ clknet_leaf_251_clock _02542_ VGND VGND VPWR VPWR decode.regfile.registers_8\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13706_ _10012_ memory.io_wb_aluresult\[15\] _09978_ memory.io_wb_reg_pc\[15\] _09995_
+ VGND VGND VPWR VPWR _10056_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_169_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17474_ decode.regfile.registers_1\[17\] net215 _12934_ VGND VGND VPWR VPWR _13422_
+ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_1_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_1_clock
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_213_Right_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14686_ execute.io_target_pc\[15\] _10682_ execute.io_target_pc\[14\] _10702_ _10728_
+ VGND VGND VPWR VPWR _10729_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_210_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_210_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19213_ _04371_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16425_ decode.regfile.registers_5\[29\] _11280_ _11139_ _11466_ _12392_ VGND VGND
+ VPWR VPWR _12393_ sky130_fd_sc_hd__a311o_1
XFILLER_0_183_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13637_ _09943_ memory.io_wb_aluresult\[6\] _09981_ memory.io_wb_readdata\[6\] VGND
+ VGND VPWR VPWR _09996_ sky130_fd_sc_hd__a22o_1
XFILLER_0_229_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19144_ _04321_ _04425_ _04270_ _04429_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_60_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16356_ _11070_ _11470_ decode.regfile.registers_10\[27\] _11382_ VGND VGND VPWR
+ VPWR _12326_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_99_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13568_ decode.io_wb_rd\[4\] decode.io_wb_regwrite VGND VGND VPWR VPWR _09933_ sky130_fd_sc_hd__and2_2
XFILLER_0_87_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15307_ decode.regfile.registers_2\[1\] _11296_ _11297_ _11121_ _11302_ VGND VGND
+ VPWR VPWR _11303_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19075_ decode.id_ex_rs1_data_reg\[1\] net247 _04005_ _04001_ VGND VGND VPWR VPWR
+ _04373_ sky130_fd_sc_hd__o211a_2
XFILLER_0_125_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16287_ decode.regfile.registers_18\[25\] _10640_ _11112_ _10651_ _10633_ VGND VGND
+ VPWR VPWR _12259_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13499_ _09880_ VGND VGND VPWR VPWR _09881_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_225_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_225_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18026_ decode.regfile.registers_10\[31\] _12600_ _03420_ _03421_ VGND VGND VPWR
+ VPWR _03422_ sky130_fd_sc_hd__a22oi_2
X_15238_ _10657_ _10957_ _11217_ _10662_ VGND VGND VPWR VPWR _11235_ sky130_fd_sc_hd__or4b_2
XFILLER_0_160_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15169_ _11165_ VGND VGND VPWR VPWR _11166_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19977_ net477 _05217_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18928_ _04171_ _04173_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__nor2_2
XFILLER_0_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18859_ net101 _03665_ _04157_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_206_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21870_ _06493_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__buf_2
XFILLER_0_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20821_ net129 _05879_ _05875_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__and3_1
XFILLER_0_221_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23540_ net2211 _07904_ _07901_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20752_ _03741_ _05671_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_214_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_214_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23471_ net15 _07861_ _07872_ _07865_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__o211a_1
X_20683_ _05621_ _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25210_ _08049_ net1294 _08041_ VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22422_ _06699_ _07010_ _07016_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_116_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_210_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26190_ _10073_ VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25141_ _10946_ _10944_ _10964_ _10665_ VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__and4b_1
X_22353_ _06649_ _06947_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__or2b_1
XFILLER_0_182_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21304_ net1112 _10878_ _06157_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__mux2_1
X_22284_ fetch.bht.bhtTable_tag\[4\]\[11\] fetch.bht.bhtTable_tag\[5\]\[11\] fetch.bht.bhtTable_tag\[6\]\[11\]
+ fetch.bht.bhtTable_tag\[7\]\[11\] _06878_ _06677_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__mux4_1
X_25072_ csr._mcycle_T_2\[28\] _08703_ _08761_ csr.mcycle\[28\] VGND VGND VPWR VPWR
+ _08762_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28900_ clknet_leaf_128_clock _01913_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24023_ net867 execute.io_target_pc\[0\] _08014_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__mux2_1
X_21235_ net842 _06115_ _09912_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold240 decode.regfile.registers_30\[7\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
X_29880_ clknet_leaf_315_clock _02893_ VGND VGND VPWR VPWR decode.regfile.registers_19\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold251 decode.regfile.registers_31\[24\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_1
Xhold262 decode.regfile.registers_25\[8\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_208_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold273 decode.regfile.registers_29\[31\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28831_ clknet_leaf_179_clock _01844_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_165_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold284 decode.regfile.registers_23\[8\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
X_21166_ _06077_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold295 decode.regfile.registers_27\[1\] VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
X_20117_ decode.id_ex_imm_reg\[17\] _10806_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__nand2_1
X_28762_ clknet_leaf_129_clock _01775_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_21097_ _06037_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__clkbuf_4
X_25974_ _08970_ _09241_ VGND VGND VPWR VPWR _09281_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_161_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27713_ clknet_leaf_19_clock _00742_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_20048_ decode.id_ex_imm_reg\[5\] _10704_ _05262_ _05264_ VGND VGND VPWR VPWR _05268_
+ sky130_fd_sc_hd__o211ai_1
X_24925_ net790 _08662_ _06318_ VGND VGND VPWR VPWR _08664_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28693_ clknet_leaf_141_clock _01706_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27644_ clknet_leaf_155_clock _00673_ VGND VGND VPWR VPWR execute.io_reg_pc\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_24856_ _06134_ net1334 _08607_ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_102 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_198_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23807_ _08057_ net2041 _08058_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_113 net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27575_ clknet_leaf_159_clock _00604_ VGND VGND VPWR VPWR csr.io_mem_pc\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_124 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24787_ _08081_ net1789 _08574_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_135 _11035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21999_ csr.mscratch\[22\] _06601_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_120_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29314_ clknet_leaf_231_clock _02327_ VGND VGND VPWR VPWR decode.regfile.registers_2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _12500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14540_ decode.control.io_opcode\[4\] decode.control.io_opcode\[5\] decode.control.io_opcode\[6\]
+ VGND VGND VPWR VPWR _10583_ sky130_fd_sc_hd__and3b_2
X_26526_ net2661 _09605_ _09612_ _09608_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__o211a_1
X_23738_ _08020_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29245_ clknet_leaf_231_clock _02258_ VGND VGND VPWR VPWR decode.regfile.registers_0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26457_ net2168 _09561_ _09572_ _09567_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__o211a_1
X_14471_ _10505_ VGND VGND VPWR VPWR _10530_ sky130_fd_sc_hd__buf_2
XFILLER_0_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23669_ _07959_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16210_ decode.regfile.registers_8\[23\] _11285_ _11365_ decode.regfile.registers_9\[23\]
+ _11382_ VGND VGND VPWR VPWR _12184_ sky130_fd_sc_hd__o221a_1
X_25408_ _08948_ _08946_ VGND VGND VPWR VPWR _08949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29176_ clknet_leaf_239_clock _02189_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__dfxtp_4
X_17190_ _12934_ VGND VGND VPWR VPWR _13145_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26388_ _10373_ _10195_ _09932_ _08903_ VGND VGND VPWR VPWR _09532_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28127_ clknet_leaf_67_clock _01149_ VGND VGND VPWR VPWR csr.io_ecause\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16141_ decode.regfile.registers_13\[21\] _11276_ VGND VGND VPWR VPWR _12117_ sky130_fd_sc_hd__nand2_1
X_25339_ _08900_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28058_ clknet_leaf_194_clock _01080_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_16072_ _11679_ decode.regfile.registers_27\[19\] _11869_ VGND VGND VPWR VPWR _12050_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_51_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15023_ _10962_ _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__a31o_1
X_27009_ clknet_leaf_342_clock _00038_ VGND VGND VPWR VPWR decode.regfile.registers_22\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_19900_ _03861_ _03863_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__or2b_1
X_19831_ _05101_ _05102_ net213 VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__and3_1
XFILLER_0_209_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19762_ _04305_ _05036_ _04371_ _04851_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_53_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16974_ _12530_ VGND VGND VPWR VPWR _12934_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_53_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18713_ net122 _03663_ _04011_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__o21ai_2
X_15925_ _11251_ _11259_ decode.regfile.registers_27\[15\] _11876_ _11906_ VGND VGND
+ VPWR VPWR _11907_ sky130_fd_sc_hd__o32a_1
XFILLER_0_95_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19693_ _04905_ _04576_ _04571_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__and3_1
XFILLER_0_189_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput8 io_fetch_data[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_0_95_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15856_ decode.regfile.registers_11\[14\] _11070_ _11470_ _11278_ VGND VGND VPWR
+ VPWR _11839_ sky130_fd_sc_hd__a31o_1
X_18644_ _03816_ _03942_ net353 VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14807_ decode.id_ex_pc_reg\[21\] _10767_ _10797_ _10802_ _10849_ VGND VGND VPWR
+ VPWR _10850_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_99_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15787_ decode.regfile.registers_7\[12\] _11378_ _11170_ decode.regfile.registers_6\[12\]
+ _11166_ VGND VGND VPWR VPWR _11772_ sky130_fd_sc_hd__a221oi_2
X_18575_ csr.io_csr_address\[3\] _09935_ _03733_ _03730_ _03736_ VGND VGND VPWR VPWR
+ _03874_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_8_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14738_ csr.io_mem_pc\[27\] csr.io_mem_pc\[28\] _10769_ VGND VGND VPWR VPWR _10781_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17526_ decode.regfile.registers_17\[18\] _12901_ _13471_ _13472_ VGND VGND VPWR
+ VPWR _13473_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_47_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17457_ _13339_ _13403_ _13404_ _13405_ VGND VGND VPWR VPWR _13406_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14669_ _10709_ _10710_ execute.io_target_pc\[2\] _10711_ VGND VGND VPWR VPWR _10712_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_129_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16408_ _11260_ _12374_ _12375_ _12376_ VGND VGND VPWR VPWR _12377_ sky130_fd_sc_hd__a31o_1
XFILLER_0_171_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17388_ _13055_ net678 _13097_ VGND VGND VPWR VPWR _13338_ sky130_fd_sc_hd__o21a_1
XFILLER_0_171_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_164_clock clknet_5_25__leaf_clock VGND VGND VPWR VPWR clknet_leaf_164_clock
+ sky130_fd_sc_hd__clkbuf_8
X_19127_ decode.id_ex_aluop_reg\[1\] decode.id_ex_aluop_reg\[3\] decode.id_ex_aluop_reg\[2\]
+ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__or3b_4
X_16339_ _12133_ net463 _12274_ _12309_ _12132_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19058_ _04354_ _04355_ _04324_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18009_ decode.regfile.registers_27\[30\] _12507_ _12520_ _12967_ _03405_ VGND VGND
+ VPWR VPWR _03406_ sky130_fd_sc_hd__o311a_1
XFILLER_0_100_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_179_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_179_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21020_ _05994_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_203_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_102_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_102_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_203_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22971_ fetch.bht.bhtTable_target_pc\[0\]\[5\] fetch.bht.bhtTable_target_pc\[1\]\[5\]
+ fetch.bht.bhtTable_target_pc\[2\]\[5\] fetch.bht.bhtTable_target_pc\[3\]\[5\] _07098_
+ _07100_ VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__mux4_1
XFILLER_0_184_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24710_ _08072_ net1798 _08531_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21922_ net526 _06545_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25690_ _08914_ _09112_ VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_195_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_195_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24641_ _08503_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21853_ csr.io_mret_vector\[5\] _09884_ _06040_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_117_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_117_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27360_ clknet_leaf_328_clock _00389_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20804_ execute.io_mem_memtoreg\[1\] _05867_ _05875_ VGND VGND VPWR VPWR _05877_
+ sky130_fd_sc_hd__and3_1
X_24572_ net1598 execute.io_target_pc\[8\] _08462_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__mux2_1
X_21784_ _06455_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__clkbuf_1
X_26311_ _09443_ _09446_ VGND VGND VPWR VPWR _09488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_212_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23523_ _03546_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27291_ clknet_leaf_8_clock _00320_ VGND VGND VPWR VPWR decode.regfile.registers_31\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_20735_ _05831_ _05813_ net2563 _05838_ _00711_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29030_ clknet_leaf_97_clock _02043_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_154_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26242_ net689 _09447_ _09449_ _09440_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_154_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23454_ net6 _07861_ _07863_ _07851_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20666_ _05791_ _05792_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22405_ fetch.bht.bhtTable_tag\[4\]\[21\] fetch.bht.bhtTable_tag\[5\]\[21\] _06809_
+ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__mux2_1
X_26173_ _09400_ _09390_ VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__nand2_1
X_23385_ fetch.bht.bhtTable_target_pc\[0\]\[29\] fetch.bht.bhtTable_target_pc\[1\]\[29\]
+ fetch.bht.bhtTable_target_pc\[2\]\[29\] fetch.bht.bhtTable_target_pc\[3\]\[29\]
+ _07669_ _07100_ VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__mux4_1
X_20597_ csr._minstret_T_3\[54\] _05578_ _05617_ csr._csr_read_data_T_8\[22\] _05559_
+ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25124_ _08790_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_167_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22336_ _06684_ _06930_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_167_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25055_ _03555_ _08748_ csr.mcycle\[23\] VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__a21oi_1
X_29932_ clknet_leaf_340_clock _02945_ VGND VGND VPWR VPWR decode.regfile.registers_21\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_22267_ _06636_ _06855_ _06861_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_163_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24006_ _08174_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__clkbuf_1
X_21218_ _06104_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22198_ _06628_ _06789_ _06699_ _06792_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__o211a_1
X_29863_ clknet_leaf_298_clock _02876_ VGND VGND VPWR VPWR decode.regfile.registers_19\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28814_ clknet_leaf_109_clock _01827_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21149_ _06062_ _06058_ net786 VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__and3_1
X_29794_ clknet_leaf_309_clock _02807_ VGND VGND VPWR VPWR decode.regfile.registers_17\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28745_ clknet_leaf_95_clock _01758_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_25957_ _08954_ _09267_ VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__nand2_1
X_13971_ _09931_ decode.io_wb_rd\[0\] VGND VGND VPWR VPWR _10240_ sky130_fd_sc_hd__and2_4
X_15710_ decode.regfile.registers_2\[10\] _11369_ _11695_ _11696_ _11152_ VGND VGND
+ VPWR VPWR _11697_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_122_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24908_ net776 _08652_ _07179_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_122_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28676_ clknet_leaf_132_clock _01689_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16690_ _11019_ _12504_ _12650_ decode.regfile.registers_10\[0\] _12654_ VGND VGND
+ VPWR VPWR _12655_ sky130_fd_sc_hd__o32a_1
XFILLER_0_198_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25888_ net2516 _09226_ _09231_ _09222_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15641_ decode.regfile.registers_15\[8\] _11037_ _11205_ VGND VGND VPWR VPWR _11630_
+ sky130_fd_sc_hd__and3_1
X_24839_ _08387_ VGND VGND VPWR VPWR _08607_ sky130_fd_sc_hd__buf_4
X_27627_ clknet_leaf_43_clock net179 VGND VGND VPWR VPWR execute.io_reg_pc\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _03658_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__clkbuf_4
X_27558_ clknet_leaf_51_clock _00587_ VGND VGND VPWR VPWR execute.io_mem_isbranch
+ sky130_fd_sc_hd__dfxtp_1
X_15572_ _11050_ decode.regfile.registers_25\[6\] _11090_ VGND VGND VPWR VPWR _11563_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_90_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17311_ decode.regfile.registers_20\[13\] _11024_ _12553_ _12823_ _12537_ VGND VGND
+ VPWR VPWR _13263_ sky130_fd_sc_hd__a41o_1
X_14523_ fetch.bht.bhtTable_tag_MPORT_en fetch.btb.io_branch _10564_ _10567_ VGND
+ VGND VPWR VPWR _10568_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_25_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26509_ _09412_ _09602_ VGND VGND VPWR VPWR _09603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18291_ _03610_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27489_ clknet_leaf_33_clock _00518_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_81_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_81_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17242_ decode.regfile.registers_7\[11\] _12611_ _12623_ decode.regfile.registers_6\[11\]
+ VGND VGND VPWR VPWR _13196_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_83_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29228_ clknet_leaf_117_clock _02241_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14454_ _10031_ _10517_ VGND VGND VPWR VPWR _10521_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_96_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29159_ clknet_leaf_196_clock _02172_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17173_ _10927_ decode.regfile.registers_24\[9\] _10933_ _12759_ _11026_ VGND VGND
+ VPWR VPWR _13129_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_25_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14385_ net592 _10477_ _10480_ _10481_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16124_ _11493_ decode.regfile.registers_22\[21\] _11450_ _10979_ _10991_ VGND VGND
+ VPWR VPWR _12100_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_52_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_96_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_96_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16055_ decode.regfile.registers_11\[19\] _11071_ _11470_ _11278_ VGND VGND VPWR
+ VPWR _12033_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_55_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15006_ decode.immGen._imm_T_24\[19\] VGND VGND VPWR VPWR _11016_ sky130_fd_sc_hd__buf_2
XFILLER_0_209_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19814_ _03705_ _04509_ _04332_ _04412_ _04700_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__a41o_1
Xhold1709 csr.mscratch\[11\] VGND VGND VPWR VPWR net1936 sky130_fd_sc_hd__dlygate4sd3_1
X_19745_ _05016_ _05018_ _03851_ _04525_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__a31o_1
X_16957_ _12695_ _12914_ _12916_ _12917_ VGND VGND VPWR VPWR _12918_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15908_ decode.regfile.registers_8\[15\] _11045_ _11175_ VGND VGND VPWR VPWR _11890_
+ sky130_fd_sc_hd__a21o_1
X_19676_ _03947_ _03944_ _04503_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_34_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_34_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16888_ decode.regfile.registers_11\[3\] _12594_ _12582_ _12550_ _12849_ VGND VGND
+ VPWR VPWR _12850_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18627_ _03659_ execute.csr_read_data_out_reg\[16\] execute.io_reg_pc\[16\] _03777_
+ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__o22a_1
X_15839_ decode.regfile.registers_21\[13\] _11267_ _11099_ _11228_ _11822_ VGND VGND
+ VPWR VPWR _11823_ sky130_fd_sc_hd__o311a_1
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18558_ memory.csr_read_data_out_reg\[30\] _09988_ _10140_ VGND VGND VPWR VPWR _03857_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_190_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_190_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17509_ decode.regfile.registers_1\[18\] _12778_ _12830_ _12882_ _13455_ VGND VGND
+ VPWR VPWR _13456_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_49_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_49_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_16_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18489_ _03709_ decode.id_ex_imm_reg\[29\] _03787_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_16_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_13 _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20520_ csr.mcycle\[11\] _05552_ _05604_ net33 _05668_ VGND VGND VPWR VPWR _05669_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_24 _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _10019_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_46 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_57 _10657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20451_ csr.msie _05517_ _05527_ _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_68 _11036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_79 _11215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23170_ fetch.bht.bhtTable_target_pc\[8\]\[16\] fetch.bht.bhtTable_target_pc\[9\]\[16\]
+ _07099_ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__mux2_1
X_20382_ _05539_ _05542_ _05543_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22121_ _06632_ _06711_ _06713_ _06715_ _06699_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_3_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput120 net120 VGND VGND VPWR VPWR io_memory_address[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput131 net131 VGND VGND VPWR VPWR io_memory_address[9] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput142 net142 VGND VGND VPWR VPWR io_memory_write_data[15] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22052_ fetch.bht.bhtTable_tag\[4\]\[22\] fetch.bht.bhtTable_tag\[5\]\[22\] _06646_
+ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_205_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput153 net153 VGND VGND VPWR VPWR io_memory_write_data[25] sky130_fd_sc_hd__clkbuf_4
Xoutput164 net164 VGND VGND VPWR VPWR io_memory_write_data[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_220_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21003_ _03582_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__clkbuf_2
X_26860_ _09387_ _09796_ VGND VGND VPWR VPWR _09805_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_4 _00707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_197_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_197_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25811_ net2081 _09183_ _09187_ _09182_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26791_ net1954 _09752_ _09765_ _09758_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28530_ clknet_leaf_218_clock _01543_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_25742_ net2123 _09139_ _09147_ _09142_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__o211a_1
X_22954_ _07401_ _07402_ _07082_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28461_ clknet_leaf_137_clock _01474_ VGND VGND VPWR VPWR decode.io_id_pc\[19\] sky130_fd_sc_hd__dfxtp_1
X_21905_ _03449_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__buf_2
XFILLER_0_223_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25673_ _08973_ _09067_ VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__nand2_1
X_22885_ _07339_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27412_ clknet_leaf_10_clock _00441_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[21\]
+ sky130_fd_sc_hd__dfxtp_4
X_24624_ _08494_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__clkbuf_1
X_28392_ clknet_leaf_58_clock _01405_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_156_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21836_ _03449_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27343_ clknet_leaf_44_clock _00372_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_24555_ net1395 execute.io_target_pc\[0\] _07335_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21767_ _06446_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23506_ net2213 _07890_ _07887_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__or3b_1
X_27274_ clknet_leaf_13_clock _00303_ VGND VGND VPWR VPWR decode.regfile.registers_30\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_20718_ decode.id_ex_rs1_data_reg\[18\] VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__inv_2
X_24486_ _08423_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21698_ csr.minstret\[22\] csr.minstret\[23\] csr.minstret\[24\] VGND VGND VPWR VPWR
+ _06400_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29013_ clknet_leaf_115_clock _02026_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26225_ _09436_ _09372_ VGND VGND VPWR VPWR _09437_ sky130_fd_sc_hd__nand2_1
X_23437_ net30 _07846_ _07853_ _07851_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20649_ net2699 _05588_ _05778_ _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14170_ _10290_ VGND VGND VPWR VPWR _10357_ sky130_fd_sc_hd__buf_2
X_26156_ net748 _09373_ _09388_ _09370_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__o211a_1
X_23368_ fetch.bht.bhtTable_target_pc\[13\]\[28\] _07099_ VGND VGND VPWR VPWR _07793_
+ sky130_fd_sc_hd__or2b_1
X_25107_ _06124_ net2049 _08778_ VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22319_ net227 _06907_ _06913_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26087_ _08933_ _09340_ VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__nand2_1
X_23299_ net223 net80 net79 _07651_ net222 VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__a41o_1
XFILLER_0_104_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25038_ csr._mcycle_T_2\[17\] _08710_ _08738_ csr.mcycle\[17\] VGND VGND VPWR VPWR
+ _08739_ sky130_fd_sc_hd__a211oi_1
X_29915_ clknet_leaf_304_clock _02928_ VGND VGND VPWR VPWR decode.regfile.registers_21\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29846_ clknet_leaf_299_clock _02859_ VGND VGND VPWR VPWR decode.regfile.registers_18\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_17860_ _12967_ _03258_ _03259_ _03260_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16811_ _12582_ _10603_ _10617_ VGND VGND VPWR VPWR _12774_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_145_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17791_ decode.regfile.registers_2\[25\] _12634_ _12629_ _03192_ VGND VGND VPWR VPWR
+ _03193_ sky130_fd_sc_hd__o211ai_2
X_29777_ clknet_leaf_294_clock _02790_ VGND VGND VPWR VPWR decode.regfile.registers_16\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26989_ _10146_ _09838_ VGND VGND VPWR VPWR _09878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19530_ _04249_ _04812_ _04813_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__o21ai_1
X_28728_ clknet_leaf_121_clock _01741_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_13954_ _10107_ _10223_ VGND VGND VPWR VPWR _10231_ sky130_fd_sc_hd__nand2_1
X_16742_ _12667_ VGND VGND VPWR VPWR _12706_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_85_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16673_ _11016_ _10597_ decode.immGen._imm_T_24\[17\] _12637_ VGND VGND VPWR VPWR
+ _12638_ sky130_fd_sc_hd__nor4_1
X_19461_ _04115_ _04442_ _04444_ net264 VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__o211a_1
X_28659_ clknet_leaf_140_clock _01672_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_13885_ _10128_ _10152_ VGND VGND VPWR VPWR _10190_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18412_ execute.io_mem_rd\[1\] net297 VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_203 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15624_ decode.regfile.registers_17\[8\] _11128_ _11106_ VGND VGND VPWR VPWR _11613_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_202_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19392_ _04415_ _04669_ _04676_ _04681_ _03595_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__o311a_2
XTAP_TAPCELL_ROW_48_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_214 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_225 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_202_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_236 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_247 net193 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15555_ _10635_ _11143_ net319 VGND VGND VPWR VPWR _11546_ sky130_fd_sc_hd__and3_1
X_18343_ execute.io_mem_rd\[0\] VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__inv_2
XINSDIODE1_258 clknet_0_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_269 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ fetch.btb.btbTable\[12\]\[1\] fetch.btb.btbTable\[13\]\[1\] fetch.btb.btbTable\[14\]\[1\]
+ fetch.btb.btbTable\[15\]\[1\] _09891_ _09888_ VGND VGND VPWR VPWR _10551_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_44_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18274_ _03601_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__clkbuf_1
X_15486_ decode.regfile.registers_19\[4\] _11453_ _11454_ _11478_ VGND VGND VPWR VPWR
+ _11479_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17225_ _13099_ _12768_ _12493_ decode.regfile.registers_29\[10\] _13179_ VGND VGND
+ VPWR VPWR _13180_ sky130_fd_sc_hd__o221a_1
X_14437_ net801 _10506_ _10511_ _10509_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput11 io_fetch_data[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 net385 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput33 io_meip VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput44 io_memory_read_data[19] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_1
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17156_ _11018_ _12977_ _12510_ decode.regfile.registers_9\[9\] VGND VGND VPWR VPWR
+ _13112_ sky130_fd_sc_hd__or4b_1
XFILLER_0_226_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput55 io_memory_read_data[29] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14368_ net661 _10463_ _10471_ _10468_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__o211a_1
Xinput66 reset VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold806 decode.regfile.registers_27\[8\] VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold817 fetch.bht.bhtTable_target_pc\[15\]\[16\] VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ _10957_ _11217_ _11085_ decode.regfile.registers_21\[20\] _11648_ VGND VGND
+ VPWR VPWR _12084_ sky130_fd_sc_hd__o32a_1
XFILLER_0_40_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold828 fetch.bht.bhtTable_tag\[1\]\[25\] VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17087_ _12505_ VGND VGND VPWR VPWR _13045_ sky130_fd_sc_hd__buf_2
Xhold839 decode.regfile.registers_27\[25\] VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14299_ _10015_ _10431_ VGND VGND VPWR VPWR _10432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_228_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16038_ _11263_ decode.regfile.registers_22\[19\] _11404_ _11264_ _11265_ VGND VGND
+ VPWR VPWR _12016_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_20_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2207 decode.regfile.registers_1\[7\] VGND VGND VPWR VPWR net2434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2218 _01130_ VGND VGND VPWR VPWR net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2229 decode.regfile.registers_25\[22\] VGND VGND VPWR VPWR net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1506 csr._mcycle_T_2\[8\] VGND VGND VPWR VPWR net1733 sky130_fd_sc_hd__clkbuf_2
Xhold1517 fetch.bht.bhtTable_tag\[14\]\[20\] VGND VGND VPWR VPWR net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1528 decode.regfile.registers_20\[20\] VGND VGND VPWR VPWR net1755 sky130_fd_sc_hd__dlygate4sd3_1
X_17989_ decode.regfile.registers_7\[30\] _12610_ _12737_ decode.regfile.registers_6\[30\]
+ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__a221oi_2
Xhold1539 fetch.bht.bhtTable_target_pc\[2\]\[16\] VGND VGND VPWR VPWR net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19728_ _04465_ _04997_ _05001_ _05002_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__a41o_2
XTAP_TAPCELL_ROW_192_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_192_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19659_ _03957_ _03960_ _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_205_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22670_ net2765 _07208_ _07220_ _07221_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21621_ csr.minstret\[6\] _06342_ csr.minstret\[7\] VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24340_ _08346_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21552_ _06296_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20503_ csr.mcycle\[9\] _05587_ _05594_ csr.minstret\[9\] VGND VGND VPWR VPWR _05654_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24271_ _08099_ net1070 _06218_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21483_ _06258_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26010_ net683 _09300_ _09302_ _09292_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23222_ _07070_ VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__buf_4
X_20434_ _05591_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23153_ net280 _07589_ _07590_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__and3_1
XFILLER_0_160_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20365_ _05527_ _03755_ _03737_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__and3_2
XFILLER_0_28_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_228_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22104_ _06640_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_149_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27961_ clknet_leaf_184_clock _00983_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_23084_ _07525_ _07406_ _07097_ VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_149_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20296_ _10806_ decode.id_ex_pc_reg\[18\] _05468_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__and3_2
XFILLER_0_41_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29700_ clknet_leaf_281_clock _02713_ VGND VGND VPWR VPWR decode.regfile.registers_14\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_224_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22035_ _06625_ _06629_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_181_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26912_ _09441_ _09794_ VGND VGND VPWR VPWR _09834_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_181_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27892_ clknet_leaf_19_clock _00921_ VGND VGND VPWR VPWR csr._mcycle_T_2\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29631_ clknet_leaf_271_clock _02644_ VGND VGND VPWR VPWR decode.regfile.registers_12\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_26843_ _09794_ VGND VGND VPWR VPWR _09795_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_215_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26774_ _09377_ _09753_ VGND VGND VPWR VPWR _09756_ sky130_fd_sc_hd__nand2_1
X_29562_ clknet_leaf_312_clock _02575_ VGND VGND VPWR VPWR decode.regfile.registers_10\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_23986_ _07959_ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__buf_4
XFILLER_0_215_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28513_ clknet_leaf_210_clock _01526_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_25725_ _08948_ _09136_ VGND VGND VPWR VPWR _09138_ sky130_fd_sc_hd__nand2_1
X_22937_ fetch.bht.bhtTable_target_pc\[8\]\[3\] fetch.bht.bhtTable_target_pc\[9\]\[3\]
+ fetch.bht.bhtTable_target_pc\[10\]\[3\] fetch.bht.bhtTable_target_pc\[11\]\[3\]
+ _07106_ _07386_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29493_ clknet_leaf_264_clock _02506_ VGND VGND VPWR VPWR decode.regfile.registers_7\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_179_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28444_ clknet_leaf_55_clock _01457_ VGND VGND VPWR VPWR decode.io_id_pc\[2\] sky130_fd_sc_hd__dfxtp_1
X_25656_ _08956_ _09092_ VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__nand2_1
X_13670_ _10025_ _10016_ VGND VGND VPWR VPWR _10026_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22868_ _07330_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24607_ net1818 execute.io_target_pc\[25\] _09897_ VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28375_ clknet_leaf_186_clock _01388_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21819_ _06480_ csr._csr_read_data_T_9\[31\] _06482_ VGND VGND VPWR VPWR _06483_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25587_ _08962_ _09049_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22799_ _07294_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15340_ _11335_ VGND VGND VPWR VPWR _11336_ sky130_fd_sc_hd__clkbuf_4
X_27326_ clknet_leaf_25_clock _00355_ VGND VGND VPWR VPWR decode.id_ex_funct3_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24538_ _08450_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_117_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15271_ _11060_ VGND VGND VPWR VPWR _11267_ sky130_fd_sc_hd__buf_2
X_27257_ clknet_leaf_9_clock _00286_ VGND VGND VPWR VPWR decode.regfile.registers_30\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_24469_ _08414_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17010_ decode.regfile.registers_2\[6\] _12835_ _12836_ decode.regfile.registers_3\[6\]
+ _12838_ VGND VGND VPWR VPWR _12969_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_108_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26208_ net2519 _09419_ _09425_ _09418_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__o211a_1
X_14222_ _10375_ VGND VGND VPWR VPWR _10387_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27188_ clknet_leaf_6_clock _00217_ VGND VGND VPWR VPWR decode.regfile.registers_28\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14153_ net2244 _10346_ _10347_ _10344_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__o211a_1
X_26139_ _09969_ VGND VGND VPWR VPWR _09377_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14084_ net2179 _10302_ _10307_ _10304_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__o211a_1
X_18961_ _03888_ _03872_ _04233_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17912_ _03308_ _03310_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18892_ _03948_ _03962_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_119_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17843_ _03242_ _12659_ _12664_ _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__a211o_1
X_29829_ clknet_leaf_303_clock _02842_ VGND VGND VPWR VPWR decode.regfile.registers_18\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17774_ _13339_ _03174_ _03175_ _03176_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__a31o_1
XFILLER_0_221_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14986_ _11001_ _11003_ _10974_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19513_ _04270_ _04332_ _03704_ _04291_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__o211a_1
X_16725_ _12604_ VGND VGND VPWR VPWR _12690_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13937_ net1577 _10213_ _10221_ _10219_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_18_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19444_ _04727_ _04729_ _04730_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_46_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13868_ _10087_ _10177_ VGND VGND VPWR VPWR _10181_ sky130_fd_sc_hd__nand2_1
X_16656_ _10607_ _12522_ _12597_ VGND VGND VPWR VPWR _12621_ sky130_fd_sc_hd__and3_1
XFILLER_0_186_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15607_ _11269_ _11595_ _11596_ VGND VGND VPWR VPWR _11597_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19375_ _04143_ _04664_ _04142_ _04496_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__o31a_1
X_16587_ _12551_ VGND VGND VPWR VPWR _12552_ sky130_fd_sc_hd__clkbuf_4
X_13799_ memory.csr_read_data_out_reg\[29\] _09988_ _10134_ VGND VGND VPWR VPWR _10135_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_186_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18326_ decode.id_ex_rs2_data_reg\[28\] _03627_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15538_ _11493_ decode.regfile.registers_24\[6\] VGND VGND VPWR VPWR _11529_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15469_ _11082_ VGND VGND VPWR VPWR _11462_ sky130_fd_sc_hd__clkbuf_4
X_18257_ _03581_ _03583_ net531 VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__and3b_1
XFILLER_0_163_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17208_ decode.regfile.registers_19\[10\] _12679_ _12545_ _13162_ VGND VGND VPWR
+ VPWR _13163_ sky130_fd_sc_hd__o211a_1
X_18188_ _10579_ _10578_ decode.control.io_opcode\[5\] decode.control.io_opcode\[4\]
+ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__or4b_1
XFILLER_0_4_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold603 csr.mscratch\[0\] VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold614 fetch.bht.bhtTable_tag\[8\]\[4\] VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17139_ _12765_ _12768_ _12493_ decode.regfile.registers_29\[8\] _13095_ VGND VGND
+ VPWR VPWR _13096_ sky130_fd_sc_hd__o221a_1
Xhold625 fetch.bht.bhtTable_target_pc\[4\]\[13\] VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold636 fetch.bht.bhtTable_target_pc\[4\]\[26\] VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 decode.regfile.registers_28\[27\] VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _01229_ VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__dlygate4sd3_1
X_20150_ _05222_ _05355_ _05228_ _00569_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold669 decode.regfile.registers_20\[3\] VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20081_ decode.id_ex_imm_reg\[12\] decode.id_ex_pc_reg\[12\] VGND VGND VPWR VPWR
+ _05296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2004 fetch.bht.bhtTable_target_pc\[10\]\[4\] VGND VGND VPWR VPWR net2231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2015 decode.regfile.registers_28\[12\] VGND VGND VPWR VPWR net2242 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2026 decode.regfile.registers_15\[5\] VGND VGND VPWR VPWR net2253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2037 decode.regfile.registers_12\[13\] VGND VGND VPWR VPWR net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1303 fetch.bht.bhtTable_tag\[2\]\[22\] VGND VGND VPWR VPWR net1530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2048 decode.regfile.registers_10\[12\] VGND VGND VPWR VPWR net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1314 fetch.bht.bhtTable_target_pc\[13\]\[28\] VGND VGND VPWR VPWR net1541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2059 decode.regfile.registers_25\[7\] VGND VGND VPWR VPWR net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 fetch.bht.bhtTable_tag\[15\]\[5\] VGND VGND VPWR VPWR net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1336 fetch.bht.bhtTable_tag\[15\]\[1\] VGND VGND VPWR VPWR net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_227_Right_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23840_ execute.io_target_pc\[15\] VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__buf_2
XFILLER_0_139_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1347 fetch.bht.bhtTable_target_pc\[9\]\[1\] VGND VGND VPWR VPWR net1574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1358 fetch.bht.bhtTable_target_pc\[10\]\[2\] VGND VGND VPWR VPWR net1585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1369 fetch.bht.bhtTable_tag\[2\]\[17\] VGND VGND VPWR VPWR net1596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23771_ _08037_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__clkbuf_1
X_20983_ _05974_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25510_ net2628 _09008_ _09013_ _09004_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__o211a_1
X_22722_ _10946_ _03520_ _07252_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__o21ai_1
X_26490_ _09577_ VGND VGND VPWR VPWR _09592_ sky130_fd_sc_hd__buf_2
XFILLER_0_36_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25441_ _06578_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22653_ csr._csr_read_data_T_8\[3\] _07208_ _07212_ _07164_ VGND VGND VPWR VPWR _01287_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28160_ clknet_leaf_64_clock _01182_ VGND VGND VPWR VPWR csr.pie sky130_fd_sc_hd__dfxtp_1
X_21604_ _03579_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__buf_4
XFILLER_0_192_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25372_ _08922_ _08923_ VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22584_ _06377_ _07165_ _07166_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__nor3_1
XFILLER_0_192_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27111_ clknet_leaf_348_clock _00140_ VGND VGND VPWR VPWR decode.regfile.registers_25\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24323_ _08085_ net1721 _08334_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28091_ clknet_leaf_185_clock _01113_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21535_ _06287_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27042_ clknet_leaf_342_clock _00071_ VGND VGND VPWR VPWR decode.regfile.registers_23\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24254_ _08302_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__clkbuf_1
X_21466_ _05246_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23205_ _07638_ _07639_ _06633_ VGND VGND VPWR VPWR _07640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20417_ _05574_ _05575_ csr.minstret\[1\] VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24185_ _08078_ net1372 _08266_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__mux2_1
X_21397_ _06145_ net1975 _06210_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23136_ fetch.bht.bhtTable_target_pc\[4\]\[14\] fetch.bht.bhtTable_target_pc\[5\]\[14\]
+ fetch.bht.bhtTable_target_pc\[6\]\[14\] fetch.bht.bhtTable_target_pc\[7\]\[14\]
+ _07099_ _07103_ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__mux4_1
XFILLER_0_219_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20348_ _05406_ _05418_ _03517_ _03551_ _05512_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__a2111oi_1
X_28993_ clknet_leaf_169_clock _02006_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23067_ _07125_ _07509_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__and2b_1
X_27944_ clknet_leaf_207_clock _00966_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20279_ _05417_ _05307_ _05460_ _05454_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22018_ net1809 _06573_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__or2_1
X_27875_ clknet_leaf_67_clock _00904_ VGND VGND VPWR VPWR csr.io_interrupt sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2560 decode.regfile.registers_30\[14\] VGND VGND VPWR VPWR net2787 sky130_fd_sc_hd__dlygate4sd3_1
X_29614_ clknet_leaf_279_clock _02627_ VGND VGND VPWR VPWR decode.regfile.registers_11\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14840_ _10813_ _10882_ _10721_ VGND VGND VPWR VPWR _10883_ sky130_fd_sc_hd__a21o_1
Xhold2571 csr._mcycle_T_2\[18\] VGND VGND VPWR VPWR net2798 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_106_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26826_ net2451 _09779_ _09785_ _09784_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_106_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1870 execute.csr_write_data_out_reg\[17\] VGND VGND VPWR VPWR net2097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1881 fetch.bht.bhtTable_target_pc\[12\]\[4\] VGND VGND VPWR VPWR net2108 sky130_fd_sc_hd__dlygate4sd3_1
X_14771_ _10812_ _10813_ VGND VGND VPWR VPWR _10814_ sky130_fd_sc_hd__xor2_1
X_29545_ clknet_leaf_273_clock _02558_ VGND VGND VPWR VPWR decode.regfile.registers_9\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_23969_ _08155_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_177_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26757_ net2363 _09736_ _09745_ _09743_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1892 fetch.bht.bhtTable_tag\[15\]\[4\] VGND VGND VPWR VPWR net2119 sky130_fd_sc_hd__dlygate4sd3_1
X_13722_ _10069_ _10016_ VGND VGND VPWR VPWR _10070_ sky130_fd_sc_hd__nand2_1
X_16510_ decode.regfile.registers_20\[31\] _11102_ _11327_ _12475_ VGND VGND VPWR
+ VPWR _12476_ sky130_fd_sc_hd__a211o_1
X_25708_ _09128_ VGND VGND VPWR VPWR _09129_ sky130_fd_sc_hd__buf_2
XFILLER_0_169_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17490_ decode.regfile.registers_17\[17\] _12719_ _12565_ _13437_ VGND VGND VPWR
+ VPWR _13438_ sky130_fd_sc_hd__o211a_1
X_26688_ net2409 _09666_ _09705_ _09702_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__o211a_1
X_29476_ clknet_leaf_263_clock _02489_ VGND VGND VPWR VPWR decode.regfile.registers_7\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28427_ clknet_leaf_247_clock _01440_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[17\]
+ sky130_fd_sc_hd__dfxtp_4
X_16441_ decode.regfile.registers_21\[29\] _11061_ _11100_ _11229_ _12408_ VGND VGND
+ VPWR VPWR _12409_ sky130_fd_sc_hd__o311a_1
X_13653_ _09942_ VGND VGND VPWR VPWR _10010_ sky130_fd_sc_hd__buf_4
X_25639_ net2759 _09082_ _09088_ _09087_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19160_ _04450_ _04453_ _04454_ _04456_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__a2bb2o_1
X_16372_ _11076_ decode.regfile.registers_27\[27\] _11869_ VGND VGND VPWR VPWR _12342_
+ sky130_fd_sc_hd__or3_1
X_28358_ clknet_leaf_216_clock _01371_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13584_ memory.csr_read_data_out_reg\[0\] _09942_ _09945_ _09948_ VGND VGND VPWR
+ VPWR _09949_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_27_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18111_ _03482_ _03480_ _03474_ net2200 VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15323_ _11279_ _11317_ _11318_ _11053_ VGND VGND VPWR VPWR _11319_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_136_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27309_ clknet_leaf_9_clock _00338_ VGND VGND VPWR VPWR decode.regfile.registers_31\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19091_ _04246_ _04373_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__nand2_1
X_28289_ clknet_leaf_86_clock _01311_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15254_ _11050_ VGND VGND VPWR VPWR _11250_ sky130_fd_sc_hd__clkbuf_4
X_18042_ _12712_ decode.regfile.registers_24\[31\] _12997_ _12998_ _11025_ VGND VGND
+ VPWR VPWR _03438_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_83_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14205_ _09950_ _10377_ VGND VGND VPWR VPWR _10378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15185_ _10628_ net324 _11042_ _11057_ VGND VGND VPWR VPWR _11182_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14136_ net494 _10332_ _10337_ _10328_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__o211a_1
X_19993_ _10684_ _05219_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18944_ _04028_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__buf_2
X_14067_ net855 _10287_ _10297_ _10291_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18875_ _04171_ _04172_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_197_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17826_ decode.regfile.registers_18\[26\] _12572_ _12562_ VGND VGND VPWR VPWR _03227_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17757_ decode.regfile.registers_8\[24\] _12726_ _03152_ _03159_ VGND VGND VPWR VPWR
+ _03160_ sky130_fd_sc_hd__o22a_1
X_14969_ _10993_ VGND VGND VPWR VPWR _10994_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_222_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16708_ _12672_ VGND VGND VPWR VPWR _12673_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17688_ _12650_ _12723_ _12669_ decode.regfile.registers_14\[22\] _03092_ VGND VGND
+ VPWR VPWR _03093_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19427_ _04155_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16639_ _12592_ VGND VGND VPWR VPWR _12604_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19358_ _04648_ _04548_ _04270_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18309_ decode.id_ex_rs2_data_reg\[20\] _03616_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__and2_1
X_19289_ _04050_ _04559_ _04051_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__o21bai_4
XTAP_TAPCELL_ROW_212_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_212_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21320_ _06170_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21251_ net1385 _06126_ _06120_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold400 decode.regfile.registers_24\[12\] VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 execute.csr_write_address_out_reg\[2\] VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 decode.regfile.registers_21\[14\] VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20202_ decode.id_ex_imm_reg\[29\] _10697_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__and2_1
Xhold433 decode.regfile.registers_27\[11\] VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold444 decode.regfile.registers_29\[12\] VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__dlygate4sd3_1
X_21182_ _05866_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__buf_2
Xhold455 decode.regfile.registers_4\[10\] VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold466 decode.regfile.registers_6\[0\] VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 fetch.bht.bhtTable_valid\[9\] VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap196 _10116_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_4
X_20133_ decode.id_ex_imm_reg\[19\] _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__or2_1
Xhold488 decode.regfile.registers_18\[16\] VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_221_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold499 decode.regfile.registers_24\[6\] VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__dlygate4sd3_1
X_25990_ _08912_ _09287_ VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20064_ _05281_ _05239_ _00557_ _05227_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__o22a_1
X_24941_ csr._mcycle_T_3\[48\] csr._mcycle_T_3\[47\] _08670_ VGND VGND VPWR VPWR _08674_
+ sky130_fd_sc_hd__and3_1
Xhold1100 fetch.bht.bhtTable_tag\[1\]\[5\] VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1111 fetch.bht.bhtTable_target_pc\[5\]\[20\] VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 fetch.bht.bhtTable_tag\[3\]\[15\] VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__dlygate4sd3_1
X_24872_ _06151_ net2076 _08388_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__mux2_1
Xhold1133 decode.regfile.registers_17\[3\] VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__dlygate4sd3_1
X_27660_ clknet_leaf_26_clock _00689_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1144 fetch.bht.bhtTable_target_pc\[6\]\[6\] VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 fetch.bht.bhtTable_target_pc\[12\]\[15\] VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1166 fetch.bht.bhtTable_tag\[6\]\[12\] VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__dlygate4sd3_1
X_23823_ _08069_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26611_ _09441_ _09621_ VGND VGND VPWR VPWR _09661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_213_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27591_ clknet_leaf_146_clock _00620_ VGND VGND VPWR VPWR execute.io_target_pc\[0\]
+ sky130_fd_sc_hd__dfxtp_4
Xhold1177 execute.csr_write_data_out_reg\[13\] VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1188 fetch.bht.bhtTable_target_pc\[0\]\[17\] VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 fetch.bht.bhtTable_target_pc\[7\]\[9\] VGND VGND VPWR VPWR net1426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_219_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29330_ clknet_leaf_226_clock _02343_ VGND VGND VPWR VPWR decode.regfile.registers_2\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_26542_ _09621_ VGND VGND VPWR VPWR _09622_ sky130_fd_sc_hd__clkbuf_4
X_23754_ _08028_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20966_ _05866_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22705_ net2684 _07235_ _07241_ _07234_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29261_ clknet_leaf_232_clock _02274_ VGND VGND VPWR VPWR decode.regfile.registers_0\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_1322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26473_ _09377_ _09579_ VGND VGND VPWR VPWR _09583_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_172_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23685_ net1556 _10820_ _07992_ VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__mux2_1
X_20897_ _05925_ _05921_ net65 VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__and3_1
XFILLER_0_222_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28212_ clknet_leaf_60_clock net807 VGND VGND VPWR VPWR csr.mscratch\[14\] sky130_fd_sc_hd__dfxtp_1
X_25424_ net197 VGND VGND VPWR VPWR _08960_ sky130_fd_sc_hd__buf_4
X_22636_ csr._minstret_T_3\[60\] csr._minstret_T_3\[59\] csr._minstret_T_3\[58\] _07196_
+ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__and4_1
X_29192_ clknet_leaf_239_clock _02205_ VGND VGND VPWR VPWR fetch.btb.btbTable\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_0__f_clock clknet_2_0_0_clock VGND VGND VPWR VPWR clknet_5_0__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28143_ clknet_leaf_193_clock _01165_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_25355_ net210 VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__buf_4
X_22567_ _06417_ _07140_ _07152_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24306_ _08068_ net1426 _08323_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21518_ _06147_ net2040 _06274_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__mux2_1
X_28074_ clknet_leaf_238_clock _01096_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25286_ _08873_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22498_ _07086_ _07089_ _07092_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_131_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27025_ clknet_leaf_333_clock _00054_ VGND VGND VPWR VPWR decode.regfile.registers_23\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24237_ _08293_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21449_ _06140_ net2036 _06230_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24168_ _08062_ net1534 _08255_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23119_ _07082_ _07558_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__nor2_1
X_28976_ clknet_leaf_105_clock _01989_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24099_ _08222_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__clkbuf_1
X_16990_ _11022_ _12568_ _12535_ _12949_ VGND VGND VPWR VPWR _12950_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_34_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27927_ clknet_leaf_33_clock _00956_ VGND VGND VPWR VPWR execute.io_mem_rd\[3\] sky130_fd_sc_hd__dfxtp_2
X_15941_ _11289_ _11920_ _11921_ VGND VGND VPWR VPWR _11922_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_129_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _03953_ _03954_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__nand2_4
X_15872_ decode.regfile.registers_12\[14\] _11194_ _11839_ _11854_ VGND VGND VPWR
+ VPWR _11855_ sky130_fd_sc_hd__o22ai_1
X_27858_ clknet_leaf_318_clock _00887_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2390 csr._minstret_T_3\[42\] VGND VGND VPWR VPWR net2617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17611_ decode.regfile.registers_19\[20\] _12678_ _02998_ _03017_ _12544_ VGND VGND
+ VPWR VPWR _03018_ sky130_fd_sc_hd__o221a_1
XFILLER_0_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14823_ _10796_ _10865_ VGND VGND VPWR VPWR _10866_ sky130_fd_sc_hd__or2_1
X_26809_ net1723 _09766_ _09775_ _09771_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18591_ _03889_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__buf_6
XFILLER_0_203_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27789_ clknet_leaf_333_clock _00818_ VGND VGND VPWR VPWR memory.io_wb_readdata\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17542_ _13215_ decode.regfile.registers_28\[18\] _13093_ VGND VGND VPWR VPWR _13489_
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_48_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29528_ clknet_leaf_314_clock _02541_ VGND VGND VPWR VPWR decode.regfile.registers_8\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14754_ csr.io_mem_pc\[21\] _10796_ VGND VGND VPWR VPWR _10797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13705_ memory.io_wb_readdata\[15\] _09981_ VGND VGND VPWR VPWR _10055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14685_ _10678_ execute.io_target_pc\[6\] VGND VGND VPWR VPWR _10728_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_138_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17473_ decode.regfile.registers_7\[17\] _12882_ _13020_ _12622_ decode.regfile.registers_6\[17\]
+ VGND VGND VPWR VPWR _13421_ sky130_fd_sc_hd__a32o_1
X_29459_ clknet_leaf_261_clock _02472_ VGND VGND VPWR VPWR decode.regfile.registers_6\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19212_ _04345_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__clkbuf_4
X_16424_ _12386_ _12390_ _12391_ VGND VGND VPWR VPWR _12392_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_28_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13636_ _09977_ VGND VGND VPWR VPWR _09995_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_172_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19143_ _04305_ _04430_ _04437_ _04439_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__o211a_1
X_16355_ decode.regfile.registers_9\[27\] _11547_ _12323_ _12324_ _11509_ VGND VGND
+ VPWR VPWR _12325_ sky130_fd_sc_hd__a221o_1
X_13567_ decode.io_wb_rd\[0\] _09931_ VGND VGND VPWR VPWR _09932_ sky130_fd_sc_hd__nor2_4
XFILLER_0_137_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15306_ _11298_ _10646_ _11299_ _11301_ VGND VGND VPWR VPWR _11302_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16286_ _12257_ decode.regfile.registers_17\[25\] _11356_ VGND VGND VPWR VPWR _12258_
+ sky130_fd_sc_hd__mux2_1
X_19074_ _04062_ _04126_ _04045_ _04070_ _04320_ _04325_ VGND VGND VPWR VPWR _04372_
+ sky130_fd_sc_hd__mux4_2
X_13498_ _09879_ VGND VGND VPWR VPWR _09880_ sky130_fd_sc_hd__buf_2
XFILLER_0_152_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18025_ decode.regfile.registers_9\[31\] _12498_ _12977_ _12510_ _12653_ VGND VGND
+ VPWR VPWR _03421_ sky130_fd_sc_hd__o41a_1
X_15237_ _11088_ decode.regfile.registers_23\[0\] _11090_ _11233_ VGND VGND VPWR VPWR
+ _11234_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_57_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15168_ _11164_ VGND VGND VPWR VPWR _11165_ sky130_fd_sc_hd__buf_2
XFILLER_0_67_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14119_ net2593 _10315_ _10326_ _10317_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_58_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19976_ net428 _05217_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15099_ _11095_ VGND VGND VPWR VPWR _11096_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18927_ _04075_ _04172_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_207_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18858_ _03658_ execute.csr_read_data_out_reg\[10\] execute.io_reg_pc\[10\] _03776_
+ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17809_ _12562_ _03210_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_66_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_1056 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18789_ _03658_ execute.csr_read_data_out_reg\[15\] execute.io_reg_pc\[15\] _03776_
+ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__o22a_1
XFILLER_0_179_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20820_ _05885_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20751_ _03737_ _05671_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_214_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23470_ _10657_ _07862_ _07859_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20682_ decode.id_ex_rs1_data_reg\[4\] decode.id_ex_ex_rs1_reg\[4\] _05056_ VGND
+ VGND VPWR VPWR _05806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22421_ _06628_ _07011_ _06635_ _07015_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_134_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_210_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25140_ _10946_ _10944_ _00461_ _08799_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22352_ fetch.bht.bhtTable_tag\[4\]\[14\] fetch.bht.bhtTable_tag\[5\]\[14\] net277
+ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_332_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_332_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21303_ _06161_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25071_ csr.mcycle\[26\] csr.mcycle\[25\] csr.mcycle\[27\] _08757_ VGND VGND VPWR
+ VPWR _08761_ sky130_fd_sc_hd__and4_1
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22283_ _06679_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24022_ _08182_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21234_ _10871_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__buf_2
Xhold230 decode.regfile.registers_31\[11\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__buf_1
Xhold241 csr._mcycle_T_3\[44\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold252 execute.io_mret_out VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_347_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_347_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold263 _03598_ VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__clkbuf_2
X_28830_ clknet_leaf_176_clock _01843_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_165_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold274 decode.regfile.registers_6\[17\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold285 csr._mcycle_T_2\[1\] VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_2
X_21165_ _06074_ _06070_ net1639 VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__and3_1
Xhold296 decode.regfile.registers_6\[13\] VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
X_20116_ _00564_ _05226_ _05326_ _05231_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__o22a_1
X_28761_ clknet_leaf_127_clock _01774_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21096_ csr.io_trapped VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__clkbuf_4
X_25973_ net2364 _09270_ _09280_ _09277_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_161_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27712_ clknet_leaf_22_clock _00741_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20047_ _00554_ _05227_ _05266_ _05267_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__a2bb2oi_1
X_24924_ net475 _08661_ _08663_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__o21a_1
X_28692_ clknet_leaf_120_clock _01705_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27643_ clknet_leaf_155_clock _00672_ VGND VGND VPWR VPWR execute.io_reg_pc\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24855_ _08615_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_124_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23806_ _07929_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__buf_4
XANTENNA_114 net2483 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24786_ _08579_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27574_ clknet_leaf_158_clock _00603_ VGND VGND VPWR VPWR csr.io_mem_pc\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_125 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21998_ csr._mcycle_T_2\[21\] _06600_ _06603_ _06592_ VGND VGND VPWR VPWR _01241_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_64_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_136 _12500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_212_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29313_ clknet_leaf_230_clock _02326_ VGND VGND VPWR VPWR decode.regfile.registers_2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23737_ net1050 csr.io_mem_pc\[31\] _08014_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26525_ _09430_ _09602_ VGND VGND VPWR VPWR _09612_ sky130_fd_sc_hd__nand2_1
XANTENNA_158 _12532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20949_ execute.io_reg_pc\[1\] _05915_ _05911_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29244_ clknet_leaf_235_clock _02257_ VGND VGND VPWR VPWR decode.regfile.registers_0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14470_ net411 _10520_ _10529_ _10522_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23668_ _07982_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26456_ _09436_ _09533_ VGND VGND VPWR VPWR _09572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22619_ _07189_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__clkbuf_2
X_25407_ _10080_ VGND VGND VPWR VPWR _08948_ sky130_fd_sc_hd__clkbuf_8
X_29175_ clknet_leaf_155_clock _02188_ VGND VGND VPWR VPWR decode.id_ex_aluop_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_26387_ net2221 _09492_ _09531_ _09525_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23599_ _07945_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16140_ _12102_ _12114_ _12115_ VGND VGND VPWR VPWR _12116_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25338_ _08891_ net2678 VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__and2_1
X_28126_ clknet_leaf_73_clock _01148_ VGND VGND VPWR VPWR csr.minstret\[31\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_134_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16071_ _11260_ _12046_ _12047_ _12048_ VGND VGND VPWR VPWR _12049_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25269_ _08864_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__clkbuf_1
X_28057_ clknet_leaf_208_clock _01079_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15022_ _11030_ VGND VGND VPWR VPWR _11031_ sky130_fd_sc_hd__buf_2
XFILLER_0_122_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27008_ clknet_leaf_342_clock _00037_ VGND VGND VPWR VPWR decode.regfile.registers_22\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19830_ _03829_ net349 _03810_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__nand3_1
XFILLER_0_20_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19761_ _04325_ _05034_ _05035_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__a21oi_1
X_28959_ clknet_leaf_180_clock _01972_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_16973_ _12829_ VGND VGND VPWR VPWR _12933_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_53_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18712_ _03657_ execute.csr_read_data_out_reg\[2\] execute.io_reg_pc\[2\] _03662_
+ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__o22a_1
X_15924_ _11075_ _11904_ _11905_ _11486_ VGND VGND VPWR VPWR _11906_ sky130_fd_sc_hd__o211a_1
X_19692_ _04963_ _04969_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 io_fetch_data[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
X_18643_ net113 _03665_ _03941_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__o21ai_1
X_15855_ decode.regfile.registers_14\[14\] _11207_ _11273_ decode.regfile.registers_15\[14\]
+ _11201_ VGND VGND VPWR VPWR _11838_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14806_ decode.id_ex_pc_reg\[19\] _10801_ _10805_ _10806_ _10848_ VGND VGND VPWR
+ VPWR _10849_ sky130_fd_sc_hd__o221a_1
X_18574_ net291 _03870_ decode.id_ex_rs2_data_reg\[23\] _03747_ _03727_ VGND VGND
+ VPWR VPWR _03873_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_204_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15786_ decode.regfile.registers_5\[12\] _11291_ _11769_ _11770_ VGND VGND VPWR VPWR
+ _11771_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_143_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17525_ decode.regfile.registers_16\[18\] _12576_ _12579_ VGND VGND VPWR VPWR _13472_
+ sky130_fd_sc_hd__o21a_1
X_14737_ _10697_ _10776_ _10778_ _10779_ VGND VGND VPWR VPWR _10780_ sky130_fd_sc_hd__o211a_1
XFILLER_0_188_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17456_ _13250_ decode.regfile.registers_24\[16\] _13170_ _13083_ _13367_ VGND VGND
+ VPWR VPWR _13405_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_200_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14668_ decode.id_ex_pc_reg\[2\] VGND VGND VPWR VPWR _10711_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16407_ _10958_ decode.regfile.registers_26\[28\] _11676_ _11338_ _10992_ VGND VGND
+ VPWR VPWR _12376_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13619_ memory.io_wb_memtoreg\[1\] _09940_ VGND VGND VPWR VPWR _09980_ sky130_fd_sc_hd__and2b_1
X_17387_ net431 _12709_ _13302_ _13337_ _13219_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__o221a_1
XFILLER_0_144_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14599_ _10640_ VGND VGND VPWR VPWR _10642_ sky130_fd_sc_hd__buf_4
XFILLER_0_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19126_ _04408_ _04414_ _04295_ _04415_ _04422_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_6_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16338_ _11646_ _11834_ _11944_ decode.regfile.registers_29\[26\] _12308_ VGND VGND
+ VPWR VPWR _12309_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19057_ _03934_ _03918_ _03989_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16269_ decode.regfile.registers_5\[25\] _11117_ _11092_ _11058_ VGND VGND VPWR VPWR
+ _12241_ sky130_fd_sc_hd__and4b_1
XFILLER_0_207_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18008_ _12968_ _03402_ _03403_ _03404_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19959_ _10678_ _03627_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_203_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22970_ csr._csr_read_data_T_8\[5\] _07416_ csr.io_mret_vector\[5\] _07417_ VGND
+ VGND VPWR VPWR _07418_ sky130_fd_sc_hd__o22a_1
XFILLER_0_214_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_199_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21921_ csr.io_mret_vector\[25\] _10773_ _06539_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_195_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24640_ net920 execute.io_target_pc\[9\] _08497_ VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__mux2_1
X_21852_ _06505_ _06494_ _06495_ _06506_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__o211a_1
X_20803_ _05876_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__clkbuf_1
X_24571_ _08467_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__clkbuf_1
X_21783_ net1062 _10777_ _06450_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23522_ net2768 _07889_ _07902_ _07893_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__o211a_1
X_26310_ net969 _09448_ _09487_ _09484_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__o211a_1
X_27290_ clknet_leaf_8_clock _00319_ VGND VGND VPWR VPWR decode.regfile.registers_31\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_20734_ _05818_ decode.id_ex_rs1_data_reg\[24\] _03585_ VGND VGND VPWR VPWR _05838_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_212_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26241_ _09025_ _09448_ VGND VGND VPWR VPWR _09449_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_83_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23453_ _10946_ _07862_ _07859_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__or3b_1
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_271_clock clknet_5_20__leaf_clock VGND VGND VPWR VPWR clknet_leaf_271_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20665_ decode.id_ex_rs1_data_reg\[0\] decode.id_ex_ex_rs1_reg\[0\] _05056_ VGND
+ VGND VPWR VPWR _05793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22404_ _06673_ _06998_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26172_ _10041_ VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__buf_4
X_23384_ fetch.bht.bhtTable_target_pc\[4\]\[29\] fetch.bht.bhtTable_target_pc\[5\]\[29\]
+ fetch.bht.bhtTable_target_pc\[6\]\[29\] fetch.bht.bhtTable_target_pc\[7\]\[29\]
+ _07669_ _07656_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__mux4_1
X_20596_ _05731_ _05734_ _05630_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__o21a_2
XFILLER_0_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25123_ _06140_ net1916 _08562_ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22335_ fetch.bht.bhtTable_tag\[4\]\[10\] fetch.bht.bhtTable_tag\[5\]\[10\] _06706_
+ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25054_ _03555_ _08747_ _08749_ _06419_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_131_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_286_clock clknet_5_20__leaf_clock VGND VGND VPWR VPWR clknet_leaf_286_clock
+ sky130_fd_sc_hd__clkbuf_8
X_29931_ clknet_leaf_337_clock _02944_ VGND VGND VPWR VPWR decode.regfile.registers_21\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22266_ _06857_ _06859_ _06860_ _06790_ _06641_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24005_ net1230 execute.io_target_pc\[23\] _08164_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__mux2_1
X_21217_ net1292 _06103_ _09912_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29862_ clknet_leaf_302_clock _02875_ VGND VGND VPWR VPWR decode.regfile.registers_19\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_22197_ _06790_ _06791_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_clock clknet_5_0__leaf_clock VGND VGND VPWR VPWR clknet_leaf_0_clock
+ sky130_fd_sc_hd__clkbuf_8
X_28813_ clknet_leaf_99_clock _01826_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_92_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21148_ _06067_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__clkbuf_1
X_29793_ clknet_leaf_309_clock _02806_ VGND VGND VPWR VPWR decode.regfile.registers_17\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28744_ clknet_leaf_99_clock _01757_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13970_ net2453 _10200_ _10239_ _10232_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__o211a_1
X_25956_ net2449 _09270_ _09271_ _09264_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__o211a_1
X_21079_ _06026_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__clkbuf_1
X_24907_ _07199_ net646 _08652_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_122_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28675_ clknet_leaf_132_clock _01688_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25887_ _08960_ _09223_ VGND VGND VPWR VPWR _09231_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_224_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_224_clock
+ sky130_fd_sc_hd__clkbuf_8
X_15640_ decode.regfile.registers_13\[8\] _11225_ _11187_ _11627_ _11628_ VGND VGND
+ VPWR VPWR _11629_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27626_ clknet_leaf_41_clock _00655_ VGND VGND VPWR VPWR execute.io_reg_pc\[3\] sky130_fd_sc_hd__dfxtp_1
X_24838_ _08606_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27557_ clknet_leaf_52_clock _00586_ VGND VGND VPWR VPWR execute.io_mem_isjump sky130_fd_sc_hd__dfxtp_1
X_15571_ _11079_ _11244_ _11261_ _11529_ _11561_ VGND VGND VPWR VPWR _11562_ sky130_fd_sc_hd__a41o_1
XFILLER_0_69_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ _08570_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17310_ _12767_ VGND VGND VPWR VPWR _13262_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14522_ _10565_ _10566_ VGND VGND VPWR VPWR _10567_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_25_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26508_ _09577_ VGND VGND VPWR VPWR _09602_ sky130_fd_sc_hd__buf_2
XFILLER_0_166_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18290_ decode.id_ex_rs2_data_reg\[11\] _03605_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27488_ clknet_leaf_157_clock _00517_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_239_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_239_clock
+ sky130_fd_sc_hd__clkbuf_8
X_29227_ clknet_leaf_139_clock _02240_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17241_ _13192_ _13193_ _13194_ VGND VGND VPWR VPWR _13195_ sky130_fd_sc_hd__o21ai_2
X_26439_ net1833 _09561_ _09562_ _09553_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__o211a_1
X_14453_ _10505_ VGND VGND VPWR VPWR _10520_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29158_ clknet_leaf_202_clock _02171_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17172_ _10938_ _12542_ _12505_ decode.regfile.registers_23\[9\] _12714_ VGND VGND
+ VPWR VPWR _13128_ sky130_fd_sc_hd__o32a_1
X_14384_ _10426_ VGND VGND VPWR VPWR _10481_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28109_ clknet_leaf_82_clock net1049 VGND VGND VPWR VPWR csr.minstret\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16123_ _11446_ decode.regfile.registers_26\[21\] _11447_ _11348_ _10993_ VGND VGND
+ VPWR VPWR _12099_ sky130_fd_sc_hd__o2111a_1
X_29089_ clknet_leaf_71_clock _02102_ VGND VGND VPWR VPWR csr._mcycle_T_3\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16054_ decode.regfile.registers_10\[19\] _10638_ _11132_ _12019_ _12031_ VGND VGND
+ VPWR VPWR _12032_ sky130_fd_sc_hd__o32a_1
XFILLER_0_84_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15005_ _11015_ _11004_ _11006_ _11007_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_55_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19813_ _04508_ _04415_ _04700_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__and3_1
XFILLER_0_209_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19744_ _05016_ _05018_ _03851_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16956_ _10928_ decode.regfile.registers_26\[4\] _12814_ _11011_ _11027_ VGND VGND
+ VPWR VPWR _12917_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_194_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15907_ _11136_ _11887_ _11888_ VGND VGND VPWR VPWR _11889_ sky130_fd_sc_hd__a21o_1
X_19675_ _04574_ _04439_ _04571_ _04949_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__a31oi_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16887_ _12847_ _12653_ _12848_ VGND VGND VPWR VPWR _12849_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18626_ memory.csr_read_data_out_reg\[16\] _09987_ _10061_ _10062_ VGND VGND VPWR
+ VPWR _03925_ sky130_fd_sc_hd__o22a_2
X_15838_ decode.regfile.registers_20\[13\] _11103_ _11327_ _11821_ VGND VGND VPWR
+ VPWR _11822_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18557_ execute.io_mem_memtoreg\[1\] execute.io_mem_memtoreg\[0\] execute.io_reg_pc\[30\]
+ _03855_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__o31a_1
X_15769_ _11679_ decode.regfile.registers_27\[11\] _11258_ VGND VGND VPWR VPWR _11755_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_190_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17508_ _12531_ _10592_ _12558_ decode.regfile.registers_0\[18\] VGND VGND VPWR VPWR
+ _13455_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18488_ net194 _03785_ _03786_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__a21boi_4
XTAP_TAPCELL_ROW_16_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_14 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17439_ decode.regfile.registers_7\[16\] _12611_ _12623_ decode.regfile.registers_6\[16\]
+ _13387_ VGND VGND VPWR VPWR _13388_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_25 _08939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_36 _10019_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_47 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _10795_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20450_ csr.minstret\[3\] _05572_ _05563_ csr._csr_read_data_T_9\[3\] VGND VGND VPWR
+ VPWR _05607_ sky130_fd_sc_hd__a22o_1
XANTENNA_69 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19109_ _03594_ _04361_ _04406_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20381_ csr.io_csr_address\[5\] _05534_ csr.io_csr_address\[6\] csr.io_csr_address\[4\]
+ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__or4b_1
XFILLER_0_125_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22120_ _06714_ _06651_ _06687_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput110 net110 VGND VGND VPWR VPWR io_memory_address[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput121 net121 VGND VGND VPWR VPWR io_memory_address[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput132 net132 VGND VGND VPWR VPWR io_memory_read sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_205_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22051_ _06645_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__buf_4
Xoutput143 net143 VGND VGND VPWR VPWR io_memory_write_data[16] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput154 net154 VGND VGND VPWR VPWR io_memory_write_data[26] sky130_fd_sc_hd__clkbuf_4
Xoutput165 net165 VGND VGND VPWR VPWR io_memory_write_data[7] sky130_fd_sc_hd__clkbuf_4
X_21002_ _05984_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_5 _00707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25810_ _08958_ _09179_ VGND VGND VPWR VPWR _09187_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_197_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26790_ _09392_ _09763_ VGND VGND VPWR VPWR _09765_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22953_ fetch.bht.bhtTable_target_pc\[8\]\[4\] fetch.bht.bhtTable_target_pc\[9\]\[4\]
+ fetch.bht.bhtTable_target_pc\[10\]\[4\] fetch.bht.bhtTable_target_pc\[11\]\[4\]
+ _07123_ _07101_ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25741_ _08964_ _09136_ VGND VGND VPWR VPWR _09147_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21904_ _06493_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_3_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28460_ clknet_leaf_148_clock _01473_ VGND VGND VPWR VPWR decode.io_id_pc\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22884_ net1223 _10771_ _07335_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__mux2_1
X_25672_ net2135 _09095_ _09106_ _09100_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__o211a_1
X_27411_ clknet_leaf_20_clock _00440_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[20\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24623_ net1008 execute.io_target_pc\[1\] _07308_ VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21835_ _06493_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__buf_2
XFILLER_0_211_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28391_ clknet_leaf_57_clock _01404_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_167_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24554_ _08458_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__clkbuf_1
X_27342_ clknet_leaf_43_clock _00371_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[15\]
+ sky130_fd_sc_hd__dfxtp_4
X_21766_ net1006 _10787_ _06439_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23505_ net92 _07889_ _07892_ _07893_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20717_ _05804_ _03596_ _05827_ net183 net2747 VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__a32o_1
X_24485_ _08111_ net2473 _08422_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27273_ clknet_leaf_12_clock _00302_ VGND VGND VPWR VPWR decode.regfile.registers_30\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21697_ _06394_ _06395_ _06396_ _06399_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29012_ clknet_leaf_119_clock _02025_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23436_ decode.immGen._imm_T_10\[0\] _07847_ _05206_ VGND VGND VPWR VPWR _07853_
+ sky130_fd_sc_hd__or3b_1
X_26224_ _10127_ VGND VGND VPWR VPWR _09436_ sky130_fd_sc_hd__buf_4
X_20648_ csr._minstret_T_3\[61\] _05556_ csr.minstret\[29\] _05658_ _05537_ VGND VGND
+ VPWR VPWR _05779_ sky130_fd_sc_hd__o221a_1
XFILLER_0_191_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26155_ _09387_ _09374_ VGND VGND VPWR VPWR _09388_ sky130_fd_sc_hd__nand2_1
X_23367_ _07075_ _07791_ _06740_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_115_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20579_ csr.minstret\[19\] _05573_ _05585_ _03554_ _05719_ VGND VGND VPWR VPWR _05720_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_225_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25106_ _08781_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__clkbuf_1
X_22318_ _06628_ _06908_ _06699_ _06912_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26086_ net641 _09343_ _09345_ _09346_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23298_ net222 net223 _07716_ VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__and3_1
X_25037_ net2542 _08735_ _06327_ _08738_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__a211oi_1
X_29914_ clknet_leaf_335_clock _02927_ VGND VGND VPWR VPWR decode.regfile.registers_21\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22249_ fetch.bht.bhtTable_tag\[12\]\[19\] fetch.bht.bhtTable_tag\[13\]\[19\] _06643_
+ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29845_ clknet_leaf_299_clock _02858_ VGND VGND VPWR VPWR decode.regfile.registers_18\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16810_ _12772_ VGND VGND VPWR VPWR _12773_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17790_ decode.regfile.registers_0\[25\] _12778_ _03191_ VGND VGND VPWR VPWR _03192_
+ sky130_fd_sc_hd__a21o_1
X_29776_ clknet_leaf_295_clock _02789_ VGND VGND VPWR VPWR decode.regfile.registers_16\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26988_ net2243 _09840_ _09877_ _06396_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_145_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28727_ clknet_leaf_132_clock _01740_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_16741_ _12487_ _12700_ _12703_ _12705_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_163_clock clknet_5_25__leaf_clock VGND VGND VPWR VPWR clknet_leaf_163_clock
+ sky130_fd_sc_hd__clkbuf_8
X_13953_ net2592 _10226_ _10230_ _10219_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__o211a_1
X_25939_ _08937_ _09253_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19460_ _04452_ _04742_ _04743_ _04526_ _04746_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__o32a_1
X_28658_ clknet_leaf_108_clock _01671_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16672_ decode.immGen._imm_T_24\[16\] _10614_ VGND VGND VPWR VPWR _12637_ sky130_fd_sc_hd__nand2_8
XFILLER_0_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13884_ net2554 _10180_ _10189_ _10188_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18411_ csr.io_csr_address\[1\] VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__buf_6
X_27609_ clknet_leaf_159_clock _00638_ VGND VGND VPWR VPWR execute.io_target_pc\[18\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_9_1253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15623_ _10957_ decode.regfile.registers_22\[8\] _11450_ _10978_ _10990_ VGND VGND
+ VPWR VPWR _11612_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_186_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_204 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19391_ _04386_ _04677_ _04678_ _04680_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_48_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28589_ clknet_leaf_103_clock _01602_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_215 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_226 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_178_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_178_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_185_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18342_ _03640_ decode.id_ex_ex_rs1_reg\[3\] VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_237 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_248 net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15554_ _11536_ _11544_ _11289_ VGND VGND VPWR VPWR _11545_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_104_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_259 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14505_ _10548_ _09917_ _09916_ _10549_ VGND VGND VPWR VPWR _10550_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18273_ decode.id_ex_rs2_data_reg\[3\] _03596_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15485_ decode.regfile.registers_18\[4\] _11455_ _11456_ _11477_ VGND VGND VPWR VPWR
+ _11478_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17224_ _12496_ _13175_ _13177_ _13178_ VGND VGND VPWR VPWR _13179_ sky130_fd_sc_hd__a31o_1
X_14436_ _09970_ _10507_ VGND VGND VPWR VPWR _10511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_101_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_101_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 net376 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_896 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput23 net387 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput34 io_memory_read_data[0] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput45 io_memory_read_data[1] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
X_17155_ decode.regfile.registers_8\[9\] _12892_ _12603_ _13110_ VGND VGND VPWR VPWR
+ _13111_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14367_ _09993_ _10464_ VGND VGND VPWR VPWR _10471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput56 io_memory_read_data[2] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xhold807 fetch.bht.bhtTable_tag\[12\]\[6\] VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16106_ decode.regfile.registers_20\[20\] _11452_ _12081_ _12082_ _11223_ VGND VGND
+ VPWR VPWR _12083_ sky130_fd_sc_hd__a221o_1
Xhold818 decode.regfile.registers_13\[8\] VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold829 fetch.bht.bhtTable_tag\[8\]\[10\] VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__dlygate4sd3_1
X_17086_ _12516_ _13040_ _13042_ _13043_ VGND VGND VPWR VPWR _13044_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14298_ _10418_ VGND VGND VPWR VPWR _10431_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_208_Right_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_116_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_116_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16037_ _11942_ decode.regfile.registers_30\[19\] _11722_ _11723_ _11724_ VGND VGND
+ VPWR VPWR _12015_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_23_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2208 fetch.bht.bhtTable_target_pc\[0\]\[31\] VGND VGND VPWR VPWR net2435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2219 decode.regfile.registers_9\[7\] VGND VGND VPWR VPWR net2446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_200_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1507 _01228_ VGND VGND VPWR VPWR net1734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1518 fetch.bht.bhtTable_tag\[14\]\[6\] VGND VGND VPWR VPWR net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_28__f_clock clknet_2_3_0_clock VGND VGND VPWR VPWR clknet_5_28__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_17988_ _03381_ _03383_ _03384_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__a21oi_2
Xhold1529 fetch.bht.bhtTable_target_pc\[10\]\[31\] VGND VGND VPWR VPWR net1756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19727_ _03639_ _04991_ _03881_ _04589_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__o31a_1
XFILLER_0_97_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16939_ _11020_ _12559_ _12534_ VGND VGND VPWR VPWR _12900_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19658_ _04935_ _04912_ _04936_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_220_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18609_ net248 VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__buf_6
XFILLER_0_94_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19589_ _04210_ _04860_ _04841_ _04870_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21620_ _05613_ csr.minstret\[5\] csr.io_inst_retired _06333_ VGND VGND VPWR VPWR
+ _06342_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21551_ _06122_ net2268 _06295_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20502_ csr.minstret\[9\] _05573_ _05585_ csr.mcycle\[9\] _05652_ VGND VGND VPWR
+ VPWR _05653_ sky130_fd_sc_hd__a221o_1
X_24270_ _08310_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21482_ _06111_ net1460 _06252_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23221_ _07107_ fetch.bht.bhtTable_target_pc\[14\]\[19\] VGND VGND VPWR VPWR _07655_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_160_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20433_ _03718_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23152_ net72 net225 net226 _07530_ net73 VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__a41o_1
XFILLER_0_144_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20364_ csr.io_csr_address\[11\] net218 _05520_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__and3b_1
XFILLER_0_141_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22103_ _06636_ _06689_ _06697_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_149_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23083_ fetch.bht.bhtTable_target_pc\[0\]\[11\] fetch.bht.bhtTable_target_pc\[1\]\[11\]
+ fetch.bht.bhtTable_target_pc\[2\]\[11\] fetch.bht.bhtTable_target_pc\[3\]\[11\]
+ _07407_ _07115_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__mux4_1
X_27960_ clknet_leaf_170_clock _00982_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_149_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20295_ _05472_ _05219_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22034_ _06628_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_181_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26911_ net2597 _09822_ _09833_ _09825_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_181_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27891_ clknet_leaf_22_clock _00920_ VGND VGND VPWR VPWR csr._mcycle_T_2\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_220_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_80_clock
+ sky130_fd_sc_hd__clkbuf_8
X_29630_ clknet_leaf_288_clock _02643_ VGND VGND VPWR VPWR decode.regfile.registers_12\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26842_ _09793_ VGND VGND VPWR VPWR _09794_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_215_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29561_ clknet_leaf_313_clock _02574_ VGND VGND VPWR VPWR decode.regfile.registers_9\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_26773_ net1731 _09752_ _09755_ _09743_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__o211a_1
X_23985_ net979 VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28512_ clknet_leaf_195_clock _01525_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25724_ net1315 _09125_ _09137_ _09129_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__o211a_1
X_22936_ _06661_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__buf_4
X_29492_ clknet_leaf_264_clock _02505_ VGND VGND VPWR VPWR decode.regfile.registers_7\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_95_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_95_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_218_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28443_ clknet_leaf_55_clock _01456_ VGND VGND VPWR VPWR decode.io_id_pc\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25655_ net2381 _09095_ _09097_ _09087_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__o211a_1
X_22867_ net910 _10795_ _07324_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24606_ _08485_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28374_ clknet_leaf_200_clock _01387_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_21818_ _06481_ csr.io_interrupt _06316_ _06470_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_175_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22798_ net1237 _10871_ _07286_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__mux2_1
X_25586_ net2379 _09052_ _09057_ _09046_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27325_ clknet_leaf_24_clock _00354_ VGND VGND VPWR VPWR decode.id_ex_funct3_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_94_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24537_ _08097_ net1531 _09902_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__mux2_1
X_21749_ net824 _10872_ _06428_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15270_ _11263_ decode.regfile.registers_22\[1\] _11093_ _11264_ _11265_ VGND VGND
+ VPWR VPWR _11266_ sky130_fd_sc_hd__o2111a_1
X_27256_ clknet_leaf_8_clock _00285_ VGND VGND VPWR VPWR decode.regfile.registers_30\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_24468_ _08095_ net1921 _08411_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26207_ _09424_ _09413_ VGND VGND VPWR VPWR _09425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14221_ net614 _10376_ _10386_ _10385_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_78_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23419_ _07834_ _07840_ _06637_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__mux2_2
X_24399_ net1189 execute.io_target_pc\[22\] _08367_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__mux2_1
X_27187_ clknet_leaf_6_clock _00216_ VGND VGND VPWR VPWR decode.regfile.registers_28\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14152_ _10031_ _10342_ VGND VGND VPWR VPWR _10347_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_33_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_33_clock
+ sky130_fd_sc_hd__clkbuf_8
X_26138_ net2170 _09373_ _09376_ _09370_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14083_ _10048_ _10299_ VGND VGND VPWR VPWR _10307_ sky130_fd_sc_hd__nand2_1
X_18960_ _04249_ _04250_ _04258_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__o21ai_1
X_26069_ net2176 _09329_ _09336_ _09333_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__o211a_1
X_17911_ decode.regfile.registers_1\[28\] _12631_ _12933_ _03309_ VGND VGND VPWR VPWR
+ _03310_ sky130_fd_sc_hd__o211ai_2
X_18891_ _04189_ _03894_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_218_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_48_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_48_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_37_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17842_ decode.regfile.registers_13\[26\] _12534_ _12588_ VGND VGND VPWR VPWR _03243_
+ sky130_fd_sc_hd__and3_1
X_29828_ clknet_leaf_303_clock _02841_ VGND VGND VPWR VPWR decode.regfile.registers_18\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17773_ _13250_ decode.regfile.registers_24\[24\] _12997_ _12998_ _13367_ VGND VGND
+ VPWR VPWR _03176_ sky130_fd_sc_hd__o2111a_1
X_29759_ clknet_leaf_311_clock _02772_ VGND VGND VPWR VPWR decode.regfile.registers_16\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14985_ _10962_ _10997_ _11002_ net2713 _10949_ VGND VGND VPWR VPWR _11003_ sky130_fd_sc_hd__a32o_1
XFILLER_0_156_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19512_ _04780_ _04789_ _04796_ _04242_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16724_ _12528_ _12684_ _12688_ VGND VGND VPWR VPWR _12689_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13936_ _10064_ _10210_ VGND VGND VPWR VPWR _10221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19443_ _04618_ _04306_ _04712_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_18_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16655_ _12619_ VGND VGND VPWR VPWR _12620_ sky130_fd_sc_hd__clkbuf_4
X_13867_ _10152_ VGND VGND VPWR VPWR _10180_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15606_ decode.regfile.registers_18\[7\] _11269_ _11271_ VGND VGND VPWR VPWR _11596_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_215_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19374_ _04126_ _04129_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__nand2_1
X_16586_ _12550_ VGND VGND VPWR VPWR _12551_ sky130_fd_sc_hd__buf_4
X_13798_ memory.io_wb_reg_pc\[29\] _09946_ _09947_ _10133_ VGND VGND VPWR VPWR _10134_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18325_ _03628_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15537_ _10962_ decode.regfile.registers_30\[6\] _11039_ _11032_ _11033_ VGND VGND
+ VPWR VPWR _11528_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18256_ _03585_ _03588_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__nor2_2
X_15468_ decode.regfile.registers_3\[4\] _11110_ _11142_ _11146_ _11460_ VGND VGND
+ VPWR VPWR _11461_ sky130_fd_sc_hd__a311o_1
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17207_ decode.regfile.registers_18\[10\] _12571_ _12561_ _13161_ VGND VGND VPWR
+ VPWR _13162_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14419_ _10128_ _10462_ VGND VGND VPWR VPWR _10500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18187_ decode.control.io_funct7\[2\] decode.control.io_funct7\[0\] _03523_ _03524_
+ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15399_ decode.regfile.registers_24\[2\] _11074_ _11352_ _11393_ VGND VGND VPWR VPWR
+ _11394_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17138_ _12496_ _13090_ _13092_ _13094_ VGND VGND VPWR VPWR _13095_ sky130_fd_sc_hd__a31o_1
Xhold604 decode.regfile.registers_22\[8\] VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 fetch.bht.bhtTable_tag\[8\]\[7\] VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 _08231_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold637 decode.regfile.registers_26\[4\] VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 fetch.bht.bhtTable_target_pc\[4\]\[15\] VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 fetch.bht.bhtTable_target_pc\[2\]\[29\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17069_ decode.regfile.registers_11\[7\] _12595_ _12587_ _12551_ _13026_ VGND VGND
+ VPWR VPWR _13027_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_111_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20080_ decode.id_ex_imm_reg\[12\] decode.id_ex_pc_reg\[12\] VGND VGND VPWR VPWR
+ _05295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2005 decode.regfile.registers_25\[17\] VGND VGND VPWR VPWR net2232 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 decode.regfile.registers_21\[30\] VGND VGND VPWR VPWR net2243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2027 decode.regfile.registers_3\[21\] VGND VGND VPWR VPWR net2254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2038 fetch.bht.bhtTable_target_pc\[0\]\[15\] VGND VGND VPWR VPWR net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1304 fetch.bht.bhtTable_target_pc\[10\]\[23\] VGND VGND VPWR VPWR net1531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_191_Right_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2049 decode.regfile.registers_20\[1\] VGND VGND VPWR VPWR net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1315 fetch.bht.bhtTable_target_pc\[9\]\[14\] VGND VGND VPWR VPWR net1542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1326 fetch.bht.bhtTable_tag\[7\]\[12\] VGND VGND VPWR VPWR net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1337 fetch.bht.bhtTable_target_pc\[6\]\[20\] VGND VGND VPWR VPWR net1564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1348 fetch.bht.bhtTable_tag\[9\]\[10\] VGND VGND VPWR VPWR net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1359 fetch.bht.bhtTable_tag\[0\]\[7\] VGND VGND VPWR VPWR net1586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23770_ _06132_ net1399 _08030_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20982_ execute.io_reg_pc\[16\] _05965_ _05973_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22721_ _10946_ _10964_ _10952_ _07249_ _07251_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__a41o_1
XFILLER_0_67_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25440_ _08970_ _08905_ VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__nand2_1
X_22652_ net2645 _07210_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_217_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21603_ csr._mcycle_T_2\[2\] _06329_ _06328_ csr.minstret\[2\] VGND VGND VPWR VPWR
+ _06330_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22583_ csr._minstret_T_3\[42\] csr._minstret_T_3\[41\] _07162_ VGND VGND VPWR VPWR
+ _07166_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25371_ _08905_ VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__buf_2
XFILLER_0_164_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27110_ clknet_leaf_348_clock _00139_ VGND VGND VPWR VPWR decode.regfile.registers_25\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_24322_ _08337_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__clkbuf_1
X_21534_ _06105_ net1693 _06284_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28090_ clknet_leaf_190_clock _01112_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_170_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24253_ _08081_ net1825 _08300_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27041_ clknet_leaf_345_clock _00070_ VGND VGND VPWR VPWR decode.regfile.registers_23\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_21465_ net12 _10673_ _10911_ _09957_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__o31a_1
XFILLER_0_65_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23204_ fetch.bht.bhtTable_target_pc\[4\]\[18\] fetch.bht.bhtTable_target_pc\[5\]\[18\]
+ fetch.bht.bhtTable_target_pc\[6\]\[18\] fetch.bht.bhtTable_target_pc\[7\]\[18\]
+ _07384_ _07113_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__mux4_1
X_20416_ _05559_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__clkbuf_4
X_24184_ _06250_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__buf_4
XFILLER_0_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21396_ _06211_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23135_ fetch.bht.bhtTable_target_pc\[0\]\[14\] fetch.bht.bhtTable_target_pc\[1\]\[14\]
+ fetch.bht.bhtTable_target_pc\[2\]\[14\] fetch.bht.bhtTable_target_pc\[3\]\[14\]
+ _07099_ _07103_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__mux4_1
X_20347_ decode.id_ex_pc_reg\[30\] _05508_ _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_73_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28992_ clknet_leaf_170_clock _02005_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23066_ fetch.bht.bhtTable_target_pc\[12\]\[10\] fetch.bht.bhtTable_target_pc\[13\]\[10\]
+ _07123_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__mux2_1
X_27943_ clknet_leaf_220_clock _00965_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20278_ _05458_ _05459_ _05420_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__o21ai_1
X_22017_ csr._mcycle_T_2\[30\] _06571_ _06613_ _06605_ VGND VGND VPWR VPWR _01250_
+ sky130_fd_sc_hd__o211a_1
X_27874_ clknet_leaf_70_clock _00903_ VGND VGND VPWR VPWR csr.io_inst_retired sky130_fd_sc_hd__dfxtp_2
XFILLER_0_179_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2550 net78 VGND VGND VPWR VPWR net2777 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29613_ clknet_leaf_279_clock _02626_ VGND VGND VPWR VPWR decode.regfile.registers_11\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_26825_ _09428_ _09776_ VGND VGND VPWR VPWR _09785_ sky130_fd_sc_hd__nand2_1
Xhold2561 decode.regfile.registers_30\[27\] VGND VGND VPWR VPWR net2788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2572 csr._mcycle_T_2\[5\] VGND VGND VPWR VPWR net2799 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1860 fetch.bht.bhtTable_target_pc\[5\]\[31\] VGND VGND VPWR VPWR net2087 sky130_fd_sc_hd__dlygate4sd3_1
X_29544_ clknet_leaf_266_clock _02557_ VGND VGND VPWR VPWR decode.regfile.registers_9\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1871 fetch.bht.bhtTable_target_pc\[8\]\[3\] VGND VGND VPWR VPWR net2098 sky130_fd_sc_hd__dlygate4sd3_1
X_14770_ csr.io_mem_pc\[10\] _10762_ VGND VGND VPWR VPWR _10813_ sky130_fd_sc_hd__nand2_1
X_26756_ _09434_ _09733_ VGND VGND VPWR VPWR _09745_ sky130_fd_sc_hd__nand2_1
X_23968_ net866 execute.io_target_pc\[5\] _08153_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__mux2_1
Xhold1882 decode.regfile.registers_18\[20\] VGND VGND VPWR VPWR net2109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1893 decode.regfile.registers_20\[14\] VGND VGND VPWR VPWR net2120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13721_ _10068_ VGND VGND VPWR VPWR _10069_ sky130_fd_sc_hd__clkbuf_8
X_25707_ _10130_ VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__clkbuf_4
X_22919_ fetch.bht.bhtTable_target_pc\[0\]\[2\] fetch.bht.bhtTable_target_pc\[1\]\[2\]
+ fetch.bht.bhtTable_target_pc\[2\]\[2\] fetch.bht.bhtTable_target_pc\[3\]\[2\] _07119_
+ _07071_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__mux4_1
XFILLER_0_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29475_ clknet_leaf_253_clock _02488_ VGND VGND VPWR VPWR decode.regfile.registers_7\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26687_ _09441_ _09664_ VGND VGND VPWR VPWR _09705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23899_ _06155_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28426_ clknet_leaf_246_clock _01439_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_16440_ decode.regfile.registers_20\[29\] _11452_ _12406_ _12407_ _11223_ VGND VGND
+ VPWR VPWR _12408_ sky130_fd_sc_hd__a221o_1
X_25638_ _08937_ _09079_ VGND VGND VPWR VPWR _09088_ sky130_fd_sc_hd__nand2_1
X_13652_ net2063 _09938_ _10009_ _09957_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28357_ clknet_leaf_237_clock _01370_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16371_ _12339_ _11486_ _12340_ VGND VGND VPWR VPWR _12341_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25569_ _08943_ _09036_ VGND VGND VPWR VPWR _09048_ sky130_fd_sc_hd__nand2_1
X_13583_ _09946_ _09947_ memory.io_wb_reg_pc\[0\] VGND VGND VPWR VPWR _09948_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18110_ _10575_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__buf_2
XFILLER_0_183_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27308_ clknet_leaf_13_clock _00337_ VGND VGND VPWR VPWR decode.regfile.registers_31\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15322_ _11314_ VGND VGND VPWR VPWR _11318_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19090_ _03635_ _03634_ _04299_ _03633_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__or4b_2
X_28288_ clknet_leaf_85_clock _01310_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_671 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18041_ _11014_ _10936_ decode.regfile.registers_23\[31\] _12995_ VGND VGND VPWR
+ VPWR _03437_ sky130_fd_sc_hd__or4_1
X_27239_ clknet_leaf_0_clock _00268_ VGND VGND VPWR VPWR decode.regfile.registers_29\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15253_ _11040_ _11241_ _11247_ _11249_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14204_ _10375_ VGND VGND VPWR VPWR _10377_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15184_ _11180_ VGND VGND VPWR VPWR _11181_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14135_ _09975_ _10333_ VGND VGND VPWR VPWR _10337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19992_ _05221_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18943_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__clkbuf_4
X_14066_ _09999_ _10288_ VGND VGND VPWR VPWR _10297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18874_ _04062_ _04065_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__and2_2
XFILLER_0_207_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17825_ decode.regfile.registers_20\[26\] _12546_ _12553_ _12554_ _12538_ VGND VGND
+ VPWR VPWR _03226_ sky130_fd_sc_hd__a41o_1
XFILLER_0_94_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17756_ _03153_ _03156_ _03157_ _03158_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__o211a_1
X_14968_ _10992_ VGND VGND VPWR VPWR _10993_ sky130_fd_sc_hd__buf_2
XFILLER_0_221_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16707_ _11019_ _12550_ _12559_ VGND VGND VPWR VPWR _12672_ sky130_fd_sc_hd__and3_2
X_13919_ net591 _10199_ _10211_ _10206_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17687_ decode.regfile.registers_13\[22\] _12774_ _03090_ _03091_ _12662_ VGND VGND
+ VPWR VPWR _03092_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14899_ decode.immGen._imm_T_24\[17\] VGND VGND VPWR VPWR _10934_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19426_ _04359_ net278 _04394_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16638_ _12602_ VGND VGND VPWR VPWR _12603_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19357_ _04647_ _04591_ _04248_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__mux2_1
X_16569_ _12533_ VGND VGND VPWR VPWR _12534_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18308_ _03619_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19288_ _04443_ _04073_ _04446_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_212_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_212_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18239_ net699 csr._mcycle_T_3\[59\] _03568_ _03573_ VGND VGND VPWR VPWR _03574_
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21250_ csr.io_mem_pc\[18\] VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__buf_2
XFILLER_0_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold401 decode.regfile.registers_14\[8\] VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold412 decode.regfile.registers_18\[13\] VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 net67 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20201_ decode.id_ex_imm_reg\[29\] _10697_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__nor2_1
Xhold434 decode.regfile.registers_30\[5\] VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21181_ _06085_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold445 decode.regfile.registers_7\[3\] VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold456 decode.regfile.registers_9\[11\] VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold467 decode.regfile.registers_28\[11\] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20132_ decode.id_ex_pc_reg\[19\] VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__buf_2
Xhold478 decode.regfile.registers_20\[15\] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold489 decode.regfile.registers_16\[3\] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_221_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20063_ _05278_ _05280_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__xor2_1
X_24940_ net2347 _08672_ _08673_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_110_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1101 fetch.bht.bhtTable_target_pc\[4\]\[12\] VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 fetch.bht.bhtTable_target_pc\[8\]\[12\] VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 fetch.bht.bhtTable_tag\[3\]\[17\] VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__dlygate4sd3_1
X_24871_ _08623_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1134 fetch.bht.bhtTable_target_pc\[10\]\[3\] VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 fetch.bht.bhtTable_target_pc\[5\]\[14\] VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1156 fetch.bht.bhtTable_target_pc\[7\]\[18\] VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__dlygate4sd3_1
X_26610_ net2455 _09649_ _09659_ _09660_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23822_ _08068_ net1311 _08058_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1167 decode.regfile.registers_4\[2\] VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27590_ clknet_leaf_149_clock _00619_ VGND VGND VPWR VPWR csr.io_mem_pc\[31\] sky130_fd_sc_hd__dfxtp_4
Xhold1178 decode.regfile.registers_1\[31\] VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 decode.regfile.registers_19\[18\] VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_219_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26541_ _09620_ VGND VGND VPWR VPWR _09621_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_219_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23753_ _06115_ net1279 _09907_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__mux2_1
X_20965_ _05964_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22704_ csr._mcycle_T_2\[26\] _07236_ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__or2_1
X_29260_ clknet_leaf_233_clock _02273_ VGND VGND VPWR VPWR decode.regfile.registers_0\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26472_ net2330 _09578_ _09581_ _09582_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23684_ _07991_ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__buf_4
XFILLER_0_165_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20896_ _05927_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_172_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28211_ clknet_leaf_82_clock net882 VGND VGND VPWR VPWR csr.mscratch\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25423_ net459 _08951_ _08959_ _08950_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22635_ csr._minstret_T_3\[59\] csr._minstret_T_3\[58\] _07196_ net1392 VGND VGND
+ VPWR VPWR _07200_ sky130_fd_sc_hd__a31oi_1
X_29191_ clknet_leaf_240_clock _02204_ VGND VGND VPWR VPWR fetch.btb.btbTable\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28142_ clknet_leaf_208_clock _01164_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22566_ csr._minstret_T_3\[38\] csr._minstret_T_3\[37\] csr._minstret_T_3\[36\] _07151_
+ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__and4_1
X_25354_ net1856 _08906_ _08911_ _07247_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24305_ _08328_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__clkbuf_1
X_21517_ _06276_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__clkbuf_1
X_28073_ clknet_leaf_222_clock _01095_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_22497_ execute.io_target_pc\[0\] _07091_ _06041_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__a21o_1
XFILLER_0_161_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25285_ _08869_ decode.regfile.registers_0\[4\] VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27024_ clknet_leaf_333_clock _00053_ VGND VGND VPWR VPWR decode.regfile.registers_23\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21448_ _06239_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__clkbuf_1
X_24236_ _08064_ net1985 _08289_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24167_ _08257_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21379_ _06202_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23118_ fetch.bht.bhtTable_target_pc\[12\]\[13\] fetch.bht.bhtTable_target_pc\[13\]\[13\]
+ fetch.bht.bhtTable_target_pc\[14\]\[13\] fetch.bht.bhtTable_target_pc\[15\]\[13\]
+ _07099_ _07101_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_92_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28975_ clknet_leaf_107_clock _01988_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_24098_ net1519 execute.io_target_pc\[4\] _08221_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold990 fetch.bht.bhtTable_target_pc\[13\]\[24\] VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23049_ fetch.bht.bhtTable_target_pc\[4\]\[9\] fetch.bht.bhtTable_target_pc\[5\]\[9\]
+ fetch.bht.bhtTable_target_pc\[6\]\[9\] fetch.bht.bhtTable_target_pc\[7\]\[9\] _07123_
+ _07111_ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__mux4_1
X_15940_ decode.regfile.registers_7\[16\] _11465_ _11466_ decode.regfile.registers_6\[16\]
+ _11281_ VGND VGND VPWR VPWR _11921_ sky130_fd_sc_hd__a221oi_1
X_27926_ clknet_leaf_42_clock _00955_ VGND VGND VPWR VPWR execute.io_mem_rd\[2\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_129_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27857_ clknet_leaf_322_clock _00886_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15871_ _11840_ _11852_ _11853_ VGND VGND VPWR VPWR _11854_ sky130_fd_sc_hd__o21a_1
XFILLER_0_215_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17610_ _12901_ _03015_ _03016_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__o21a_1
Xhold2380 decode.regfile.registers_23\[24\] VGND VGND VPWR VPWR net2607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14822_ _10800_ _10765_ _10795_ VGND VGND VPWR VPWR _10865_ sky130_fd_sc_hd__a21oi_1
X_26808_ _09410_ _09763_ VGND VGND VPWR VPWR _09775_ sky130_fd_sc_hd__nand2_1
Xhold2391 decode.regfile.registers_11\[23\] VGND VGND VPWR VPWR net2618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18590_ _03706_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27788_ clknet_leaf_334_clock _00817_ VGND VGND VPWR VPWR memory.io_wb_readdata\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1690 fetch.bht.bhtTable_tag\[8\]\[22\] VGND VGND VPWR VPWR net1917 sky130_fd_sc_hd__dlygate4sd3_1
X_17541_ _13091_ _13176_ decode.regfile.registers_27\[18\] _13487_ VGND VGND VPWR
+ VPWR _13488_ sky130_fd_sc_hd__or4_1
X_29527_ clknet_leaf_266_clock _02540_ VGND VGND VPWR VPWR decode.regfile.registers_8\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_14753_ csr.io_mem_pc\[19\] _10795_ _10765_ VGND VGND VPWR VPWR _10796_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26739_ net1544 _09723_ _09735_ _09730_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_103_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13704_ net687 _10027_ _10054_ _10020_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_138_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17472_ decode.regfile.registers_13\[17\] _12927_ _12588_ _12663_ VGND VGND VPWR
+ VPWR _13420_ sky130_fd_sc_hd__a31o_1
X_29458_ clknet_leaf_261_clock _02471_ VGND VGND VPWR VPWR decode.regfile.registers_6\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_14684_ _10707_ execute.io_target_pc\[9\] _10725_ execute.io_target_pc\[25\] _10726_
+ VGND VGND VPWR VPWR _10727_ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19211_ _04477_ _04491_ _04492_ _04502_ _04506_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__a32o_1
XFILLER_0_128_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28409_ clknet_leaf_170_clock _01422_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_1
X_16423_ _11043_ decode.regfile.registers_4\[29\] _11503_ _10629_ _11083_ VGND VGND
+ VPWR VPWR _12391_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_6_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13635_ net1572 _09938_ _09994_ _09957_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__o211a_1
X_29389_ clknet_leaf_258_clock _02402_ VGND VGND VPWR VPWR decode.regfile.registers_4\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19142_ _04438_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_60_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16354_ decode.regfile.registers_8\[27\] _11045_ _11174_ VGND VGND VPWR VPWR _12324_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_229_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13566_ decode.io_wb_rd\[1\] VGND VGND VPWR VPWR _09931_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15305_ _11300_ decode.regfile.registers_0\[1\] VGND VGND VPWR VPWR _11301_ sky130_fd_sc_hd__nand2_1
X_19073_ _04290_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16285_ decode.regfile.registers_16\[25\] _11122_ _12239_ _12256_ VGND VGND VPWR
+ VPWR _12257_ sky130_fd_sc_hd__o22a_1
X_13497_ csr.io_mem_pc\[4\] VGND VGND VPWR VPWR _09879_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18024_ _12603_ _03419_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15236_ decode.regfile.registers_22\[0\] _11096_ _11230_ _11232_ VGND VGND VPWR VPWR
+ _11233_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15167_ net319 _11041_ _11143_ VGND VGND VPWR VPWR _11164_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14118_ _10136_ _10286_ VGND VGND VPWR VPWR _10326_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_58_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19975_ net2620 _05217_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__nor2_1
X_15098_ _11048_ _11093_ _11094_ _10976_ VGND VGND VPWR VPWR _11095_ sky130_fd_sc_hd__and4_1
XFILLER_0_157_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18926_ _03637_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__clkbuf_4
X_14049_ _10285_ VGND VGND VPWR VPWR _10286_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18857_ memory.csr_read_data_out_reg\[10\] _10010_ _10028_ _10029_ VGND VGND VPWR
+ VPWR _04156_ sky130_fd_sc_hd__o22a_2
XFILLER_0_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17808_ decode.regfile.registers_18\[25\] _12566_ _03188_ _03209_ VGND VGND VPWR
+ VPWR _03210_ sky130_fd_sc_hd__o22a_1
XFILLER_0_171_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18788_ _10056_ _10055_ _10010_ memory.csr_read_data_out_reg\[15\] VGND VGND VPWR
+ VPWR _04087_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_59_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17739_ _02990_ _03068_ decode.regfile.registers_27\[23\] _13487_ VGND VGND VPWR
+ VPWR _03143_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20750_ _05627_ _05671_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19409_ _04503_ _04696_ _04697_ _04242_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__o31a_1
XFILLER_0_92_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20681_ _05630_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22420_ _06690_ _07012_ _06672_ _07014_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22351_ _06672_ _06945_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21302_ net1204 _10817_ _06157_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_130_Left_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25070_ net1947 _08759_ _08760_ _06327_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22282_ _06642_ _06870_ _06876_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24021_ net1007 execute.io_target_pc\[31\] _07960_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21233_ _06114_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold220 csr._mcycle_T_3\[63\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold231 decode.regfile.registers_30\[9\] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold242 decode.regfile.registers_31\[18\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold253 decode.regfile.registers_12\[7\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 decode.regfile.registers_24\[9\] VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
X_21164_ _06076_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_165_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold275 csr._mcycle_T_3\[52\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold286 _01185_ VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold297 csr._mcycle_T_3\[39\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
X_20115_ _05321_ _05325_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__xnor2_1
X_28760_ clknet_leaf_121_clock _01773_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21095_ _06036_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_1170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25972_ _08968_ _09241_ VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_161_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27711_ clknet_leaf_20_clock _00740_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20046_ _05222_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__inv_2
X_24923_ _06318_ _08662_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_217_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28691_ clknet_leaf_140_clock _01704_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27642_ clknet_leaf_45_clock _00671_ VGND VGND VPWR VPWR execute.io_reg_pc\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24854_ _06132_ net1261 _08607_ VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23805_ execute.io_target_pc\[4\] VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27573_ clknet_leaf_159_clock _00602_ VGND VGND VPWR VPWR csr.io_mem_pc\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_104 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24785_ _08078_ net1229 _08574_ VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_115 net2754 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ net2390 _06601_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__or2_1
XANTENNA_126 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29312_ clknet_leaf_244_clock _02325_ VGND VGND VPWR VPWR decode.regfile.registers_2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_137 _12532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26524_ net2574 _09605_ _09611_ _09608_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__o211a_1
X_23736_ _08019_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _12532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20948_ _05955_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29243_ clknet_leaf_232_clock _02256_ VGND VGND VPWR VPWR decode.regfile.registers_0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26455_ net2721 _09561_ _09571_ _09567_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__o211a_1
X_23667_ net798 _10773_ _07972_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__mux2_1
X_20879_ _05858_ _09956_ net45 VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__and3_1
XFILLER_0_181_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25406_ net2744 _08928_ _08947_ _08927_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22618_ csr._minstret_T_3\[54\] csr._minstret_T_3\[53\] csr._minstret_T_3\[52\] _07185_
+ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__and4_1
X_29174_ clknet_leaf_155_clock _02187_ VGND VGND VPWR VPWR decode.id_ex_aluop_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26386_ _09443_ _09490_ VGND VGND VPWR VPWR _09531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23598_ _06128_ net1974 _07941_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28125_ clknet_leaf_78_clock _01147_ VGND VGND VPWR VPWR csr.minstret\[30\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_23_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25337_ _08899_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22549_ csr._minstret_T_3\[33\] csr._minstret_T_3\[32\] csr.minstret\[30\] csr.minstret\[31\]
+ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28056_ clknet_leaf_203_clock _01078_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16070_ _11436_ decode.regfile.registers_26\[19\] _11676_ _11338_ _11564_ VGND VGND
+ VPWR VPWR _12048_ sky130_fd_sc_hd__o2111a_1
X_25268_ _08107_ net1255 _09906_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15021_ _10667_ _10954_ _10997_ decode.control.io_funct7\[6\] _10973_ VGND VGND VPWR
+ VPWR _11030_ sky130_fd_sc_hd__o311a_1
X_27007_ clknet_leaf_342_clock _00036_ VGND VGND VPWR VPWR decode.regfile.registers_22\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_24219_ _08113_ net2087 _06251_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25199_ net422 _08828_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16972_ _12630_ VGND VGND VPWR VPWR _12932_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19760_ _03888_ _04320_ _04265_ _04249_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__o211a_1
X_28958_ clknet_leaf_131_clock _01971_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15923_ decode.regfile.registers_25\[15\] _11483_ _11484_ decode.regfile.registers_24\[15\]
+ VGND VGND VPWR VPWR _11905_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_53_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18711_ _09967_ _09968_ memory.csr_read_data_out_reg\[2\] _09942_ VGND VGND VPWR
+ VPWR _04010_ sky130_fd_sc_hd__o2bb2a_2
X_19691_ _04546_ _04966_ _04303_ _04967_ _04968_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__o311a_1
X_27909_ clknet_leaf_18_clock _00938_ VGND VGND VPWR VPWR csr._mcycle_T_2\[30\] sky130_fd_sc_hd__dfxtp_2
X_28889_ clknet_leaf_127_clock _01902_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_18642_ _03658_ execute.csr_read_data_out_reg\[21\] execute.io_reg_pc\[21\] _03776_
+ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__o22a_1
X_15854_ decode.regfile.registers_18\[14\] _11225_ _11113_ _10988_ _10976_ VGND VGND
+ VPWR VPWR _11837_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_204_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14805_ _10845_ _10846_ _10847_ VGND VGND VPWR VPWR _10848_ sky130_fd_sc_hd__and3_1
X_18573_ _03868_ _03700_ _03688_ decode.id_ex_rs1_data_reg\[23\] _03871_ VGND VGND
+ VPWR VPWR _03872_ sky130_fd_sc_hd__o221a_4
XFILLER_0_118_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15785_ _11044_ decode.regfile.registers_4\[12\] _10648_ _10631_ _11084_ VGND VGND
+ VPWR VPWR _11770_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_188_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17524_ decode.regfile.registers_15\[18\] _12585_ _13469_ _13470_ _12673_ VGND VGND
+ VPWR VPWR _13471_ sky130_fd_sc_hd__a221o_1
X_14736_ _10777_ _10684_ VGND VGND VPWR VPWR _10779_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17455_ _13081_ _13168_ decode.regfile.registers_23\[16\] _13041_ VGND VGND VPWR
+ VPWR _13404_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14667_ decode.id_ex_pc_reg\[13\] VGND VGND VPWR VPWR _10710_ sky130_fd_sc_hd__buf_2
XFILLER_0_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16406_ decode.regfile.registers_25\[28\] _11333_ _11336_ decode.regfile.registers_24\[28\]
+ VGND VGND VPWR VPWR _12375_ sky130_fd_sc_hd__o22a_1
XFILLER_0_223_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13618_ _09977_ _09978_ memory.io_wb_reg_pc\[4\] VGND VGND VPWR VPWR _09979_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17386_ _12492_ decode.regfile.registers_29\[14\] _13303_ _13336_ _12702_ VGND VGND
+ VPWR VPWR _13337_ sky130_fd_sc_hd__o221a_1
XFILLER_0_144_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14598_ _10640_ decode.id_ex_ex_rd_reg\[0\] VGND VGND VPWR VPWR _10641_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19125_ _04349_ _04420_ _04421_ _04414_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_70_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16337_ _11396_ _12305_ _12306_ _12307_ VGND VGND VPWR VPWR _12308_ sky130_fd_sc_hd__a31o_1
X_13549_ _09914_ _09890_ _09917_ net398 VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19056_ _04205_ net190 _04233_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16268_ decode.regfile.registers_13\[25\] _11275_ _11278_ decode.regfile.registers_12\[25\]
+ VGND VGND VPWR VPWR _12240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18007_ _12494_ decode.regfile.registers_26\[30\] _13002_ _11010_ _11026_ VGND VGND
+ VPWR VPWR _03404_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_207_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15219_ _11104_ VGND VGND VPWR VPWR _11216_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16199_ decode.regfile.registers_11\[23\] _11071_ _11204_ _11187_ VGND VGND VPWR
+ VPWR _12173_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19958_ _10705_ _03599_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18909_ _03929_ _03933_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_203_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_203_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19889_ _03789_ _03790_ _03803_ _05123_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_199_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21920_ _06553_ _06543_ _06544_ _06554_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_195_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21851_ csr._mcycle_T_2\[4\] _06497_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20802_ execute.io_mem_memtoreg\[0\] _05867_ _05875_ VGND VGND VPWR VPWR _05876_
+ sky130_fd_sc_hd__and3_1
X_21782_ _06454_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24570_ net878 execute.io_target_pc\[7\] _08462_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23521_ net2178 _07890_ _07901_ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20733_ _05831_ _05808_ decode.id_ex_rs1_data_reg\[23\] _05837_ _00514_ VGND VGND
+ VPWR VPWR _00742_ sky130_fd_sc_hd__a32o_1
XFILLER_0_148_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26240_ _09446_ VGND VGND VPWR VPWR _09448_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23452_ _10670_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__buf_2
X_20664_ decode.id_ex_funct3_reg\[0\] decode.id_ex_funct3_reg\[1\] _03587_ VGND VGND
+ VPWR VPWR _05792_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_154_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22403_ fetch.bht.bhtTable_tag\[0\]\[21\] fetch.bht.bhtTable_tag\[1\]\[21\] fetch.bht.bhtTable_tag\[2\]\[21\]
+ fetch.bht.bhtTable_tag\[3\]\[21\] _06617_ _06622_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23383_ _07805_ _07806_ _07081_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__mux2_1
X_26171_ net2342 _09395_ _09399_ _09394_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_208_Left_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20595_ net2390 _05593_ _05625_ _05732_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__o32a_1
XFILLER_0_2_1281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25122_ _08789_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__clkbuf_1
X_22334_ fetch.bht.bhtTable_tag\[6\]\[10\] fetch.bht.bhtTable_tag\[7\]\[10\] _06680_
+ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22265_ fetch.bht.bhtTable_tag\[8\]\[17\] fetch.bht.bhtTable_tag\[9\]\[17\] fetch.bht.bhtTable_tag\[10\]\[17\]
+ fetch.bht.bhtTable_tag\[11\]\[17\] _06691_ _06677_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__mux4_1
X_25053_ net2774 _08710_ _08748_ _03555_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__a211oi_1
X_29930_ clknet_leaf_340_clock _02943_ VGND VGND VPWR VPWR decode.regfile.registers_21\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24004_ _08173_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__clkbuf_1
X_21216_ _10821_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__buf_2
XFILLER_0_108_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29861_ clknet_leaf_303_clock _02874_ VGND VGND VPWR VPWR decode.regfile.registers_19\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_22196_ fetch.bht.bhtTable_tag\[8\]\[5\] fetch.bht.bhtTable_tag\[9\]\[5\] fetch.bht.bhtTable_tag\[10\]\[5\]
+ fetch.bht.bhtTable_tag\[11\]\[5\] _06644_ _06730_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__mux4_1
XFILLER_0_228_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28812_ clknet_leaf_88_clock _01825_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_21147_ _06062_ _06058_ net2317 VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__and3_1
X_29792_ clknet_leaf_310_clock _02805_ VGND VGND VPWR VPWR decode.regfile.registers_17\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28743_ clknet_leaf_118_clock _01756_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25955_ _08952_ _09267_ VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__nand2_1
X_21078_ execute.csr_read_data_out_reg\[27\] _06025_ _03583_ VGND VGND VPWR VPWR _06026_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_217_Left_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20029_ decode.id_ex_imm_reg\[3\] _10747_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__o21ai_1
X_24906_ csr._mcycle_T_3\[36\] csr._mcycle_T_3\[35\] csr._mcycle_T_3\[34\] _08647_
+ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28674_ clknet_leaf_133_clock _01687_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25886_ net2506 _09226_ _09230_ _09222_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_87_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27625_ clknet_leaf_54_clock _00654_ VGND VGND VPWR VPWR execute.io_reg_pc\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24837_ _06115_ net1586 _08422_ VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27556_ clknet_leaf_52_clock _00585_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dfxtp_2
X_15570_ decode.regfile.registers_23\[6\] _11262_ _11530_ _11560_ _11335_ VGND VGND
+ VPWR VPWR _11561_ sky130_fd_sc_hd__o221a_1
X_24768_ _08062_ net1979 _08563_ VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__mux2_1
Xrebuffer90 _04396_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_1
XFILLER_0_56_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14521_ _10550_ _10554_ _10559_ _10563_ VGND VGND VPWR VPWR _10566_ sky130_fd_sc_hd__nor4_1
X_26507_ net2412 _09592_ _09601_ _09595_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__o211a_1
X_23719_ _08010_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_25_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27487_ clknet_leaf_33_clock _00516_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24699_ _08533_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29226_ clknet_leaf_106_clock _02239_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17240_ decode.regfile.registers_4\[11\] _12548_ _13145_ decode.regfile.registers_5\[11\]
+ _12614_ VGND VGND VPWR VPWR _13194_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26438_ _09420_ _09558_ VGND VGND VPWR VPWR _09562_ sky130_fd_sc_hd__nand2_1
X_14452_ net441 _10506_ _10519_ _10509_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_226_Left_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29157_ clknet_leaf_212_clock _02170_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17171_ decode.regfile.registers_22\[9\] _13100_ _13125_ _13126_ _12687_ VGND VGND
+ VPWR VPWR _13127_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26369_ _09426_ _09515_ VGND VGND VPWR VPWR _09522_ sky130_fd_sc_hd__nand2_1
X_14383_ _10042_ _10474_ VGND VGND VPWR VPWR _10480_ sky130_fd_sc_hd__nand2_1
X_28108_ clknet_leaf_82_clock net2445 VGND VGND VPWR VPWR csr.minstret\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16122_ _11942_ net2784 _12095_ _12096_ _12097_ VGND VGND VPWR VPWR _12098_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_88_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29088_ clknet_leaf_71_clock _02101_ VGND VGND VPWR VPWR csr._mcycle_T_3\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28039_ clknet_leaf_183_clock _01061_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16053_ _12020_ _12029_ _12030_ VGND VGND VPWR VPWR _12031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_1344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15004_ _11014_ VGND VGND VPWR VPWR _11015_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_55_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19812_ _04693_ _04879_ _05075_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_47_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19743_ _04974_ _04972_ _04995_ _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__a31oi_2
X_16955_ _12915_ decode.regfile.registers_25\[4\] _12506_ _12812_ VGND VGND VPWR VPWR
+ _12916_ sky130_fd_sc_hd__or4_1
XFILLER_0_224_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15906_ decode.regfile.registers_7\[15\] _11465_ _11466_ decode.regfile.registers_6\[15\]
+ _11165_ VGND VGND VPWR VPWR _11888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19674_ _04942_ _04943_ _04948_ _04951_ _04952_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__o41a_4
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16886_ decode.regfile.registers_10\[3\] _12652_ _12791_ VGND VGND VPWR VPWR _12848_
+ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_331_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_331_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_216_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15837_ decode.regfile.registers_19\[13\] _11406_ _11798_ _11820_ _11219_ VGND VGND
+ VPWR VPWR _11821_ sky130_fd_sc_hd__o221a_1
X_18625_ _03918_ _03923_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15768_ _11260_ _11751_ _11752_ _11753_ VGND VGND VPWR VPWR _11754_ sky130_fd_sc_hd__a31o_1
X_18556_ execute.csr_read_data_out_reg\[30\] _03659_ net123 _03666_ VGND VGND VPWR
+ VPWR _03855_ sky130_fd_sc_hd__o22a_1
XFILLER_0_220_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14719_ csr.io_mem_pc\[7\] csr.io_mem_pc\[8\] csr.io_mem_pc\[9\] _10761_ VGND VGND
+ VPWR VPWR _10762_ sky130_fd_sc_hd__and4_1
X_17507_ decode.regfile.registers_8\[18\] _10593_ _12549_ _12592_ _12606_ VGND VGND
+ VPWR VPWR _13454_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_190_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_346_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_346_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18487_ _03759_ _03779_ decode.id_ex_rs2_data_reg\[29\] _03747_ _03727_ VGND VGND
+ VPWR VPWR _03786_ sky130_fd_sc_hd__o221a_1
XFILLER_0_170_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15699_ _11446_ decode.regfile.registers_26\[10\] _11447_ _10981_ _11448_ VGND VGND
+ VPWR VPWR _11686_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_59_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17438_ _13381_ _13385_ _13386_ VGND VGND VPWR VPWR _13387_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_15 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_26 _08939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 _10019_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_48 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17369_ decode.regfile.registers_9\[14\] _12602_ _13310_ _13319_ VGND VGND VPWR VPWR
+ _13320_ sky130_fd_sc_hd__o22a_1
XANTENNA_59 _10795_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19108_ _04346_ _04362_ _04370_ _04387_ _04405_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__o311a_1
X_20380_ csr.io_csr_address\[11\] csr.io_csr_address\[10\] csr.io_csr_address\[9\]
+ csr.io_csr_address\[8\] VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__nand4_1
XFILLER_0_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_209_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_209_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19039_ _04324_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput100 net100 VGND VGND VPWR VPWR io_memory_address[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput111 net111 VGND VGND VPWR VPWR io_memory_address[1] sky130_fd_sc_hd__clkbuf_4
Xoutput122 net122 VGND VGND VPWR VPWR io_memory_address[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22050_ _06644_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__buf_4
XFILLER_0_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput133 net133 VGND VGND VPWR VPWR io_memory_size[0] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput144 net144 VGND VGND VPWR VPWR io_memory_write_data[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput155 net155 VGND VGND VPWR VPWR io_memory_write_data[27] sky130_fd_sc_hd__clkbuf_4
Xoutput166 net166 VGND VGND VPWR VPWR io_memory_write_data[8] sky130_fd_sc_hd__clkbuf_4
X_21001_ execute.io_reg_pc\[25\] _05977_ _05973_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_6 _00932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_197_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25740_ net2706 _09139_ _09146_ _09142_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__o211a_1
X_22952_ fetch.bht.bhtTable_target_pc\[12\]\[4\] fetch.bht.bhtTable_target_pc\[13\]\[4\]
+ fetch.bht.bhtTable_target_pc\[14\]\[4\] fetch.bht.bhtTable_target_pc\[15\]\[4\]
+ _07123_ _07101_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21903_ csr.io_mret_vector\[20\] _10795_ _06539_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25671_ _08970_ _09067_ VGND VGND VPWR VPWR _09106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_222_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22883_ _07338_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27410_ clknet_leaf_10_clock _00439_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[19\]
+ sky130_fd_sc_hd__dfxtp_4
X_24622_ _08493_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28390_ clknet_leaf_143_clock _01403_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_4
X_21834_ _06492_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_214_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27341_ clknet_leaf_45_clock _00370_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_24553_ _08113_ net1756 _09902_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21765_ _06445_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23504_ _04459_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_1112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27272_ clknet_leaf_12_clock _00301_ VGND VGND VPWR VPWR decode.regfile.registers_30\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_20716_ _05818_ decode.id_ex_rs1_data_reg\[17\] _05710_ VGND VGND VPWR VPWR _05827_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_175_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24484_ _08387_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__clkbuf_8
X_21696_ _06320_ _06365_ _06397_ _06398_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_163_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29011_ clknet_leaf_139_clock _02024_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26223_ net2652 _09419_ _09435_ _09418_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23435_ net29 _07846_ _07852_ _07851_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20647_ _05526_ _05536_ _05618_ csr._csr_read_data_T_8\[29\] _05777_ VGND VGND VPWR
+ VPWR _05778_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26154_ _10007_ VGND VGND VPWR VPWR _09387_ sky130_fd_sc_hd__buf_4
X_23366_ fetch.bht.bhtTable_target_pc\[8\]\[28\] fetch.bht.bhtTable_target_pc\[9\]\[28\]
+ fetch.bht.bhtTable_target_pc\[10\]\[28\] fetch.bht.bhtTable_target_pc\[11\]\[28\]
+ _07119_ _07071_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__mux4_1
X_20578_ _05541_ csr.io_mret_vector\[19\] _05602_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_115_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25105_ _06122_ net1603 _08778_ VGND VGND VPWR VPWR _08781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22317_ _06909_ _06685_ _06631_ _06911_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__a211o_1
X_26085_ _09263_ VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_186_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23297_ execute.io_target_pc\[23\] _07090_ _06041_ _06038_ VGND VGND VPWR VPWR _07727_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_186_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25036_ csr.mcycle\[16\] csr.mcycle\[15\] _08733_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29913_ clknet_leaf_305_clock _02926_ VGND VGND VPWR VPWR decode.regfile.registers_20\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_22248_ fetch.bht.bhtTable_tag\[8\]\[19\] fetch.bht.bhtTable_tag\[9\]\[19\] fetch.bht.bhtTable_tag\[10\]\[19\]
+ fetch.bht.bhtTable_tag\[11\]\[19\] _06616_ _06621_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__mux4_2
X_22179_ fetch.bht.bhtTable_tag\[2\]\[25\] fetch.bht.bhtTable_tag\[3\]\[25\] _06619_
+ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__mux2_1
X_29844_ clknet_leaf_299_clock _02857_ VGND VGND VPWR VPWR decode.regfile.registers_18\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29775_ clknet_leaf_294_clock _02788_ VGND VGND VPWR VPWR decode.regfile.registers_16\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_26987_ _10141_ _09838_ VGND VGND VPWR VPWR _09877_ sky130_fd_sc_hd__nand2_1
XFILLER_0_218_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_145_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16740_ _12704_ VGND VGND VPWR VPWR _12705_ sky130_fd_sc_hd__clkbuf_4
X_28726_ clknet_leaf_127_clock _01739_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13952_ _10102_ _10223_ VGND VGND VPWR VPWR _10230_ sky130_fd_sc_hd__nand2_1
X_25938_ net2080 _09256_ _09260_ _09250_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28657_ clknet_leaf_104_clock _01670_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_16671_ net215 VGND VGND VPWR VPWR _12636_ sky130_fd_sc_hd__clkbuf_8
X_13883_ _10122_ _10177_ VGND VGND VPWR VPWR _10189_ sky130_fd_sc_hd__nand2_1
X_25869_ net1090 _09213_ _09220_ _09209_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15622_ _10959_ decode.regfile.registers_26\[8\] _11447_ _11348_ _10993_ VGND VGND
+ VPWR VPWR _11611_ sky130_fd_sc_hd__o2111a_1
X_18410_ _03708_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__buf_8
X_27608_ clknet_leaf_158_clock _00637_ VGND VGND VPWR VPWR execute.io_target_pc\[17\]
+ sky130_fd_sc_hd__dfxtp_4
X_19390_ _03639_ _04345_ _04306_ _04679_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__or4_1
X_28588_ clknet_leaf_101_clock _01601_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_205 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_216 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_227 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18341_ execute.io_mem_rd\[3\] VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__inv_2
X_27539_ clknet_leaf_45_clock net357 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_2
X_15553_ _11146_ _11542_ _11543_ VGND VGND VPWR VPWR _11544_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_104_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_238 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_249 net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14504_ fetch.btb.btbTable\[4\]\[1\] fetch.btb.btbTable\[5\]\[1\] fetch.btb.btbTable\[6\]\[1\]
+ fetch.btb.btbTable\[7\]\[1\] _09891_ _09888_ VGND VGND VPWR VPWR _10549_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_13_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _03600_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15484_ _10955_ _11215_ _11216_ _11476_ VGND VGND VPWR VPWR _11477_ sky130_fd_sc_hd__o31a_1
XFILLER_0_204_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1088 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17223_ _12701_ decode.regfile.registers_28\[10\] _13093_ VGND VGND VPWR VPWR _13178_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29209_ clknet_leaf_162_clock _02222_ VGND VGND VPWR VPWR fetch.btb.btbTable\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14435_ net539 _10506_ _10510_ _10509_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput13 io_fetch_data[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput24 net375 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17154_ _13107_ _13108_ _13109_ VGND VGND VPWR VPWR _13110_ sky130_fd_sc_hd__a21o_1
XFILLER_0_226_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput35 io_memory_read_data[10] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
X_14366_ net536 _10463_ _10470_ _10468_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__o211a_1
Xinput46 io_memory_read_data[20] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
Xinput57 io_memory_read_data[30] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
X_16105_ decode.regfile.registers_19\[20\] _11049_ _11215_ _11217_ _11454_ VGND VGND
+ VPWR VPWR _12082_ sky130_fd_sc_hd__o41a_1
XFILLER_0_220_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold808 fetch.bht.bhtTable_target_pc\[12\]\[20\] VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold819 fetch.bht.bhtTable_tag\[10\]\[13\] VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__dlygate4sd3_1
X_17085_ _10927_ decode.regfile.registers_24\[7\] _10933_ _12759_ _12862_ VGND VGND
+ VPWR VPWR _13043_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14297_ net541 _10419_ _10430_ _10427_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16036_ _11761_ net469 _11983_ _12014_ _11760_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__o221a_1
XFILLER_0_161_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2209 csr._mcycle_T_2\[8\] VGND VGND VPWR VPWR net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1508 fetch.bht.bhtTable_target_pc\[14\]\[23\] VGND VGND VPWR VPWR net1735 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17987_ decode.regfile.registers_4\[30\] _12548_ _13145_ decode.regfile.registers_5\[30\]
+ _12625_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__a221oi_1
Xhold1519 fetch.bht.bhtTable_tag\[5\]\[6\] VGND VGND VPWR VPWR net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_270_clock clknet_5_20__leaf_clock VGND VGND VPWR VPWR clknet_leaf_270_clock
+ sky130_fd_sc_hd__clkbuf_8
X_19726_ _04408_ _04992_ _04993_ _04445_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16938_ decode.regfile.registers_15\[4\] _12874_ _12875_ _12898_ VGND VGND VPWR VPWR
+ _12899_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_205_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19657_ _04199_ _04200_ _03937_ _03903_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__o31a_1
X_16869_ decode.regfile.registers_1\[3\] decode.regfile.registers_0\[3\] _12631_ VGND
+ VGND VPWR VPWR _12831_ sky130_fd_sc_hd__mux2_1
X_18608_ _03751_ net304 net240 _03784_ decode.id_ex_rs2_data_reg\[17\] VGND VGND VPWR
+ VPWR _03907_ sky130_fd_sc_hd__a311o_4
XFILLER_0_149_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_285_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_285_clock
+ sky130_fd_sc_hd__clkbuf_8
X_19588_ _04496_ _04862_ _04863_ _04869_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18539_ _03709_ decode.id_ex_imm_reg\[25\] _03837_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21550_ _06283_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_151_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20501_ _05541_ csr.io_mret_vector\[9\] _05602_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21481_ _06257_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23220_ execute.io_target_pc\[19\] _10757_ _10970_ _06037_ VGND VGND VPWR VPWR _07654_
+ sky130_fd_sc_hd__a211o_1
X_20432_ csr.io_mret_vector\[2\] _05580_ _05581_ net1913 VGND VGND VPWR VPWR _05590_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23151_ net73 _07582_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__nand2_1
X_20363_ _05525_ _03721_ net293 VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__and3_4
XFILLER_0_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_223_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_223_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_228_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22102_ _06693_ _06695_ _06696_ _06673_ _06641_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_228_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23082_ _07522_ _07523_ _07082_ VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20294_ _05418_ _05331_ _05470_ _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_149_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22033_ _06627_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__buf_4
XFILLER_0_140_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26910_ _09438_ _09794_ VGND VGND VPWR VPWR _09833_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_181_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27890_ clknet_leaf_23_clock _00919_ VGND VGND VPWR VPWR csr._mcycle_T_2\[11\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_181_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26841_ net331 _10149_ _10196_ _09935_ VGND VGND VPWR VPWR _09793_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_71_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_238_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_238_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_177_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29560_ clknet_leaf_313_clock _02573_ VGND VGND VPWR VPWR decode.regfile.registers_9\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26772_ _09450_ _09753_ VGND VGND VPWR VPWR _09755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_215_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23984_ net978 execute.io_target_pc\[13\] _08153_ VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28511_ clknet_leaf_196_clock _01524_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25723_ _08945_ _09136_ VGND VGND VPWR VPWR _09137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_225_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22935_ fetch.bht.bhtTable_target_pc\[12\]\[3\] fetch.bht.bhtTable_target_pc\[13\]\[3\]
+ fetch.bht.bhtTable_target_pc\[14\]\[3\] fetch.bht.bhtTable_target_pc\[15\]\[3\]
+ _07384_ _07113_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__mux4_1
X_29491_ clknet_leaf_264_clock _02504_ VGND VGND VPWR VPWR decode.regfile.registers_7\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28442_ clknet_leaf_54_clock _01455_ VGND VGND VPWR VPWR decode.io_id_pc\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_140_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25654_ _08954_ _09092_ VGND VGND VPWR VPWR _09097_ sky130_fd_sc_hd__nand2_1
X_22866_ _07329_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_179_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24605_ net1440 execute.io_target_pc\[24\] _09897_ VGND VGND VPWR VPWR _08485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28373_ clknet_leaf_199_clock _01386_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21817_ _06038_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__buf_4
XFILLER_0_196_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25585_ _08960_ _09049_ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__nand2_1
X_22797_ _07293_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27324_ clknet_leaf_25_clock _00353_ VGND VGND VPWR VPWR decode.id_ex_funct3_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_24536_ _08449_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21748_ _06436_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_117_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_159_Left_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27255_ clknet_leaf_9_clock _00284_ VGND VGND VPWR VPWR decode.regfile.registers_30\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_24467_ _08413_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21679_ net1093 _06329_ csr.minstret\[22\] VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26206_ net193 VGND VGND VPWR VPWR _09424_ sky130_fd_sc_hd__buf_4
X_14220_ _10008_ _10377_ VGND VGND VPWR VPWR _10386_ sky130_fd_sc_hd__nand2_1
X_23418_ _06633_ _07835_ _07837_ _07839_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__o22a_1
X_27186_ clknet_leaf_352_clock _00215_ VGND VGND VPWR VPWR decode.regfile.registers_28\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24398_ _08376_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14151_ _10331_ VGND VGND VPWR VPWR _10346_ sky130_fd_sc_hd__buf_2
X_26137_ _08982_ _09374_ VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__nand2_1
X_23349_ net85 _07706_ _07707_ _07775_ _07705_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__o311a_1
XFILLER_0_132_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14082_ net1113 _10302_ _10306_ _10304_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__o211a_1
X_26068_ _08914_ _09330_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__nand2_1
X_25019_ csr._mcycle_T_2\[11\] _08712_ _08725_ csr.mcycle\[11\] VGND VGND VPWR VPWR
+ _08726_ sky130_fd_sc_hd__a211o_1
X_17910_ _12530_ _12616_ _12557_ decode.regfile.registers_0\[28\] VGND VGND VPWR VPWR
+ _03309_ sky130_fd_sc_hd__a31o_1
X_18890_ _03888_ _03893_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Left_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17841_ decode.regfile.registers_12\[26\] _12542_ _12723_ _03229_ _03241_ VGND VGND
+ VPWR VPWR _03242_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_7_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29827_ clknet_leaf_307_clock _02840_ VGND VGND VPWR VPWR decode.regfile.registers_18\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14984_ _10667_ _10950_ _10952_ _10969_ VGND VGND VPWR VPWR _11002_ sky130_fd_sc_hd__nor4_1
XFILLER_0_22_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17772_ _11014_ _10936_ decode.regfile.registers_23\[24\] _12995_ VGND VGND VPWR
+ VPWR _03175_ sky130_fd_sc_hd__or4_1
X_29758_ clknet_leaf_310_clock _02771_ VGND VGND VPWR VPWR decode.regfile.registers_16\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19511_ _04302_ _04794_ _04795_ _04425_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_57_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28709_ clknet_leaf_136_clock _01722_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13935_ net1887 _10213_ _10220_ _10219_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__o211a_1
X_16723_ decode.regfile.registers_22\[0\] _12528_ _12687_ VGND VGND VPWR VPWR _12688_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29689_ clknet_leaf_289_clock _02702_ VGND VGND VPWR VPWR decode.regfile.registers_13\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19442_ _04511_ _04509_ _04515_ _04633_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_18_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16654_ _12522_ _12530_ _12616_ VGND VGND VPWR VPWR _12619_ sky130_fd_sc_hd__and3_2
XFILLER_0_201_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13866_ net2414 _10167_ _10179_ _10175_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15605_ decode.regfile.registers_17\[7\] _11357_ _11594_ VGND VGND VPWR VPWR _11595_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16585_ _12549_ VGND VGND VPWR VPWR _12550_ sky130_fd_sc_hd__clkbuf_4
X_19373_ _04635_ _04142_ _04143_ _04637_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__or4_4
XFILLER_0_215_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13797_ _10060_ memory.io_wb_aluresult\[29\] _10004_ memory.io_wb_readdata\[29\]
+ _10005_ VGND VGND VPWR VPWR _10133_ sky130_fd_sc_hd__a221o_1
X_15536_ _11344_ net582 _11492_ _11527_ _11249_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__o221a_1
X_18324_ decode.id_ex_rs2_data_reg\[27\] _03627_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18255_ _03587_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15467_ decode.regfile.registers_2\[4\] _11190_ _11148_ _11151_ _11459_ VGND VGND
+ VPWR VPWR _11460_ sky130_fd_sc_hd__o311a_1
XFILLER_0_127_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17206_ decode.regfile.registers_17\[10\] _12579_ _12565_ _13160_ VGND VGND VPWR
+ VPWR _13161_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14418_ net557 _10490_ _10499_ _10494_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__o211a_1
X_18186_ _10943_ decode.control.io_funct3\[0\] VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15398_ decode.regfile.registers_23\[2\] _11086_ _11353_ _11392_ _11335_ VGND VGND
+ VPWR VPWR _11393_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17137_ _12701_ decode.regfile.registers_28\[8\] _13093_ VGND VGND VPWR VPWR _13094_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14349_ net602 _10420_ _10459_ _10453_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__o211a_1
Xhold605 fetch.bht.bhtTable_target_pc\[8\]\[25\] VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 csr.minstret\[23\] VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_2_1_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_1_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold627 fetch.bht.bhtTable_tag\[1\]\[21\] VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 fetch.bht.bhtTable_target_pc\[2\]\[14\] VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold649 decode.regfile.registers_1\[13\] VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17068_ _13023_ _13024_ _13025_ VGND VGND VPWR VPWR _13026_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16019_ decode.regfile.registers_8\[18\] _11280_ _11175_ _11131_ VGND VGND VPWR VPWR
+ _11998_ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2006 fetch.bht.bhtTable_target_pc\[14\]\[30\] VGND VGND VPWR VPWR net2233 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2017 decode.regfile.registers_27\[10\] VGND VGND VPWR VPWR net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2028 net97 VGND VGND VPWR VPWR net2255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2039 decode.regfile.registers_7\[18\] VGND VGND VPWR VPWR net2266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1305 fetch.bht.bhtTable_target_pc\[7\]\[0\] VGND VGND VPWR VPWR net1532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1316 decode.regfile.registers_21\[8\] VGND VGND VPWR VPWR net1543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 fetch.bht.bhtTable_tag\[5\]\[0\] VGND VGND VPWR VPWR net1554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1338 fetch.bht.bhtTable_tag\[15\]\[11\] VGND VGND VPWR VPWR net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 fetch.bht.bhtTable_target_pc\[13\]\[20\] VGND VGND VPWR VPWR net1576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19709_ _04290_ _04594_ _04879_ _04985_ _04595_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__a32o_1
XFILLER_0_174_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20981_ _03582_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22720_ _03524_ _03539_ _07250_ _03458_ decode.control.io_opcode\[5\] VGND VGND VPWR
+ VPWR _07251_ sky130_fd_sc_hd__o311a_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22651_ net2662 _07208_ _07211_ _07164_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_217_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21602_ _06320_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__clkbuf_4
X_25370_ _10014_ VGND VGND VPWR VPWR _08922_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22582_ csr._minstret_T_3\[41\] _07160_ net2617 VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24321_ _08083_ net1658 _08334_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21533_ _06286_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27040_ clknet_leaf_342_clock _00069_ VGND VGND VPWR VPWR decode.regfile.registers_23\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24252_ _08301_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21464_ net1 _10673_ _10911_ _09957_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__o31a_1
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_162_clock clknet_5_24__leaf_clock VGND VGND VPWR VPWR clknet_leaf_162_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23203_ fetch.bht.bhtTable_target_pc\[0\]\[18\] fetch.bht.bhtTable_target_pc\[1\]\[18\]
+ fetch.bht.bhtTable_target_pc\[2\]\[18\] fetch.bht.bhtTable_target_pc\[3\]\[18\]
+ _07098_ _07113_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20415_ _05573_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24183_ _08265_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__clkbuf_1
X_21395_ _06143_ net2182 _06210_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23134_ _07345_ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20346_ _05508_ decode.id_ex_pc_reg\[30\] _05411_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_73_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28991_ clknet_leaf_182_clock _02004_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23065_ _07506_ _07507_ _07406_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__mux2_1
X_27942_ clknet_leaf_165_clock _00964_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20277_ _10694_ _05452_ _10710_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_177_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_177_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22016_ net1251 _06573_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__or2_1
XFILLER_0_216_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27873_ clknet_leaf_327_clock _00902_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2540 decode.io_id_pc\[0\] VGND VGND VPWR VPWR net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2551 net76 VGND VGND VPWR VPWR net2778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29612_ clknet_leaf_276_clock _02625_ VGND VGND VPWR VPWR decode.regfile.registers_11\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1098 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26824_ net1991 _09779_ _09783_ _09784_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__o211a_1
Xhold2562 csr._mcycle_T_2\[14\] VGND VGND VPWR VPWR net2789 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2573 csr._mcycle_T_2\[31\] VGND VGND VPWR VPWR net2800 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_100_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_100_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_32_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1850 fetch.bht.bhtTable_tag\[0\]\[11\] VGND VGND VPWR VPWR net2077 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1861 decode.regfile.registers_20\[17\] VGND VGND VPWR VPWR net2088 sky130_fd_sc_hd__dlygate4sd3_1
X_26755_ net2367 _09736_ _09744_ _09743_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__o211a_1
X_29543_ clknet_leaf_273_clock _02556_ VGND VGND VPWR VPWR decode.regfile.registers_9\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_23967_ _08154_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__clkbuf_1
Xhold1872 decode.regfile.registers_13\[27\] VGND VGND VPWR VPWR net2099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1883 decode.regfile.registers_29\[4\] VGND VGND VPWR VPWR net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1894 fetch.bht.bhtTable_tag\[9\]\[22\] VGND VGND VPWR VPWR net2121 sky130_fd_sc_hd__dlygate4sd3_1
X_13720_ memory.csr_read_data_out_reg\[17\] _09986_ _10066_ _10067_ VGND VGND VPWR
+ VPWR _10068_ sky130_fd_sc_hd__a2bb2o_4
X_25706_ _08931_ _09122_ VGND VGND VPWR VPWR _09127_ sky130_fd_sc_hd__nand2_1
X_22918_ fetch.bht.bhtTable_target_pc\[4\]\[2\] fetch.bht.bhtTable_target_pc\[5\]\[2\]
+ fetch.bht.bhtTable_target_pc\[6\]\[2\] fetch.bht.bhtTable_target_pc\[7\]\[2\] _07107_
+ _07071_ VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__mux4_1
X_26686_ net2234 _09692_ _09704_ _09702_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__o211a_1
X_29474_ clknet_leaf_253_clock _02487_ VGND VGND VPWR VPWR decode.regfile.registers_7\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_23898_ _08118_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25637_ net2426 _09082_ _09086_ _09087_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__o211a_1
X_28425_ clknet_leaf_246_clock _01438_ VGND VGND VPWR VPWR decode.immGen._imm_T_24\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_13651_ _10008_ _09951_ VGND VGND VPWR VPWR _10009_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22849_ _07320_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_115_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_115_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_195_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28356_ clknet_leaf_184_clock _01369_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16370_ _10959_ decode.regfile.registers_26\[27\] _11349_ _10980_ _11347_ VGND VGND
+ VPWR VPWR _12340_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_183_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25568_ net755 _09039_ _09047_ _09046_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__o211a_1
X_13582_ _09940_ _09939_ VGND VGND VPWR VPWR _09947_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_155_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15321_ _11181_ _11312_ _11316_ VGND VGND VPWR VPWR _11317_ sky130_fd_sc_hd__o21ai_1
X_27307_ clknet_leaf_14_clock _00336_ VGND VGND VPWR VPWR decode.regfile.registers_31\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24519_ _08078_ net2151 _08439_ VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28287_ clknet_leaf_85_clock _01309_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25499_ net2601 _08995_ _09007_ _09004_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18040_ decode.regfile.registers_22\[31\] _12527_ _03434_ _03435_ _12686_ VGND VGND
+ VPWR VPWR _03436_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27238_ clknet_leaf_364_clock _00267_ VGND VGND VPWR VPWR decode.regfile.registers_29\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_15252_ _11248_ VGND VGND VPWR VPWR _11249_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14203_ _10375_ VGND VGND VPWR VPWR _10376_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27169_ clknet_leaf_362_clock _00198_ VGND VGND VPWR VPWR decode.regfile.registers_27\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_15183_ _11179_ VGND VGND VPWR VPWR _11180_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14134_ net482 _10332_ _10336_ _10328_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19991_ _10697_ _05214_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_176_Left_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18942_ _03635_ _03634_ _03633_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__and3b_1
X_14065_ net1005 _10287_ _10296_ _10291_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18873_ _04070_ _04073_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__nand2_4
XFILLER_0_197_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17824_ _13451_ net496 _13492_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17755_ decode.regfile.registers_4\[24\] _10609_ _12882_ _12614_ VGND VGND VPWR VPWR
+ _03158_ sky130_fd_sc_hd__or4_1
X_14967_ _10991_ VGND VGND VPWR VPWR _10992_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16706_ _11021_ _12491_ _12667_ decode.regfile.registers_14\[0\] _12670_ VGND VGND
+ VPWR VPWR _12671_ sky130_fd_sc_hd__o32a_1
XFILLER_0_57_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13918_ _10015_ _10210_ VGND VGND VPWR VPWR _10211_ sky130_fd_sc_hd__nand2_1
X_17686_ _12498_ _12489_ _12510_ decode.regfile.registers_12\[22\] _12590_ VGND VGND
+ VPWR VPWR _03091_ sky130_fd_sc_hd__o32a_1
X_14898_ _10933_ _10577_ _10673_ _10911_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__nor4_1
XFILLER_0_162_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_185_Left_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19425_ _04710_ _04241_ _04712_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__and3_1
X_13849_ _10042_ _10164_ VGND VGND VPWR VPWR _10170_ sky130_fd_sc_hd__nand2_1
X_16637_ _12601_ VGND VGND VPWR VPWR _12602_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19356_ _04254_ _04126_ _04327_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__o21a_1
X_16568_ _12532_ VGND VGND VPWR VPWR _12533_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18307_ decode.id_ex_rs2_data_reg\[19\] _03616_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15519_ _11508_ _11510_ VGND VGND VPWR VPWR _11511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16499_ _11289_ _12463_ _12464_ VGND VGND VPWR VPWR _12465_ sky130_fd_sc_hd__o21ai_1
X_19287_ _04075_ _04172_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_212_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18238_ _03569_ _03570_ _03571_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_212_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18169_ _03512_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold402 decode.regfile.registers_28\[9\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 io_fetch_data[11] VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_225_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_194_Left_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20200_ _00576_ _05227_ _05398_ _05267_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21180_ _06074_ _06082_ net1476 VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__and3_1
Xhold424 decode.regfile.registers_20\[8\] VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_94_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_94_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold435 csr._csr_read_data_T_9\[3\] VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold446 decode.regfile.registers_3\[9\] VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold457 fetch.bht.bhtTable_valid\[11\] VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20131_ decode.id_ex_imm_reg\[19\] decode.id_ex_pc_reg\[19\] VGND VGND VPWR VPWR
+ _05339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold468 decode.regfile.registers_7\[14\] VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold479 decode.regfile.registers_28\[8\] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap198 _10086_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_221_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20062_ decode.id_ex_imm_reg\[8\] decode.id_ex_pc_reg\[8\] _05279_ VGND VGND VPWR
+ VPWR _05280_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1102 fetch.bht.bhtTable_target_pc\[14\]\[21\] VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 fetch.bht.bhtTable_tag\[3\]\[22\] VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__dlygate4sd3_1
X_24870_ _06149_ net1849 _08388_ VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1124 fetch.bht.bhtTable_target_pc\[9\]\[22\] VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 fetch.bht.bhtTable_tag\[10\]\[15\] VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_12__f_clock clknet_2_1_0_clock VGND VGND VPWR VPWR clknet_5_12__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
Xhold1146 fetch.bht.bhtTable_tag\[5\]\[25\] VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__dlygate4sd3_1
X_23821_ execute.io_target_pc\[9\] VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__buf_2
XFILLER_0_174_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1157 net74 VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1168 fetch.bht.bhtTable_target_pc\[11\]\[0\] VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1179 fetch.bht.bhtTable_target_pc\[9\]\[7\] VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26540_ _10149_ _10196_ _03672_ VGND VGND VPWR VPWR _09620_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_219_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23752_ _08027_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_219_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_32_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20964_ execute.io_reg_pc\[8\] _05915_ _05961_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22703_ net2402 _07235_ _07240_ _07234_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__o211a_1
X_26471_ _09566_ VGND VGND VPWR VPWR _09582_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_66_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23683_ _07990_ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ _05925_ _05921_ net64 VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28210_ clknet_leaf_61_clock net1779 VGND VGND VPWR VPWR csr.mscratch\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25422_ _08958_ _08946_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29190_ clknet_leaf_239_clock _02203_ VGND VGND VPWR VPWR fetch.btb.btbTable\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_22634_ _03579_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__buf_4
XFILLER_0_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28141_ clknet_leaf_210_clock _01163_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25353_ _08910_ _08907_ VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_47_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_47_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22565_ csr._minstret_T_3\[39\] csr._minstret_T_3\[35\] csr._minstret_T_3\[34\] VGND
+ VGND VPWR VPWR _07151_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24304_ _08066_ net1980 _08323_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__mux2_1
X_21516_ _06145_ net2060 _06274_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__mux2_1
X_28072_ clknet_leaf_235_clock _01094_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25284_ _08872_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22496_ _07090_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27023_ clknet_leaf_331_clock _00052_ VGND VGND VPWR VPWR decode.regfile.registers_23\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_24235_ _08292_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21447_ _06138_ net1674 _06230_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24166_ _08060_ net1616 _08255_ VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21378_ _06126_ net1553 _06199_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23117_ _07122_ _07556_ _07127_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__o21ai_1
X_20329_ _05378_ _05412_ _03517_ _05498_ _03551_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_92_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24097_ _06426_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__clkbuf_8
X_28974_ clknet_leaf_110_clock _01987_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold980 _01239_ VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold991 fetch.bht.bhtTable_tag\[4\]\[15\] VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23048_ fetch.bht.bhtTable_target_pc\[0\]\[9\] fetch.bht.bhtTable_target_pc\[1\]\[9\]
+ fetch.bht.bhtTable_target_pc\[2\]\[9\] fetch.bht.bhtTable_target_pc\[3\]\[9\] _07108_
+ _07125_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_34_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27925_ clknet_leaf_34_clock _00954_ VGND VGND VPWR VPWR execute.io_mem_rd\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_229_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ _11070_ _11167_ decode.regfile.registers_10\[14\] _11381_ VGND VGND VPWR
+ VPWR _11853_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_30_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27856_ clknet_leaf_317_clock _00885_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2370 decode.regfile.registers_20\[29\] VGND VGND VPWR VPWR net2597 sky130_fd_sc_hd__dlygate4sd3_1
X_14821_ decode.id_ex_pc_reg\[22\] VGND VGND VPWR VPWR _10864_ sky130_fd_sc_hd__clkbuf_4
Xhold2381 csr.minstret\[2\] VGND VGND VPWR VPWR net2608 sky130_fd_sc_hd__dlygate4sd3_1
X_26807_ net663 _09766_ _09774_ _09771_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2392 decode.regfile.registers_19\[26\] VGND VGND VPWR VPWR net2619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24999_ csr._mcycle_T_2\[4\] _08712_ _08709_ csr.mcycle\[3\] csr.mcycle\[4\] VGND
+ VGND VPWR VPWR _08713_ sky130_fd_sc_hd__a221oi_1
X_27787_ clknet_leaf_334_clock _00816_ VGND VGND VPWR VPWR memory.io_wb_readdata\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1680 fetch.bht.bhtTable_target_pc\[6\]\[1\] VGND VGND VPWR VPWR net1907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14752_ csr.io_mem_pc\[20\] VGND VGND VPWR VPWR _10795_ sky130_fd_sc_hd__buf_4
Xhold1691 execute.csr_write_address_out_reg\[8\] VGND VGND VPWR VPWR net1918 sky130_fd_sc_hd__dlygate4sd3_1
X_17540_ _12506_ VGND VGND VPWR VPWR _13487_ sky130_fd_sc_hd__clkbuf_2
X_29526_ clknet_leaf_266_clock _02539_ VGND VGND VPWR VPWR decode.regfile.registers_8\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_26738_ _09415_ _09733_ VGND VGND VPWR VPWR _09735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13703_ _10053_ _10016_ VGND VGND VPWR VPWR _10054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17471_ decode.regfile.registers_15\[17\] _12555_ _10619_ _12589_ _13031_ VGND VGND
+ VPWR VPWR _13419_ sky130_fd_sc_hd__a41o_1
X_14683_ _10725_ execute.io_target_pc\[25\] _10721_ execute.io_target_pc\[10\] VGND
+ VGND VPWR VPWR _10726_ sky130_fd_sc_hd__o2bb2a_1
X_26669_ _09424_ _09689_ VGND VGND VPWR VPWR _09695_ sky130_fd_sc_hd__nand2_1
X_29457_ clknet_leaf_260_clock _02470_ VGND VGND VPWR VPWR decode.regfile.registers_6\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19210_ _04245_ _04503_ _04505_ _04009_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28408_ clknet_leaf_113_clock _01421_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_4
X_16422_ decode.regfile.registers_2\[29\] _11503_ _11148_ _11152_ _12389_ VGND VGND
+ VPWR VPWR _12390_ sky130_fd_sc_hd__o311a_1
X_13634_ _09993_ _09951_ VGND VGND VPWR VPWR _09994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29388_ clknet_leaf_259_clock _02401_ VGND VGND VPWR VPWR decode.regfile.registers_4\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19141_ _03635_ _03634_ _04056_ _03633_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__and4b_1
XFILLER_0_55_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16353_ _11289_ _12321_ _12322_ VGND VGND VPWR VPWR _12323_ sky130_fd_sc_hd__o21ai_2
X_28339_ clknet_leaf_206_clock _01352_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13565_ net331 VGND VGND VPWR VPWR _09930_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_60_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_229_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15304_ _11153_ VGND VGND VPWR VPWR _11300_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_212_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19072_ _04369_ _04357_ _04291_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16284_ _10649_ _10625_ _11052_ _12240_ _12255_ VGND VGND VPWR VPWR _12256_ sky130_fd_sc_hd__o32a_1
XFILLER_0_212_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15235_ _11231_ VGND VGND VPWR VPWR _11232_ sky130_fd_sc_hd__clkbuf_4
X_18023_ decode.regfile.registers_8\[31\] _12892_ _03410_ _03418_ VGND VGND VPWR VPWR
+ _03419_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_81_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15166_ decode.regfile.registers_5\[0\] _10638_ _11139_ _11161_ _11162_ VGND VGND
+ VPWR VPWR _11163_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14117_ net2717 _10315_ _10325_ _10317_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_58_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19974_ _10682_ _05217_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15097_ _10652_ VGND VGND VPWR VPWR _11094_ sky130_fd_sc_hd__clkbuf_4
X_14048_ _09930_ _10195_ _09932_ _09933_ VGND VGND VPWR VPWR _10285_ sky130_fd_sc_hd__and4b_1
X_18925_ _03867_ _03882_ _03965_ _04223_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__o31a_1
XFILLER_0_181_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18856_ _04153_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__and2_2
XFILLER_0_94_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17807_ decode.regfile.registers_16\[25\] _12576_ _12719_ _03208_ VGND VGND VPWR
+ VPWR _03209_ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18787_ _04081_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__xnor2_1
X_15999_ _11679_ decode.regfile.registers_27\[17\] _11869_ VGND VGND VPWR VPWR _11979_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_206_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17738_ _12968_ _03139_ _03140_ _03141_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__a31o_1
XFILLER_0_221_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17669_ _13451_ net450 _13492_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__o21a_1
XFILLER_0_175_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19408_ _04409_ _04413_ net311 VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_214_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20680_ decode.id_ex_funct3_reg\[1\] VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19339_ _04546_ _04303_ _04626_ _04630_ _04515_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__o311a_1
XFILLER_0_70_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22350_ fetch.bht.bhtTable_tag\[0\]\[14\] fetch.bht.bhtTable_tag\[1\]\[14\] fetch.bht.bhtTable_tag\[2\]\[14\]
+ fetch.bht.bhtTable_tag\[3\]\[14\] _06616_ _06621_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21301_ _06160_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__clkbuf_1
X_22281_ _06632_ _06871_ _06873_ _06875_ _06636_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24020_ _08181_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21232_ net1879 _06113_ _09912_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold210 decode.control.io_funct7\[0\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold221 execute.csr_write_address_out_reg\[11\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 decode.regfile.registers_1\[23\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 decode.control.io_funct7\[6\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 decode.regfile.registers_23\[10\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold265 decode.regfile.registers_23\[9\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
X_21163_ _06074_ _06070_ execute.csr_write_data_out_reg\[25\] VGND VGND VPWR VPWR
+ _06076_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_165_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold276 decode.regfile.registers_19\[10\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold287 decode.regfile.registers_31\[10\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__buf_1
XFILLER_0_111_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20114_ decode.id_ex_imm_reg\[15\] _10681_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__o21ai_1
Xhold298 _08658_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21094_ _10019_ _06035_ _06025_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__and3_1
X_25971_ net2350 _09270_ _09279_ _09277_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20045_ _05262_ _05265_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__xor2_1
X_24922_ csr._mcycle_T_3\[42\] csr._mcycle_T_3\[41\] _08659_ VGND VGND VPWR VPWR _08662_
+ sky130_fd_sc_hd__and3_1
X_27710_ clknet_leaf_20_clock _00739_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_28690_ clknet_leaf_107_clock _01703_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24853_ _08614_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__clkbuf_1
X_27641_ clknet_leaf_155_clock _00670_ VGND VGND VPWR VPWR execute.io_reg_pc\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23804_ _08056_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_124_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27572_ clknet_leaf_161_clock _00601_ VGND VGND VPWR VPWR csr.io_mem_pc\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_124_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24784_ _08578_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_105 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21996_ csr._mcycle_T_2\[20\] _06600_ _06602_ _06592_ VGND VGND VPWR VPWR _01240_
+ sky130_fd_sc_hd__o211a_1
XANTENNA_116 _04981_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29311_ clknet_leaf_244_clock _02324_ VGND VGND VPWR VPWR decode.regfile.registers_2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_26523_ _09428_ _09602_ VGND VGND VPWR VPWR _09611_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_127 _10631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23735_ net1326 _10777_ _08014_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_138 _12551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20947_ net2752 _05915_ _05911_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_120_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29242_ clknet_leaf_243_clock _02255_ VGND VGND VPWR VPWR decode.regfile.registers_0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_26454_ _09434_ _09558_ VGND VGND VPWR VPWR _09571_ sky130_fd_sc_hd__nand2_1
X_23666_ _07981_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20878_ _05917_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__clkbuf_1
X_25405_ _08945_ _08946_ VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29173_ clknet_leaf_184_clock _02186_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_22617_ csr._minstret_T_3\[53\] csr._minstret_T_3\[52\] _07185_ net2212 VGND VGND
+ VPWR VPWR _07188_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_187_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26385_ net1859 _09492_ _09530_ _09525_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__o211a_1
X_23597_ _07944_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28124_ clknet_leaf_80_clock _01146_ VGND VGND VPWR VPWR csr.minstret\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_148_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25336_ _08891_ net2674 VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22548_ _06377_ _07138_ _07139_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_23_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28055_ clknet_leaf_196_clock _01077_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25267_ _08863_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22479_ fetch.bht.bhtTable_target_pc\[12\]\[0\] fetch.bht.bhtTable_target_pc\[13\]\[0\]
+ fetch.bht.bhtTable_target_pc\[14\]\[0\] fetch.bht.bhtTable_target_pc\[15\]\[0\]
+ _07069_ _07072_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_94_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15020_ _10969_ VGND VGND VPWR VPWR _11029_ sky130_fd_sc_hd__buf_2
X_27006_ clknet_leaf_341_clock _00035_ VGND VGND VPWR VPWR decode.regfile.registers_22\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_24218_ _08283_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25198_ _09880_ _09883_ _08801_ VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24149_ net1270 execute.io_target_pc\[29\] _06427_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28957_ clknet_leaf_178_clock _01970_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16971_ _11017_ _12539_ _12502_ decode.regfile.registers_8\[5\] VGND VGND VPWR VPWR
+ _12931_ sky130_fd_sc_hd__or4b_1
XFILLER_0_120_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18710_ _04008_ _03976_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27908_ clknet_leaf_70_clock _00937_ VGND VGND VPWR VPWR csr._mcycle_T_2\[29\] sky130_fd_sc_hd__dfxtp_2
X_15922_ decode.regfile.registers_23\[15\] _11088_ _11877_ _11903_ VGND VGND VPWR
+ VPWR _11904_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_53_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19690_ _04294_ _04371_ _04301_ _04770_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__or4_1
X_28888_ clknet_leaf_122_clock _01901_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18641_ _10090_ _10089_ memory.csr_read_data_out_reg\[21\] _10010_ VGND VGND VPWR
+ VPWR _03940_ sky130_fd_sc_hd__o2bb2a_1
X_15853_ _10956_ decode.regfile.registers_22\[14\] _11093_ _11264_ _11265_ VGND VGND
+ VPWR VPWR _11836_ sky130_fd_sc_hd__o2111a_1
X_27839_ clknet_leaf_326_clock _00868_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_14804_ _10805_ _10806_ VGND VGND VPWR VPWR _10847_ sky130_fd_sc_hd__nand2_1
X_18572_ _03768_ _03769_ _03770_ _03870_ _03670_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__o41a_2
XFILLER_0_203_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15784_ decode.regfile.registers_3\[12\] _11111_ _11167_ _11146_ _11768_ VGND VGND
+ VPWR VPWR _11769_ sky130_fd_sc_hd__a311o_1
X_17523_ _11020_ _12491_ _12666_ decode.regfile.registers_14\[18\] _12670_ VGND VGND
+ VPWR VPWR _13470_ sky130_fd_sc_hd__o32a_1
X_29509_ clknet_5_22__leaf_clock _02522_ VGND VGND VPWR VPWR decode.regfile.registers_8\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_14735_ _10684_ _10777_ VGND VGND VPWR VPWR _10778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_203_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14666_ execute.io_target_pc\[13\] VGND VGND VPWR VPWR _10709_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17454_ decode.regfile.registers_22\[16\] _13100_ _13402_ _13289_ VGND VGND VPWR
+ VPWR _13403_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16405_ _11088_ _12372_ _12373_ VGND VGND VPWR VPWR _12374_ sky130_fd_sc_hd__a21o_1
X_13617_ _09961_ VGND VGND VPWR VPWR _09978_ sky130_fd_sc_hd__buf_4
XFILLER_0_229_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14597_ _10639_ VGND VGND VPWR VPWR _10640_ sky130_fd_sc_hd__buf_4
X_17385_ decode.regfile.registers_27\[14\] _12507_ _12520_ _12495_ _13335_ VGND VGND
+ VPWR VPWR _13336_ sky130_fd_sc_hd__o311a_1
XFILLER_0_223_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19124_ _04412_ _03704_ _04332_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13548_ _09914_ _09887_ _09917_ net392 VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__a31o_1
X_16336_ _11756_ decode.regfile.registers_28\[26\] _11871_ _11681_ _11448_ VGND VGND
+ VPWR VPWR _12307_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_229_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19055_ _04350_ _04351_ _04352_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16267_ decode.regfile.registers_14\[25\] _11206_ _11272_ decode.regfile.registers_15\[25\]
+ _11201_ VGND VGND VPWR VPWR _12239_ sky130_fd_sc_hd__a221o_1
XFILLER_0_152_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18006_ _10938_ decode.regfile.registers_25\[30\] _12505_ _12811_ VGND VGND VPWR
+ VPWR _03403_ sky130_fd_sc_hd__or4_1
X_15218_ _11125_ VGND VGND VPWR VPWR _11215_ sky130_fd_sc_hd__buf_4
XFILLER_0_72_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16198_ decode.regfile.registers_14\[23\] _11360_ _11274_ decode.regfile.registers_15\[23\]
+ _11202_ VGND VGND VPWR VPWR _12172_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15149_ _11145_ VGND VGND VPWR VPWR _11146_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_1193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19957_ net1266 _03599_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18908_ _04204_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_203_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19888_ _04799_ _04798_ _04805_ _04729_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_203_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18839_ _03715_ _03725_ _04135_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__or3b_1
XFILLER_0_223_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_195_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21850_ csr.io_mret_vector\[4\] _09881_ _06040_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20801_ _03582_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21781_ net2093 csr.io_mem_pc\[29\] _06450_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23520_ decode.id_ex_memread_reg VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_1175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20732_ _05056_ _05836_ csr.mcycle\[23\] _05537_ _05748_ VGND VGND VPWR VPWR _05837_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_158_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_186_Right_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23451_ _03546_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20663_ decode.id_ex_funct3_reg\[1\] _03594_ _05569_ VGND VGND VPWR VPWR _05791_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_163_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22402_ _06790_ _06992_ _06994_ _06996_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_154_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26170_ _09398_ _09390_ VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23382_ fetch.bht.bhtTable_target_pc\[8\]\[29\] fetch.bht.bhtTable_target_pc\[9\]\[29\]
+ fetch.bht.bhtTable_target_pc\[10\]\[29\] fetch.bht.bhtTable_target_pc\[11\]\[29\]
+ _07669_ _07656_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20594_ _05627_ csr.io_mret_vector\[21\] _05603_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25121_ _06138_ net2038 _08562_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22333_ net72 _06927_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25052_ csr.mcycle\[20\] _03554_ csr.mcycle\[21\] _08742_ VGND VGND VPWR VPWR _08748_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_103_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22264_ _06858_ _06650_ _06686_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24003_ net1247 execute.io_target_pc\[22\] _08164_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__mux2_1
X_21215_ _06102_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__clkbuf_1
X_29860_ clknet_leaf_303_clock _02873_ VGND VGND VPWR VPWR decode.regfile.registers_19\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_22195_ _00002_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__clkbuf_8
X_28811_ clknet_leaf_94_clock _01824_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_21146_ _06066_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29791_ clknet_leaf_309_clock _02804_ VGND VGND VPWR VPWR decode.regfile.registers_17\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28742_ clknet_leaf_94_clock _01755_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21077_ _05864_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__buf_4
X_25954_ _09241_ VGND VGND VPWR VPWR _09270_ sky130_fd_sc_hd__buf_2
XFILLER_0_214_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20028_ _04018_ _10711_ _05241_ _05243_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__o211ai_2
X_24905_ csr._mcycle_T_3\[35\] _08649_ net645 VGND VGND VPWR VPWR _08651_ sky130_fd_sc_hd__a21oi_1
X_28673_ clknet_leaf_174_clock _01686_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_25885_ _08958_ _09223_ VGND VGND VPWR VPWR _09230_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_122_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27624_ clknet_leaf_48_clock _00653_ VGND VGND VPWR VPWR execute.io_reg_pc\[1\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_87_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24836_ _08605_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24767_ _08569_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27555_ clknet_leaf_52_clock _00584_ VGND VGND VPWR VPWR execute.io_mem_memwrite
+ sky130_fd_sc_hd__dfxtp_1
X_21979_ csr.mscratch\[13\] _06588_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__or2_1
Xrebuffer80 net199 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__buf_1
X_14520_ _09900_ fetch.btb.io_branch VGND VGND VPWR VPWR _10565_ sky130_fd_sc_hd__nand2_2
Xrebuffer91 net317 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__buf_1
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23718_ net787 _10787_ _08003_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__mux2_1
X_26506_ _09410_ _09589_ VGND VGND VPWR VPWR _09601_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27486_ clknet_leaf_38_clock _00515_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_2
X_24698_ _08060_ net1199 _08531_ VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29225_ clknet_leaf_105_clock _02238_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14451_ _10025_ _10517_ VGND VGND VPWR VPWR _10519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23649_ net1473 _10868_ _07972_ VGND VGND VPWR VPWR _07973_ sky130_fd_sc_hd__mux2_1
X_26437_ _09533_ VGND VGND VPWR VPWR _09561_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17170_ decode.regfile.registers_21\[9\] _12682_ _12806_ VGND VGND VPWR VPWR _13126_
+ sky130_fd_sc_hd__o21a_1
X_29156_ clknet_leaf_205_clock _02169_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26368_ net2718 _09518_ _09521_ _09512_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14382_ net464 _10477_ _10479_ _10468_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16121_ _10994_ VGND VGND VPWR VPWR _12097_ sky130_fd_sc_hd__buf_2
X_28107_ clknet_leaf_82_clock _01129_ VGND VGND VPWR VPWR csr.minstret\[12\] sky130_fd_sc_hd__dfxtp_1
X_25319_ _08880_ net2663 VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29087_ clknet_leaf_72_clock _02100_ VGND VGND VPWR VPWR csr._mcycle_T_3\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26299_ net2700 _09475_ _09481_ _09471_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16052_ decode.regfile.registers_8\[19\] _11044_ _11174_ VGND VGND VPWR VPWR _12030_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_228_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28038_ clknet_leaf_168_clock _01060_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15003_ _11013_ VGND VGND VPWR VPWR _11014_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_161_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19811_ _05082_ _05083_ _04589_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_23_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19742_ _04982_ _04993_ _04992_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__a21bo_1
X_16954_ _10595_ VGND VGND VPWR VPWR _12915_ sky130_fd_sc_hd__buf_2
XFILLER_0_194_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15905_ _11880_ _11886_ VGND VGND VPWR VPWR _11887_ sky130_fd_sc_hd__nand2_1
X_19673_ _04805_ _04538_ _04728_ _04883_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__a31o_1
XFILLER_0_217_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16885_ decode.regfile.registers_9\[3\] _12606_ _12845_ _12846_ VGND VGND VPWR VPWR
+ _12847_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_218_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18624_ _03919_ _03920_ _03921_ _03922_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_154_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15836_ _11225_ _11125_ _11216_ _11819_ VGND VGND VPWR VPWR _11820_ sky130_fd_sc_hd__o31a_1
XFILLER_0_220_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18555_ _03703_ _03766_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__xor2_4
XFILLER_0_204_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15767_ _11436_ decode.regfile.registers_26\[11\] _11676_ _10980_ _11564_ VGND VGND
+ VPWR VPWR _11753_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17506_ _12712_ decode.regfile.registers_24\[18\] VGND VGND VPWR VPWR _13453_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_190_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14718_ csr.io_mem_pc\[5\] csr.io_mem_pc\[6\] _09928_ VGND VGND VPWR VPWR _10761_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18486_ _03715_ _03725_ net204 VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_190_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15698_ _11571_ decode.regfile.registers_30\[10\] _11039_ _11032_ _11033_ VGND VGND
+ VPWR VPWR _11685_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_16_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17437_ decode.regfile.registers_4\[16\] _12548_ _13145_ decode.regfile.registers_5\[16\]
+ _12614_ VGND VGND VPWR VPWR _13386_ sky130_fd_sc_hd__a221oi_1
X_14649_ decode.id_ex_pc_reg\[19\] VGND VGND VPWR VPWR _10692_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_16 _03944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 _08939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_38 _10019_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17368_ _12611_ _13317_ _13318_ VGND VGND VPWR VPWR _13319_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19107_ _04390_ _04397_ _04404_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__or3_2
XFILLER_0_166_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16319_ _11690_ _12289_ VGND VGND VPWR VPWR _12290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17299_ _12516_ _13248_ _13249_ _13251_ VGND VGND VPWR VPWR _13252_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_209_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_209_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19038_ _04332_ _04333_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_209_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput101 net101 VGND VGND VPWR VPWR io_memory_address[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput112 net112 VGND VGND VPWR VPWR io_memory_address[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput123 net123 VGND VGND VPWR VPWR io_memory_address[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput134 net134 VGND VGND VPWR VPWR io_memory_size[1] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput145 net145 VGND VGND VPWR VPWR io_memory_write_data[18] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_205_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput156 net156 VGND VGND VPWR VPWR io_memory_write_data[28] sky130_fd_sc_hd__clkbuf_4
X_21000_ _05983_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__clkbuf_1
Xoutput167 net167 VGND VGND VPWR VPWR io_memory_write_data[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_7 _00932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_215_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22951_ csr._csr_read_data_T_8\[4\] _06039_ csr.io_mret_vector\[4\] _06463_ VGND
+ VGND VPWR VPWR _07400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21902_ _06540_ _06519_ _06520_ _06541_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_3_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25670_ net2595 _09095_ _09105_ _09100_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__o211a_1
X_22882_ net1804 _10759_ _07335_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24621_ net1063 execute.io_target_pc\[0\] _07308_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21833_ _06457_ _06459_ _06472_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27340_ clknet_leaf_43_clock _00369_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[13\]
+ sky130_fd_sc_hd__dfxtp_4
X_24552_ _08457_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_156_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21764_ net1218 csr.io_mem_pc\[21\] _06439_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23503_ net1377 _07890_ _07887_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__or3b_1
X_27271_ clknet_leaf_13_clock _00300_ VGND VGND VPWR VPWR decode.regfile.registers_30\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20715_ _00514_ _05703_ _05826_ net182 net2691 VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__a32o_1
X_24483_ _08421_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__clkbuf_1
X_21695_ csr.minstret\[25\] csr.minstret\[26\] csr.io_inst_retired _06380_ VGND VGND
+ VPWR VPWR _06398_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29010_ clknet_leaf_104_clock _02023_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26222_ _09434_ _09413_ VGND VGND VPWR VPWR _09435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23434_ _10579_ _07847_ _05206_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20646_ csr.mscratch\[29\] _05591_ _05611_ _05672_ _05776_ VGND VGND VPWR VPWR _05777_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_117_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26153_ net1982 _09373_ _09386_ _09370_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__o211a_1
X_23365_ _06795_ _07783_ _07789_ _07064_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20577_ csr.mscratch\[19\] _05592_ _05611_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_115_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25104_ _08780_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22316_ _06730_ _06910_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__and2b_1
X_26084_ _08931_ _09340_ VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23296_ _07722_ _07723_ _07724_ _07725_ _07371_ _07127_ VGND VGND VPWR VPWR _07726_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_186_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25035_ csr._mcycle_T_2\[16\] _08704_ net2541 VGND VGND VPWR VPWR _08737_ sky130_fd_sc_hd__a21oi_1
X_29912_ clknet_leaf_304_clock _02925_ VGND VGND VPWR VPWR decode.regfile.registers_20\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22247_ _06685_ _06839_ _06687_ _06841_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_104_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29843_ clknet_leaf_296_clock _02856_ VGND VGND VPWR VPWR decode.regfile.registers_18\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_22178_ _06661_ _06770_ _06629_ _06772_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__a211oi_1
X_21129_ _06050_ _06046_ net2348 VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_50_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29774_ clknet_leaf_293_clock _02787_ VGND VGND VPWR VPWR decode.regfile.registers_16\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26986_ net504 _09866_ _09876_ _06396_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_89_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28725_ clknet_leaf_116_clock _01738_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13951_ net2538 _10226_ _10229_ _10219_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__o211a_1
X_25937_ _08935_ _09253_ VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_222_Right_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28656_ clknet_leaf_120_clock _01669_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_16670_ _11016_ _10597_ decode.immGen._imm_T_24\[17\] VGND VGND VPWR VPWR _12635_
+ sky130_fd_sc_hd__nor3_1
X_13882_ net1695 _10180_ _10187_ _10188_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__o211a_1
X_25868_ _08941_ _09210_ VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27607_ clknet_leaf_158_clock _00636_ VGND VGND VPWR VPWR execute.io_target_pc\[16\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_9_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15621_ _11571_ decode.regfile.registers_30\[8\] _11039_ _11032_ _11033_ VGND VGND
+ VPWR VPWR _11610_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_201_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24819_ _08111_ net2233 _08596_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__mux2_1
X_28587_ clknet_leaf_94_clock _01600_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25799_ net2540 _09170_ _09180_ _09169_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_206 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_217 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _03638_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__buf_4
XFILLER_0_90_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27538_ clknet_leaf_155_clock _00567_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_29_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_228 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15552_ decode.regfile.registers_4\[6\] _10636_ _11138_ VGND VGND VPWR VPWR _11543_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_239 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14503_ fetch.btb.btbTable\[0\]\[1\] fetch.btb.btbTable\[1\]\[1\] fetch.btb.btbTable\[2\]\[1\]
+ fetch.btb.btbTable\[3\]\[1\] _09891_ _09888_ VGND VGND VPWR VPWR _10548_ sky130_fd_sc_hd__mux4_1
XFILLER_0_194_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ decode.regfile.registers_17\[4\] _10652_ _11112_ _11118_ _11475_ VGND VGND
+ VPWR VPWR _11476_ sky130_fd_sc_hd__a41o_1
XFILLER_0_56_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18271_ decode.id_ex_rs2_data_reg\[2\] _03596_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27469_ clknet_leaf_54_clock _00498_ VGND VGND VPWR VPWR csr.io_csr_address\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_13_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29208_ clknet_leaf_157_clock _02221_ VGND VGND VPWR VPWR fetch.btb.btbTable\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_17222_ _13091_ _13176_ decode.regfile.registers_27\[10\] _13050_ VGND VGND VPWR
+ VPWR _13177_ sky130_fd_sc_hd__or4_1
XFILLER_0_154_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14434_ _09964_ _10507_ VGND VGND VPWR VPWR _10510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput14 io_fetch_data[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
X_29139_ clknet_leaf_79_clock _02152_ VGND VGND VPWR VPWR csr.mcycle\[23\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput25 net374 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14365_ _09984_ _10464_ VGND VGND VPWR VPWR _10470_ sky130_fd_sc_hd__nand2_1
X_17153_ decode.regfile.registers_7\[9\] _10617_ _13020_ _12888_ VGND VGND VPWR VPWR
+ _13109_ sky130_fd_sc_hd__a31o_1
Xinput36 io_memory_read_data[11] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput47 io_memory_read_data[21] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
XFILLER_0_141_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput58 io_memory_read_data[31] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_1
X_16104_ _10989_ _10977_ _10956_ _11114_ _12080_ VGND VGND VPWR VPWR _12081_ sky130_fd_sc_hd__a41o_1
XFILLER_0_126_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17084_ _11015_ _10937_ decode.regfile.registers_23\[7\] _13041_ VGND VGND VPWR VPWR
+ _13042_ sky130_fd_sc_hd__or4_1
Xhold809 fetch.bht.bhtTable_tag\[4\]\[14\] VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ _10008_ _10420_ VGND VGND VPWR VPWR _10430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16035_ _11445_ _12012_ _12013_ VGND VGND VPWR VPWR _12014_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17986_ decode.regfile.registers_1\[30\] _12932_ _12830_ _03382_ VGND VGND VPWR VPWR
+ _03383_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_200_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1509 fetch.bht.bhtTable_tag\[14\]\[0\] VGND VGND VPWR VPWR net1736 sky130_fd_sc_hd__dlygate4sd3_1
X_19725_ _04995_ _04999_ _05000_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16937_ _12659_ _12896_ _12897_ VGND VGND VPWR VPWR _12898_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19656_ _04204_ _04206_ _04201_ _03938_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_192_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16868_ _12829_ VGND VGND VPWR VPWR _12830_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_0_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18607_ _03797_ _03905_ _03785_ _10068_ _03889_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__a221oi_4
X_15819_ decode.regfile.registers_3\[13\] _11157_ _11140_ _11145_ VGND VGND VPWR VPWR
+ _11803_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19587_ _04860_ _04832_ _04864_ _04868_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__o31a_1
XFILLER_0_172_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16799_ _12492_ decode.regfile.registers_29\[1\] _12711_ _12762_ _12702_ VGND VGND
+ VPWR VPWR _12763_ sky130_fd_sc_hd__o221a_1
XFILLER_0_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18538_ _03759_ _03832_ _03727_ _03836_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__o211a_2
XFILLER_0_88_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18469_ decode.id_ex_ex_rs1_reg\[0\] _03642_ _03647_ _03646_ _03648_ VGND VGND VPWR
+ VPWR _03768_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_185_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20500_ csr.mscratch\[9\] _05592_ _05611_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21480_ _06109_ net2055 _06252_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20431_ _05586_ _05588_ csr.mcycle\[2\] VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23150_ net72 _07536_ _07537_ _07588_ _07535_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__o311a_1
X_20362_ csr.io_csr_address\[2\] net358 VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22101_ fetch.bht.bhtTable_tag\[8\]\[7\] fetch.bht.bhtTable_tag\[9\]\[7\] fetch.bht.bhtTable_tag\[10\]\[7\]
+ fetch.bht.bhtTable_tag\[11\]\[7\] _06674_ _06675_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_228_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_998 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_228_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23081_ fetch.bht.bhtTable_target_pc\[8\]\[11\] fetch.bht.bhtTable_target_pc\[9\]\[11\]
+ fetch.bht.bhtTable_target_pc\[10\]\[11\] fetch.bht.bhtTable_target_pc\[11\]\[11\]
+ _07123_ _07111_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20293_ _10806_ _05468_ _05416_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_110_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22032_ _06626_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_181_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26840_ net2222 _09753_ _09792_ _09784_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23983_ _08162_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__clkbuf_1
X_26771_ net2497 _09752_ _09754_ _09743_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28510_ clknet_leaf_196_clock _01523_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22934_ _07066_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__clkbuf_8
X_25722_ _09110_ VGND VGND VPWR VPWR _09136_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_108_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29490_ clknet_leaf_264_clock _02503_ VGND VGND VPWR VPWR decode.regfile.registers_7\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28441_ clknet_leaf_54_clock _01454_ VGND VGND VPWR VPWR decode.control.io_funct7\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22865_ net848 _10800_ _07324_ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25653_ net2672 _09095_ _09096_ _09087_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24604_ _08484_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21816_ _06461_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__clkbuf_4
X_28372_ clknet_leaf_213_clock _01385_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_25584_ net2641 _09052_ _09056_ _09046_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22796_ net1034 csr.io_mem_pc\[12\] _07286_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24535_ _08095_ net1926 _08439_ VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27323_ clknet_leaf_26_clock _00352_ VGND VGND VPWR VPWR decode.id_ex_ex_rs1_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21747_ net1076 _10871_ _06428_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24466_ _08093_ net1808 _08411_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27254_ clknet_leaf_32_clock _00283_ VGND VGND VPWR VPWR decode.regfile.registers_30\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_21678_ _06385_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23417_ _07838_ _07070_ _07080_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__a21o_1
XFILLER_0_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26205_ net2400 _09419_ _09423_ _09418_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20629_ _05627_ csr.io_mret_vector\[26\] _05603_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27185_ clknet_leaf_352_clock _00214_ VGND VGND VPWR VPWR decode.regfile.registers_28\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24397_ net1776 execute.io_target_pc\[21\] _08367_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14150_ net484 _10332_ _10345_ _10344_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_330_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_330_clock
+ sky130_fd_sc_hd__clkbuf_8
X_26136_ net2441 _09373_ _09375_ _09370_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__o211a_1
X_23348_ _07619_ _07573_ _07620_ _07774_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14081_ _10042_ _10299_ VGND VGND VPWR VPWR _10306_ sky130_fd_sc_hd__nand2_1
X_26067_ net2621 _09329_ _09335_ _09333_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__o211a_1
X_23279_ _07100_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25018_ _06331_ _08724_ _08725_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__nor3_1
XFILLER_0_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_345_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_345_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_37_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17840_ _12654_ _03239_ _03240_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__a21oi_2
X_29826_ clknet_leaf_307_clock _02839_ VGND VGND VPWR VPWR decode.regfile.registers_18\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17771_ decode.regfile.registers_22\[24\] _13100_ _03173_ _13289_ VGND VGND VPWR
+ VPWR _03174_ sky130_fd_sc_hd__a211o_1
X_29757_ clknet_leaf_309_clock _02770_ VGND VGND VPWR VPWR decode.regfile.registers_16\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14983_ _10950_ _10952_ _11000_ decode.control.io_funct7\[6\] VGND VGND VPWR VPWR
+ _11001_ sky130_fd_sc_hd__o31a_1
X_26969_ _10091_ _09862_ VGND VGND VPWR VPWR _09868_ sky130_fd_sc_hd__nand2_1
X_19510_ _04083_ _04084_ _04081_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__a21oi_1
X_28708_ clknet_leaf_131_clock _01721_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16722_ _12686_ VGND VGND VPWR VPWR _12687_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13934_ _10058_ _10210_ VGND VGND VPWR VPWR _10220_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29688_ clknet_leaf_289_clock _02701_ VGND VGND VPWR VPWR decode.regfile.registers_13\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19441_ _04728_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__buf_6
XFILLER_0_92_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28639_ clknet_leaf_176_clock _01652_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16653_ _12617_ VGND VGND VPWR VPWR _12618_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13865_ _10081_ _10177_ VGND VGND VPWR VPWR _10179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15604_ decode.regfile.registers_16\[7\] _11359_ _11574_ _11593_ _11127_ VGND VGND
+ VPWR VPWR _11594_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19372_ _04142_ _04143_ _04639_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__o21ai_1
X_16584_ _12548_ VGND VGND VPWR VPWR _12549_ sky130_fd_sc_hd__buf_4
X_13796_ net676 _10083_ _10129_ _10132_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18323_ _03594_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__buf_4
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15535_ _11346_ _11253_ _11064_ decode.regfile.registers_29\[5\] _11526_ VGND VGND
+ VPWR VPWR _11527_ sky130_fd_sc_hd__o221a_1
XFILLER_0_96_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18254_ _03586_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15466_ _11300_ decode.regfile.registers_0\[4\] _11155_ _11458_ VGND VGND VPWR VPWR
+ _11459_ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17205_ _11021_ _12567_ _12586_ _13159_ VGND VGND VPWR VPWR _13160_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14417_ _10122_ _10487_ VGND VGND VPWR VPWR _10499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_835 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18185_ decode.control.io_funct7\[6\] decode.control.io_funct7\[4\] decode.control.io_funct7\[3\]
+ decode.control.io_funct7\[1\] VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15397_ decode.regfile.registers_21\[2\] _11060_ _11098_ _11227_ _11391_ VGND VGND
+ VPWR VPWR _11392_ sky130_fd_sc_hd__o311a_1
X_17136_ _12697_ VGND VGND VPWR VPWR _13093_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14348_ _10142_ _10418_ VGND VGND VPWR VPWR _10459_ sky130_fd_sc_hd__nand2_1
Xhold606 fetch.bht.bhtTable_target_pc\[8\]\[29\] VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold617 _01140_ VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold628 decode.regfile.registers_26\[6\] VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 fetch.bht.bhtTable_target_pc\[2\]\[5\] VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14279_ _10418_ VGND VGND VPWR VPWR _10420_ sky130_fd_sc_hd__clkbuf_4
X_17067_ decode.regfile.registers_10\[7\] _12790_ _12792_ VGND VGND VPWR VPWR _13025_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16018_ _10648_ _10624_ _11084_ _11989_ _11996_ VGND VGND VPWR VPWR _11997_ sky130_fd_sc_hd__o32a_1
XFILLER_0_0_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_223_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 decode.regfile.registers_17\[29\] VGND VGND VPWR VPWR net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2018 fetch.bht.bhtTable_tag\[5\]\[16\] VGND VGND VPWR VPWR net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2029 csr._csr_read_data_T_8\[18\] VGND VGND VPWR VPWR net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1306 decode.regfile.registers_16\[2\] VGND VGND VPWR VPWR net1533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 decode.regfile.registers_18\[19\] VGND VGND VPWR VPWR net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1328 decode.regfile.registers_5\[17\] VGND VGND VPWR VPWR net1555 sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ _10938_ decode.regfile.registers_25\[29\] _12505_ _12811_ VGND VGND VPWR
+ VPWR _03367_ sky130_fd_sc_hd__or4_1
XFILLER_0_224_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1339 fetch.bht.bhtTable_tag\[13\]\[14\] VGND VGND VPWR VPWR net1566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19708_ _04984_ _04897_ _04268_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20980_ _05972_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19639_ _04918_ _04875_ _04247_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_1254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22650_ csr._mcycle_T_2\[2\] _07210_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21601_ csr.minstret\[0\] csr.minstret\[1\] _06323_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_217_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22581_ csr._minstret_T_3\[41\] _07160_ _07163_ _07164_ VGND VGND VPWR VPWR _01263_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_174_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24320_ _08336_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21532_ _06103_ net2083 _06284_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24251_ _08078_ net1653 _08300_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21463_ _06247_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23202_ _07635_ _07636_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20414_ _05572_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__clkbuf_4
X_24182_ _08076_ net1626 _08255_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21394_ _06186_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__buf_4
XFILLER_0_114_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23133_ net225 _07536_ _07537_ _07572_ _07535_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__o311a_1
XFILLER_0_113_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20345_ _05403_ _05418_ _03517_ _03551_ _05510_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_4_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28990_ clknet_leaf_173_clock _02003_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23064_ fetch.bht.bhtTable_target_pc\[0\]\[10\] fetch.bht.bhtTable_target_pc\[1\]\[10\]
+ fetch.bht.bhtTable_target_pc\[2\]\[10\] fetch.bht.bhtTable_target_pc\[3\]\[10\]
+ _07407_ _07115_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__mux4_1
X_27941_ clknet_leaf_235_clock _00963_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20276_ _10694_ _10710_ _05452_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22015_ csr._mcycle_T_2\[29\] _06600_ _06612_ _06605_ VGND VGND VPWR VPWR _01249_
+ sky130_fd_sc_hd__o211a_1
X_27872_ clknet_leaf_327_clock _00901_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2530 csr._csr_read_data_T_8\[29\] VGND VGND VPWR VPWR net2757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29611_ clknet_leaf_276_clock _02624_ VGND VGND VPWR VPWR decode.regfile.registers_11\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2541 net69 VGND VGND VPWR VPWR net2768 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26823_ _09701_ VGND VGND VPWR VPWR _09784_ sky130_fd_sc_hd__buf_4
XFILLER_0_192_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2552 net85 VGND VGND VPWR VPWR net2779 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2563 csr._mcycle_T_2\[5\] VGND VGND VPWR VPWR net2790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2574 csr._minstret_T_3\[58\] VGND VGND VPWR VPWR net2801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1840 decode.regfile.registers_2\[29\] VGND VGND VPWR VPWR net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29542_ clknet_leaf_267_clock _02555_ VGND VGND VPWR VPWR decode.regfile.registers_9\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26754_ _09432_ _09733_ VGND VGND VPWR VPWR _09744_ sky130_fd_sc_hd__nand2_1
Xhold1851 decode.regfile.registers_28\[16\] VGND VGND VPWR VPWR net2078 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23966_ net986 execute.io_target_pc\[4\] _08153_ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__mux2_1
Xhold1862 fetch.bht.bhtTable_tag\[5\]\[2\] VGND VGND VPWR VPWR net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1873 fetch.bht.bhtTable_target_pc\[6\]\[8\] VGND VGND VPWR VPWR net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1884 fetch.bht.bhtTable_target_pc\[9\]\[16\] VGND VGND VPWR VPWR net2111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1895 decode.io_id_pc\[27\] VGND VGND VPWR VPWR net2122 sky130_fd_sc_hd__dlygate4sd3_1
X_25705_ net599 _09125_ _09126_ _09115_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__o211a_1
X_22917_ _07367_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__buf_4
X_29473_ clknet_leaf_252_clock _02486_ VGND VGND VPWR VPWR decode.regfile.registers_7\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_23897_ net1083 _08055_ _06179_ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__mux2_1
X_26685_ _09438_ _09664_ VGND VGND VPWR VPWR _09704_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28424_ clknet_leaf_47_clock _01437_ VGND VGND VPWR VPWR decode.control.io_funct3\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_22848_ net964 _10812_ _09898_ VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__mux2_1
X_25636_ _08990_ VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__buf_2
X_13650_ _10007_ VGND VGND VPWR VPWR _10008_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28355_ clknet_leaf_168_clock _01368_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13581_ _09939_ _09940_ VGND VGND VPWR VPWR _09946_ sky130_fd_sc_hd__nand2b_2
X_22779_ _06153_ net1611 _07276_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25567_ _08941_ _09036_ VGND VGND VPWR VPWR _09047_ sky130_fd_sc_hd__nand2_1
X_15320_ _10649_ _10631_ _11052_ decode.regfile.registers_11\[1\] _11315_ VGND VGND
+ VPWR VPWR _11316_ sky130_fd_sc_hd__o32a_1
X_27306_ clknet_leaf_13_clock _00335_ VGND VGND VPWR VPWR decode.regfile.registers_31\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24518_ _08440_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28286_ clknet_leaf_86_clock _01308_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25498_ _08948_ _09005_ VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27237_ clknet_leaf_364_clock _00266_ VGND VGND VPWR VPWR decode.regfile.registers_29\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_15251_ _10994_ _10981_ _10960_ _11215_ _10973_ VGND VGND VPWR VPWR _11248_ sky130_fd_sc_hd__o41a_2
X_24449_ _08076_ net1497 _08400_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14202_ _10374_ VGND VGND VPWR VPWR _10375_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15182_ _10629_ _11178_ net324 _11058_ VGND VGND VPWR VPWR _11179_ sky130_fd_sc_hd__and4_2
XFILLER_0_227_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27168_ clknet_leaf_359_clock _00197_ VGND VGND VPWR VPWR decode.regfile.registers_27\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_14133_ _09970_ _10333_ VGND VGND VPWR VPWR _10336_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26119_ net1952 _09356_ _09364_ _09359_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__o211a_1
X_19990_ net2722 _05219_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27099_ clknet_leaf_348_clock _00128_ VGND VGND VPWR VPWR decode.regfile.registers_25\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_284_clock clknet_5_20__leaf_clock VGND VGND VPWR VPWR clknet_leaf_284_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14064_ _09993_ _10288_ VGND VGND VPWR VPWR _10296_ sky130_fd_sc_hd__nand2_1
X_18941_ _03636_ _03767_ _04224_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__or4b_4
XFILLER_0_123_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18872_ _04062_ _04065_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29809_ clknet_leaf_295_clock _02822_ VGND VGND VPWR VPWR decode.regfile.registers_17\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_17823_ net509 _12872_ _03185_ _03224_ _03073_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_299_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_299_clock
+ sky130_fd_sc_hd__clkbuf_8
X_17754_ decode.regfile.registers_5\[24\] _12509_ _12614_ _12735_ VGND VGND VPWR VPWR
+ _03157_ sky130_fd_sc_hd__o31a_1
X_14966_ _10990_ VGND VGND VPWR VPWR _10991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16705_ _12669_ VGND VGND VPWR VPWR _12670_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13917_ _10198_ VGND VGND VPWR VPWR _10210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17685_ _12792_ _03088_ _03089_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__a21o_1
X_14897_ _10604_ VGND VGND VPWR VPWR _10933_ sky130_fd_sc_hd__buf_4
XFILLER_0_187_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19424_ _04474_ _04243_ net312 _04711_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_222_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_222_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16636_ _11016_ _10605_ decode.immGen._imm_T_24\[17\] _12509_ VGND VGND VPWR VPWR
+ _12601_ sky130_fd_sc_hd__or4_2
XFILLER_0_159_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13848_ net685 _10167_ _10169_ _10162_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19355_ _04017_ _04015_ _04016_ _04282_ _04289_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__a311o_1
XFILLER_0_128_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16567_ _12531_ VGND VGND VPWR VPWR _12532_ sky130_fd_sc_hd__buf_4
XFILLER_0_18_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13779_ _10117_ _10075_ VGND VGND VPWR VPWR _10118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18306_ _03618_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__clkbuf_1
X_15518_ decode.regfile.registers_11\[5\] _11180_ _11509_ decode.regfile.registers_10\[5\]
+ _11186_ VGND VGND VPWR VPWR _11510_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_73_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19286_ _04579_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_84_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16498_ decode.regfile.registers_7\[31\] _11308_ _11169_ decode.regfile.registers_6\[31\]
+ _11133_ VGND VGND VPWR VPWR _12464_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_127_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_237_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_237_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_212_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18237_ csr._mcycle_T_3\[49\] csr._mcycle_T_3\[48\] csr._mcycle_T_3\[47\] csr._mcycle_T_3\[46\]
+ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_212_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15449_ _11346_ _11253_ _11064_ decode.regfile.registers_29\[3\] _11442_ VGND VGND
+ VPWR VPWR _11443_ sky130_fd_sc_hd__o221a_1
XFILLER_0_66_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_212_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18168_ _03463_ _03464_ _10921_ decode.control.io_funct7\[3\] VGND VGND VPWR VPWR
+ _03512_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_170_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold403 decode.regfile.registers_27\[12\] VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17119_ decode.regfile.registers_18\[8\] _12572_ _12562_ _13075_ VGND VGND VPWR VPWR
+ _13076_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold414 decode.regfile.registers_10\[11\] VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold425 decode.regfile.registers_28\[17\] VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ _03469_ _03467_ _03474_ net2459 VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_106_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold436 decode.regfile.registers_19\[16\] VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold447 decode.regfile.registers_2\[11\] VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__dlygate4sd3_1
X_20130_ _00566_ _05226_ _05338_ _05239_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__o22a_1
Xhold458 decode.regfile.registers_23\[11\] VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 decode.regfile.registers_27\[24\] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap188 _03821_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_4
XFILLER_0_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap199 _03745_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_221_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20061_ _05270_ _05272_ _05276_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_141_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1103 fetch.bht.bhtTable_target_pc\[5\]\[19\] VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1114 decode.regfile.registers_19\[19\] VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1125 fetch.bht.bhtTable_target_pc\[4\]\[21\] VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1136 fetch.bht.bhtTable_target_pc\[7\]\[21\] VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__dlygate4sd3_1
X_23820_ _08067_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1147 decode.regfile.registers_24\[2\] VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 fetch.bht.bhtTable_tag\[8\]\[12\] VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 fetch.bht.bhtTable_tag\[11\]\[0\] VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23751_ _06113_ net1357 _09907_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__mux2_1
X_20963_ _05963_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_219_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22702_ net526 _07236_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23682_ _09885_ _09894_ _09917_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__and3_4
XFILLER_0_36_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26470_ _09450_ _09579_ VGND VGND VPWR VPWR _09581_ sky130_fd_sc_hd__nand2_1
XFILLER_0_215_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20894_ _05926_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_172_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22633_ net2780 net1524 _07196_ _07198_ _06336_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__a311oi_1
XTAP_TAPCELL_ROW_172_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25421_ net200 VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__buf_4
XFILLER_0_222_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28140_ clknet_leaf_195_clock _01162_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25352_ _09969_ VGND VGND VPWR VPWR _08910_ sky130_fd_sc_hd__clkbuf_4
X_22564_ csr._minstret_T_3\[38\] _07147_ net2291 VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24303_ _08327_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__clkbuf_1
X_21515_ _06275_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28071_ clknet_leaf_222_clock _01093_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25283_ _08869_ net2558 VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22495_ _10757_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24234_ _08062_ net1371 _08289_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27022_ clknet_leaf_333_clock _00051_ VGND VGND VPWR VPWR decode.regfile.registers_22\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21446_ _06238_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_20_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24165_ _08256_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21377_ _06201_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23116_ fetch.bht.bhtTable_target_pc\[8\]\[13\] fetch.bht.bhtTable_target_pc\[9\]\[13\]
+ fetch.bht.bhtTable_target_pc\[10\]\[13\] fetch.bht.bhtTable_target_pc\[11\]\[13\]
+ _07555_ _07114_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__mux4_1
X_20328_ _05496_ _05497_ _05411_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__a21oi_1
X_28973_ clknet_leaf_103_clock _01986_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_24096_ _08220_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__clkbuf_1
Xhold970 decode.regfile.registers_15\[10\] VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold981 decode.regfile.registers_27\[27\] VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold992 fetch.bht.bhtTable_target_pc\[8\]\[16\] VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__dlygate4sd3_1
X_23047_ _07489_ _07490_ _07406_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27924_ clknet_leaf_37_clock _00953_ VGND VGND VPWR VPWR execute.io_mem_rd\[0\] sky130_fd_sc_hd__dfxtp_1
X_20259_ _10730_ decode.id_ex_pc_reg\[8\] _05433_ _10706_ VGND VGND VPWR VPWR _05445_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_129_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27855_ clknet_leaf_321_clock _00884_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_129_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2360 decode.regfile.registers_2\[23\] VGND VGND VPWR VPWR net2587 sky130_fd_sc_hd__dlygate4sd3_1
X_14820_ _10787_ _10767_ VGND VGND VPWR VPWR _10863_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26806_ _09408_ _09763_ VGND VGND VPWR VPWR _09774_ sky130_fd_sc_hd__nand2_1
Xhold2371 decode.regfile.registers_20\[24\] VGND VGND VPWR VPWR net2598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2382 decode.regfile.registers_9\[15\] VGND VGND VPWR VPWR net2609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2393 _10675_ VGND VGND VPWR VPWR net2620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27786_ clknet_leaf_322_clock _00815_ VGND VGND VPWR VPWR memory.io_wb_readdata\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24998_ _08703_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__clkbuf_4
Xhold1670 fetch.bht.bhtTable_target_pc\[0\]\[11\] VGND VGND VPWR VPWR net1897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29525_ clknet_leaf_265_clock _02538_ VGND VGND VPWR VPWR decode.regfile.registers_8\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1681 fetch.bht.bhtTable_target_pc\[15\]\[28\] VGND VGND VPWR VPWR net1908 sky130_fd_sc_hd__dlygate4sd3_1
X_14751_ _10791_ _10792_ _10790_ VGND VGND VPWR VPWR _10794_ sky130_fd_sc_hd__o21ai_1
X_26737_ net859 _09723_ _09734_ _09730_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23949_ net773 _08107_ _06156_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__mux2_1
Xhold1692 fetch.bht.bhtTable_tag\[9\]\[23\] VGND VGND VPWR VPWR net1919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13702_ _10052_ VGND VGND VPWR VPWR _10053_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17470_ decode.regfile.registers_18\[17\] _10924_ _12569_ _11023_ _11008_ VGND VGND
+ VPWR VPWR _13418_ sky130_fd_sc_hd__o2111a_1
X_29456_ clknet_leaf_261_clock _02469_ VGND VGND VPWR VPWR decode.regfile.registers_6\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14682_ decode.id_ex_pc_reg\[25\] VGND VGND VPWR VPWR _10725_ sky130_fd_sc_hd__inv_2
X_26668_ net1717 _09692_ _09694_ _09688_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28407_ clknet_leaf_113_clock _01420_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_4
X_16421_ _12387_ _11371_ _10646_ _11298_ _12388_ VGND VGND VPWR VPWR _12389_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_129_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25619_ _08918_ _09069_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__nand2_1
X_13633_ _09992_ VGND VGND VPWR VPWR _09993_ sky130_fd_sc_hd__buf_4
X_29387_ clknet_leaf_258_clock _02400_ VGND VGND VPWR VPWR decode.regfile.registers_4\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26599_ net2642 _09649_ _09654_ _09648_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19140_ _04244_ _04433_ _04435_ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_17_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28338_ clknet_leaf_221_clock _01351_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16352_ decode.regfile.registers_7\[27\] _11465_ _11466_ decode.regfile.registers_6\[27\]
+ _11166_ VGND VGND VPWR VPWR _12322_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_94_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13564_ decode.io_wb_rd\[2\] VGND VGND VPWR VPWR _09929_ sky130_fd_sc_hd__buf_6
XFILLER_0_183_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_229_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15303_ decode.regfile.registers_1\[1\] _11116_ _11137_ _11157_ VGND VGND VPWR VPWR
+ _11299_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_229_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19071_ _04365_ _04368_ _04269_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_229_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28269_ clknet_leaf_64_clock _01291_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16283_ _11143_ _11035_ _12254_ VGND VGND VPWR VPWR _12255_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18022_ _10603_ _12615_ _03411_ _03412_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__o32a_1
X_15234_ _10989_ _10976_ _10955_ _11093_ VGND VGND VPWR VPWR _11231_ sky130_fd_sc_hd__and4_1
XFILLER_0_151_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15165_ _11044_ decode.regfile.registers_4\[0\] _10648_ _10630_ _11084_ VGND VGND
+ VPWR VPWR _11162_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_50_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14116_ _10128_ _10286_ VGND VGND VPWR VPWR _10325_ sky130_fd_sc_hd__nand2_1
X_19973_ _03588_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__clkbuf_4
X_15096_ _11092_ VGND VGND VPWR VPWR _11093_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18924_ _04214_ _03854_ _04215_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__and4_1
X_14047_ net2368 _10244_ _10284_ _10275_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18855_ _04149_ _04152_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17806_ _12585_ _03205_ _03206_ _03207_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_98_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18786_ _04083_ _04084_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__nand2_1
X_15998_ _11976_ _11486_ _11977_ VGND VGND VPWR VPWR _11978_ sky130_fd_sc_hd__a21o_1
XFILLER_0_221_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_206_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17737_ _02986_ decode.regfile.registers_26\[23\] _13002_ _13484_ _02987_ VGND VGND
+ VPWR VPWR _03141_ sky130_fd_sc_hd__o2111a_1
Xclkbuf_leaf_161_clock clknet_5_24__leaf_clock VGND VGND VPWR VPWR clknet_leaf_161_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14949_ _10976_ VGND VGND VPWR VPWR _10977_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17668_ net600 _12872_ _03032_ _03072_ _03073_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__o221a_1
X_19407_ _04291_ _04420_ _04695_ _04345_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_35_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16619_ _10611_ _10618_ _12583_ VGND VGND VPWR VPWR _12584_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_214_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17599_ decode.regfile.registers_7\[20\] _12610_ _12623_ decode.regfile.registers_6\[20\]
+ _12843_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_163_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_176_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_176_clock
+ sky130_fd_sc_hd__clkbuf_8
X_19338_ _04345_ _04629_ _04242_ _04442_ _04610_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_156_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19269_ _04401_ _04560_ _04561_ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21300_ net1450 _10881_ _06157_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22280_ _06874_ _06623_ _06628_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21231_ csr.io_mem_pc\[12\] VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__buf_2
XFILLER_0_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold200 decode.regfile.registers_31\[12\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 decode.regfile.registers_31\[15\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold222 decode.control.io_funct7\[1\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 decode.regfile.registers_27\[5\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 decode.regfile.registers_3\[8\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold255 decode.regfile.registers_27\[2\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
X_21162_ _06075_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold266 decode.regfile.registers_27\[6\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold277 decode.regfile.registers_21\[29\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold288 decode.regfile.registers_1\[29\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
X_20113_ _05309_ _05323_ _05314_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__nand3_1
XFILLER_0_229_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_114_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_114_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold299 csr._mcycle_T_2\[25\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkbuf_2
X_21093_ csr.mtie csr.ie csr.mtip _09924_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25970_ _08966_ _09267_ VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20044_ decode.id_ex_imm_reg\[5\] _10704_ _05264_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__o21ai_2
X_24921_ csr._mcycle_T_3\[41\] csr._mcycle_T_3\[40\] csr._mcycle_T_3\[39\] _08656_
+ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__and4_1
XFILLER_0_147_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27640_ clknet_leaf_155_clock _00669_ VGND VGND VPWR VPWR execute.io_reg_pc\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_24852_ _06130_ net2073 _08607_ VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_129_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_129_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23803_ _08055_ net1822 _07952_ VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__mux2_1
X_27571_ clknet_leaf_161_clock _00600_ VGND VGND VPWR VPWR csr.io_mem_pc\[12\] sky130_fd_sc_hd__dfxtp_4
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24783_ _08076_ net1949 _08574_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__mux2_1
X_21995_ net2006 _06601_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_124_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29310_ clknet_leaf_244_clock _02323_ VGND VGND VPWR VPWR decode.regfile.registers_2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26522_ net1920 _09605_ _09610_ _09608_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__o211a_1
XANTENNA_128 _10638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23734_ _08018_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_139 _12650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20946_ _05954_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29241_ clknet_leaf_175_clock _02254_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_26453_ decode.regfile.registers_14\[26\] _09561_ _09570_ _09567_ VGND VGND VPWR
+ VPWR _02729_ sky130_fd_sc_hd__o211a_1
X_23665_ net1038 _10772_ _07972_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__mux2_1
X_20877_ _05858_ _09956_ net34 VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__and3_1
XFILLER_0_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25404_ _08905_ VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_27_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29172_ clknet_leaf_168_clock _02185_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_22616_ net2781 net1512 _07185_ _07187_ _06336_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_154_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23596_ _06126_ net1944 _07941_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__mux2_1
X_26384_ _09441_ _09490_ VGND VGND VPWR VPWR _09530_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28123_ clknet_leaf_90_clock _01145_ VGND VGND VPWR VPWR csr.minstret\[28\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_153_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25335_ _08898_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__clkbuf_1
X_22547_ csr._minstret_T_3\[33\] csr._minstret_T_3\[32\] csr.minstret\[31\] _06420_
+ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_23_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28054_ clknet_leaf_200_clock _01076_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_25266_ _08105_ net1737 _09906_ VGND VGND VPWR VPWR _08863_ sky130_fd_sc_hd__mux2_1
X_22478_ fetch.bht.bhtTable_target_pc\[8\]\[0\] fetch.bht.bhtTable_target_pc\[9\]\[0\]
+ fetch.bht.bhtTable_target_pc\[10\]\[0\] fetch.bht.bhtTable_target_pc\[11\]\[0\]
+ _07069_ _07072_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_224_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27005_ clknet_leaf_337_clock _00034_ VGND VGND VPWR VPWR decode.regfile.registers_22\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24217_ _08111_ net2249 _06251_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__mux2_1
X_21429_ _06229_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_62_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25197_ _08827_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24148_ _08247_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28956_ clknet_leaf_181_clock _01969_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24079_ net1079 execute.io_target_pc\[27\] _07991_ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16970_ decode.regfile.registers_9\[5\] _12776_ _12604_ _12532_ _12598_ VGND VGND
+ VPWR VPWR _12930_ sky130_fd_sc_hd__a41o_1
XFILLER_0_229_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27907_ clknet_leaf_18_clock _00936_ VGND VGND VPWR VPWR csr._mcycle_T_2\[28\] sky130_fd_sc_hd__dfxtp_4
X_15921_ decode.regfile.registers_21\[15\] _11062_ _11100_ _11229_ _11902_ VGND VGND
+ VPWR VPWR _11903_ sky130_fd_sc_hd__o311a_1
XFILLER_0_21_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28887_ clknet_leaf_117_clock _01900_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18640_ _03912_ _03924_ _03936_ _03937_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__a311o_1
X_15852_ _11493_ decode.regfile.registers_24\[14\] VGND VGND VPWR VPWR _11835_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27838_ clknet_leaf_326_clock _00867_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2190 decode.regfile.registers_22\[25\] VGND VGND VPWR VPWR net2417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14803_ _10764_ _10809_ _10681_ VGND VGND VPWR VPWR _10846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18571_ execute.io_reg_pc\[23\] _03777_ _03665_ net115 _03869_ VGND VGND VPWR VPWR
+ _03870_ sky130_fd_sc_hd__o221a_1
X_15783_ decode.regfile.registers_2\[12\] _10647_ _11149_ _11152_ _11767_ VGND VGND
+ VPWR VPWR _11768_ sky130_fd_sc_hd__o311a_1
X_27769_ clknet_leaf_324_clock _00798_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17522_ decode.regfile.registers_13\[18\] _12775_ _13467_ _13468_ _12664_ VGND VGND
+ VPWR VPWR _13469_ sky130_fd_sc_hd__a221o_1
X_29508_ clknet_leaf_267_clock _02521_ VGND VGND VPWR VPWR decode.regfile.registers_8\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14734_ csr.io_mem_pc\[30\] VGND VGND VPWR VPWR _10777_ sky130_fd_sc_hd__buf_4
XFILLER_0_118_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_93_clock clknet_5_10__leaf_clock VGND VGND VPWR VPWR clknet_leaf_93_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_157_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17453_ decode.regfile.registers_21\[16\] _12716_ _13378_ _13401_ _12806_ VGND VGND
+ VPWR VPWR _13402_ sky130_fd_sc_hd__o221a_1
X_29439_ clknet_leaf_248_clock _02452_ VGND VGND VPWR VPWR decode.regfile.registers_6\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14665_ _10705_ execute.io_target_pc\[5\] _10707_ execute.io_target_pc\[9\] VGND
+ VGND VPWR VPWR _10708_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_131_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16404_ _10991_ _11065_ _11080_ _11232_ decode.regfile.registers_23\[28\] VGND VGND
+ VPWR VPWR _12373_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13616_ _09960_ VGND VGND VPWR VPWR _09977_ sky130_fd_sc_hd__clkbuf_4
X_17384_ _12694_ _13332_ _13333_ _13334_ VGND VGND VPWR VPWR _13335_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14596_ _10638_ VGND VGND VPWR VPWR _10639_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19123_ _04269_ _04417_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_172_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16335_ _11679_ decode.regfile.registers_27\[26\] _11869_ VGND VGND VPWR VPWR _12306_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_55_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13547_ _09914_ _09894_ _09917_ net394 VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19054_ _04246_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__clkbuf_4
X_16266_ _11493_ decode.regfile.registers_24\[25\] VGND VGND VPWR VPWR _12238_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_11_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18005_ _12515_ _03399_ _03400_ _03401_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__a31o_1
XFILLER_0_180_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15217_ _11106_ _11212_ _11213_ VGND VGND VPWR VPWR _11214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16197_ _10957_ decode.regfile.registers_22\[23\] _11450_ _10978_ _10990_ VGND VGND
+ VPWR VPWR _12171_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_31_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_199_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15148_ _11144_ VGND VGND VPWR VPWR _11145_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_207_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_207_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19956_ _10748_ _03599_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__nor2_1
X_15079_ _11049_ VGND VGND VPWR VPWR _11076_ sky130_fd_sc_hd__clkbuf_4
X_18907_ _03898_ _03899_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_203_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19887_ _04856_ _05134_ _05156_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_leaf_46_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_46_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_203_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18838_ _04133_ _03914_ _03687_ decode.id_ex_rs1_data_reg\[9\] _04136_ VGND VGND
+ VPWR VPWR _04137_ sky130_fd_sc_hd__o221a_4
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18769_ memory.csr_read_data_out_reg\[6\] _10010_ _09997_ VGND VGND VPWR VPWR _04068_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20800_ _05874_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21780_ _06453_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20731_ decode.id_ex_rs1_data_reg\[23\] VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23450_ net5 _07846_ _07860_ _07851_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__o211a_1
X_20662_ _05788_ _05790_ _03595_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22401_ _06995_ _06675_ _06686_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23381_ fetch.bht.bhtTable_target_pc\[12\]\[29\] fetch.bht.bhtTable_target_pc\[13\]\[29\]
+ fetch.bht.bhtTable_target_pc\[14\]\[29\] fetch.bht.bhtTable_target_pc\[15\]\[29\]
+ _07068_ _07656_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__mux4_1
XFILLER_0_163_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20593_ csr.minstret\[21\] _05574_ _05586_ csr.mcycle\[21\] VGND VGND VPWR VPWR _05732_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25120_ _08788_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__clkbuf_1
X_22332_ _06920_ _06922_ _06924_ _06926_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_6_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25051_ csr.mcycle\[20\] _03554_ csr.mcycle\[21\] _08644_ VGND VGND VPWR VPWR _08747_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_104_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22263_ fetch.bht.bhtTable_tag\[14\]\[17\] fetch.bht.bhtTable_tag\[15\]\[17\] _06809_
+ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24002_ _08172_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__clkbuf_1
X_21214_ net879 _06101_ _09912_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__mux2_1
X_22194_ fetch.bht.bhtTable_tag\[12\]\[5\] fetch.bht.bhtTable_tag\[13\]\[5\] fetch.bht.bhtTable_tag\[14\]\[5\]
+ fetch.bht.bhtTable_tag\[15\]\[5\] _06700_ _06651_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_203_Right_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28810_ clknet_leaf_98_clock _01823_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21145_ _06062_ _06058_ net2097 VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__and3_1
X_29790_ clknet_leaf_310_clock _02803_ VGND VGND VPWR VPWR decode.regfile.registers_17\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_28741_ clknet_leaf_135_clock _01754_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25953_ net2062 _09256_ _09269_ _09264_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__o211a_1
X_21076_ _06024_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20027_ _05248_ _05249_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__and2b_1
X_24904_ net1898 _08649_ _08650_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__o21a_1
X_28672_ clknet_leaf_171_clock _01685_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25884_ net2461 _09226_ _09229_ _09222_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__o211a_1
X_27623_ clknet_leaf_48_clock _00652_ VGND VGND VPWR VPWR execute.io_reg_pc\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24835_ _06113_ net1400 _08422_ VGND VGND VPWR VPWR _08605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27554_ clknet_leaf_25_clock _00583_ VGND VGND VPWR VPWR execute.io_mem_regwrite
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24766_ _08060_ net1701 _08563_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__mux2_1
X_21978_ csr._mcycle_T_2\[12\] _06587_ _06591_ _06592_ VGND VGND VPWR VPWR _01232_
+ sky130_fd_sc_hd__o211a_1
Xrebuffer70 _03710_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_1
X_26505_ net1699 _09592_ _09600_ _09595_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__o211a_1
Xrebuffer81 _03751_ VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_189_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23717_ _08009_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer92 _11069_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__buf_1
XFILLER_0_95_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20929_ _09955_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27485_ clknet_leaf_24_clock _00514_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_1
X_24697_ _08532_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29224_ clknet_leaf_120_clock _02237_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26436_ net2326 _09548_ _09560_ _09553_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__o211a_1
X_14450_ net435 _10506_ _10518_ _10509_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__o211a_1
X_23648_ _07960_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29155_ clknet_leaf_221_clock _02168_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26367_ _09424_ _09515_ VGND VGND VPWR VPWR _09521_ sky130_fd_sc_hd__nand2_1
X_14381_ _10036_ _10474_ VGND VGND VPWR VPWR _10479_ sky130_fd_sc_hd__nand2_1
X_23579_ _07934_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_1086 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28106_ clknet_leaf_75_clock _01128_ VGND VGND VPWR VPWR csr.minstret\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_70_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16120_ _10981_ VGND VGND VPWR VPWR _12096_ sky130_fd_sc_hd__buf_2
X_25318_ _08889_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29086_ clknet_leaf_72_clock _02099_ VGND VGND VPWR VPWR csr._mcycle_T_3\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26298_ _09430_ _09472_ VGND VGND VPWR VPWR _09481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_228_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28037_ clknet_leaf_183_clock _01059_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16051_ _11084_ _11297_ _11534_ decode.regfile.registers_6\[19\] _12028_ VGND VGND
+ VPWR VPWR _12029_ sky130_fd_sc_hd__o221a_1
X_25249_ _08854_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15002_ _10599_ VGND VGND VPWR VPWR _11013_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19810_ _03810_ _03639_ _04667_ _03814_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16953_ _12516_ _12911_ _12912_ _12913_ VGND VGND VPWR VPWR _12914_ sky130_fd_sc_hd__a31o_1
X_19741_ _04931_ _04929_ _05015_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__o21bai_2
X_28939_ clknet_leaf_93_clock _01952_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15904_ _11881_ _11884_ _11885_ VGND VGND VPWR VPWR _11886_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_218_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19672_ _04508_ _04492_ _04536_ _04950_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__a31o_1
X_16884_ _11017_ _12502_ _12509_ decode.regfile.registers_8\[3\] _12725_ VGND VGND
+ VPWR VPWR _12846_ sky130_fd_sc_hd__o32a_1
XFILLER_0_95_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18623_ _03889_ decode.id_ex_imm_reg\[18\] VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__and2_1
X_15835_ _11818_ decode.regfile.registers_17\[13\] _11356_ VGND VGND VPWR VPWR _11819_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18554_ _03839_ _03851_ _03852_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__and3_1
X_15766_ decode.regfile.registers_25\[11\] _11333_ _11336_ decode.regfile.registers_24\[11\]
+ VGND VGND VPWR VPWR _11752_ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17505_ _13451_ net2272 _13097_ VGND VGND VPWR VPWR _13452_ sky130_fd_sc_hd__o21a_1
XFILLER_0_213_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14717_ csr.io_mem_pc\[26\] VGND VGND VPWR VPWR _10760_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_190_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18485_ _03734_ _03782_ _03783_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_190_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ _11344_ net441 _11645_ _11684_ _11249_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17436_ decode.regfile.registers_2\[16\] _12634_ _12628_ _13384_ VGND VGND VPWR VPWR
+ _13385_ sky130_fd_sc_hd__o211ai_4
X_14648_ _10688_ _10689_ execute.io_target_pc\[4\] _10690_ VGND VGND VPWR VPWR _10691_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_16_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_17 _04655_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_28 _08939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17367_ _11016_ _12539_ _12502_ decode.regfile.registers_7\[14\] _12644_ VGND VGND
+ VPWR VPWR _13318_ sky130_fd_sc_hd__o32a_1
XANTENNA_39 _10101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14579_ _10604_ decode.id_ex_ex_rd_reg\[1\] decode.id_ex_ex_rd_reg\[3\] _10606_ _10621_
+ VGND VGND VPWR VPWR _10622_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19106_ _04398_ _04399_ _04400_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16318_ decode.regfile.registers_11\[26\] _11364_ _12277_ _12288_ VGND VGND VPWR
+ VPWR _12289_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_67_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17298_ _13250_ decode.regfile.registers_24\[12\] _13170_ _13083_ _12862_ VGND VGND
+ VPWR VPWR _13251_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19037_ _04249_ _04335_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_209_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16249_ decode.regfile.registers_16\[24\] _11123_ _12205_ _12221_ VGND VGND VPWR
+ VPWR _12222_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_209_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput102 net102 VGND VGND VPWR VPWR io_memory_address[11] sky130_fd_sc_hd__clkbuf_4
Xoutput113 net113 VGND VGND VPWR VPWR io_memory_address[21] sky130_fd_sc_hd__clkbuf_4
Xoutput124 net124 VGND VGND VPWR VPWR io_memory_address[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput135 net135 VGND VGND VPWR VPWR io_memory_write sky130_fd_sc_hd__clkbuf_4
Xoutput146 net146 VGND VGND VPWR VPWR io_memory_write_data[19] sky130_fd_sc_hd__clkbuf_4
Xoutput157 net157 VGND VGND VPWR VPWR io_memory_write_data[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_8 _01445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19939_ _05203_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22950_ net92 _07348_ _07399_ _03580_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__a211o_1
XFILLER_0_177_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21901_ csr._mcycle_T_2\[19\] _06521_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22881_ _07337_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24620_ _08492_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__clkbuf_1
X_21832_ csr.io_mret_vector\[0\] csr.io_mem_pc\[0\] _06040_ VGND VGND VPWR VPWR _06491_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21763_ _06444_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__clkbuf_1
X_24551_ _08111_ net2092 _09902_ VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23502_ net89 _07889_ _07891_ _07879_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__o211a_1
X_20714_ _05813_ decode.id_ex_rs1_data_reg\[16\] VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__nand2_1
X_27270_ clknet_leaf_14_clock _00299_ VGND VGND VPWR VPWR decode.regfile.registers_30\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_24482_ _08109_ net1429 _08411_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__mux2_1
X_21694_ _05691_ csr.minstret\[16\] _06391_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26221_ net195 VGND VGND VPWR VPWR _09434_ sky130_fd_sc_hd__buf_4
X_20645_ csr.minstret\[29\] _05572_ _05582_ csr.mcycle\[29\] _05775_ VGND VGND VPWR
+ VPWR _05776_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23433_ net28 _07846_ _07850_ _07851_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23364_ _06795_ _07783_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__nand2_1
X_26152_ _09385_ _09374_ VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20576_ _05717_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25103_ _06119_ net1606 _08778_ VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22315_ fetch.bht.bhtTable_tag\[8\]\[0\] fetch.bht.bhtTable_tag\[9\]\[0\] _06643_
+ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23295_ fetch.bht.bhtTable_target_pc\[8\]\[23\] fetch.bht.bhtTable_target_pc\[9\]\[23\]
+ fetch.bht.bhtTable_target_pc\[10\]\[23\] fetch.bht.bhtTable_target_pc\[11\]\[23\]
+ _07708_ _07103_ VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26083_ net556 _09343_ _09344_ _09333_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_186_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22246_ _06684_ _06840_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_186_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25034_ _08736_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29911_ clknet_leaf_340_clock _02924_ VGND VGND VPWR VPWR decode.regfile.registers_20\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29842_ clknet_leaf_299_clock _02855_ VGND VGND VPWR VPWR decode.regfile.registers_18\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_22177_ _06624_ _06771_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21128_ _06056_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29773_ clknet_leaf_295_clock _02786_ VGND VGND VPWR VPWR decode.regfile.registers_16\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_26985_ _10135_ _09838_ VGND VGND VPWR VPWR _09876_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28724_ clknet_leaf_117_clock _01737_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13950_ _10097_ _10223_ VGND VGND VPWR VPWR _10229_ sky130_fd_sc_hd__nand2_1
X_25936_ net937 _09256_ _09259_ _09250_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__o211a_1
X_21059_ execute.csr_read_data_out_reg\[18\] _06014_ _06010_ VGND VGND VPWR VPWR _06016_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_145_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28655_ clknet_leaf_111_clock _01668_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13881_ _10131_ VGND VGND VPWR VPWR _10188_ sky130_fd_sc_hd__clkbuf_4
X_25867_ net2371 _09213_ _09219_ _09209_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27606_ clknet_leaf_151_clock _00635_ VGND VGND VPWR VPWR execute.io_target_pc\[15\]
+ sky130_fd_sc_hd__dfxtp_4
X_15620_ _11344_ net434 _11572_ _11609_ _11249_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__o221a_1
X_24818_ _08561_ VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__clkbuf_8
X_28586_ clknet_leaf_98_clock _01599_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25798_ _08945_ _09179_ VGND VGND VPWR VPWR _09180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_207 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27537_ clknet_leaf_155_clock _00566_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_2
X_15551_ decode.regfile.registers_3\[6\] _11152_ _11537_ _11541_ VGND VGND VPWR VPWR
+ _11542_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_218 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24749_ _08111_ net2219 _06283_ VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_229 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14502_ net775 _10507_ _10547_ _10546_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18270_ net490 _03599_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27468_ clknet_leaf_53_clock _00497_ VGND VGND VPWR VPWR csr.io_csr_address\[2\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_13_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ decode.regfile.registers_16\[4\] _11359_ _11457_ _11474_ _11126_ VGND VGND
+ VPWR VPWR _11475_ sky130_fd_sc_hd__o221a_1
XFILLER_0_189_1159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29207_ clknet_leaf_240_clock _02220_ VGND VGND VPWR VPWR fetch.btb.btbTable\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_17221_ _12667_ VGND VGND VPWR VPWR _13176_ sky130_fd_sc_hd__buf_2
X_26419_ _09400_ _09545_ VGND VGND VPWR VPWR _09551_ sky130_fd_sc_hd__nand2_1
X_14433_ net580 _10506_ _10508_ _10509_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27399_ clknet_leaf_29_clock _00428_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29138_ clknet_leaf_78_clock _02151_ VGND VGND VPWR VPWR csr.mcycle\[22\] sky130_fd_sc_hd__dfxtp_1
X_17152_ decode.regfile.registers_6\[9\] _10602_ _12626_ _12645_ VGND VGND VPWR VPWR
+ _13108_ sky130_fd_sc_hd__o31a_1
XFILLER_0_135_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput15 io_fetch_data[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14364_ net553 _10463_ _10469_ _10468_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__o211a_1
Xinput26 io_fetch_data[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput37 io_memory_read_data[12] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
XFILLER_0_135_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16103_ _12079_ decode.regfile.registers_18\[20\] _11455_ VGND VGND VPWR VPWR _12080_
+ sky130_fd_sc_hd__mux2_1
Xinput48 io_memory_read_data[22] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
Xinput59 io_memory_read_data[3] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_2
X_29069_ clknet_leaf_200_clock _02082_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17083_ _12519_ VGND VGND VPWR VPWR _13041_ sky130_fd_sc_hd__clkbuf_2
X_14295_ net698 _10419_ _10429_ _10427_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16034_ _11489_ decode.regfile.registers_28\[18\] decode.regfile.registers_29\[18\]
+ _11255_ _11245_ VGND VGND VPWR VPWR _12013_ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17985_ _12934_ _10592_ _12558_ decode.regfile.registers_0\[30\] VGND VGND VPWR VPWR
+ _03382_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_200_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16936_ decode.regfile.registers_13\[4\] _12659_ _12670_ VGND VGND VPWR VPWR _12897_
+ sky130_fd_sc_hd__o21ai_1
X_19724_ _03894_ _04195_ _04998_ _04496_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_196_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16867_ _10591_ _10605_ _10934_ _10607_ VGND VGND VPWR VPWR _12829_ sky130_fd_sc_hd__nand4_4
X_19655_ _04192_ _04929_ _04931_ _04933_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_0_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18606_ net108 _03665_ _03904_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__o21ai_2
X_15818_ decode.regfile.registers_5\[13\] _11178_ _11138_ VGND VGND VPWR VPWR _11802_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_133_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19586_ _04198_ _04865_ net213 _04867_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16798_ decode.regfile.registers_27\[1\] _12507_ _12520_ _12495_ _12761_ VGND VGND
+ VPWR VPWR _12762_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_9_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18537_ decode.id_ex_rs2_data_reg\[25\] _03747_ _03833_ _03764_ VGND VGND VPWR VPWR
+ _03836_ sky130_fd_sc_hd__o22a_1
X_15749_ decode.regfile.registers_5\[11\] _11291_ _11733_ _11734_ VGND VGND VPWR VPWR
+ _11735_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_181_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18468_ _03639_ _03705_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17419_ _13339_ _13365_ _13366_ _13368_ VGND VGND VPWR VPWR _13369_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_151_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18399_ _03693_ _03695_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__nor3_4
XFILLER_0_43_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20430_ _05587_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__buf_4
XFILLER_0_145_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20361_ _03737_ _03741_ _03755_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22100_ _06694_ _06690_ _06627_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23080_ fetch.bht.bhtTable_target_pc\[12\]\[11\] fetch.bht.bhtTable_target_pc\[13\]\[11\]
+ fetch.bht.bhtTable_target_pc\[14\]\[11\] fetch.bht.bhtTable_target_pc\[15\]\[11\]
+ _07069_ _07111_ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_228_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20292_ _10681_ decode.id_ex_pc_reg\[16\] _10806_ _05462_ VGND VGND VPWR VPWR _05470_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_110_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22031_ _00002_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_227_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_181_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26770_ _10245_ _09753_ VGND VGND VPWR VPWR _09754_ sky130_fd_sc_hd__nand2_1
X_23982_ net1672 execute.io_target_pc\[12\] _08153_ VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__mux2_1
X_25721_ net1555 _09125_ _09135_ _09129_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__o211a_1
X_22933_ net89 _07343_ _07344_ _07383_ _06566_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_108_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28440_ clknet_leaf_54_clock _01453_ VGND VGND VPWR VPWR decode.control.io_funct7\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_196_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25652_ _08952_ _09092_ VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22864_ _07328_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_140_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1057 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24603_ net1257 execute.io_target_pc\[23\] _09897_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28371_ clknet_leaf_207_clock _01384_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_21815_ _06316_ _06472_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_80_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25583_ _08958_ _09049_ VGND VGND VPWR VPWR _09056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22795_ _07292_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27322_ clknet_leaf_34_clock _00351_ VGND VGND VPWR VPWR decode.id_ex_ex_rs1_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_4
X_24534_ _08448_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21746_ _06435_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27253_ clknet_leaf_30_clock _00282_ VGND VGND VPWR VPWR decode.regfile.registers_30\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_24465_ _08412_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__clkbuf_1
X_21677_ _10019_ _06382_ _06384_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26204_ _09422_ _09413_ VGND VGND VPWR VPWR _09423_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23416_ fetch.bht.bhtTable_target_pc\[6\]\[31\] fetch.bht.bhtTable_target_pc\[7\]\[31\]
+ _07066_ VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20628_ csr.minstret\[26\] _05573_ _05585_ csr.mcycle\[26\] VGND VGND VPWR VPWR _05762_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27184_ clknet_leaf_6_clock _00213_ VGND VGND VPWR VPWR decode.regfile.registers_28\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_3__f_clock clknet_2_0_0_clock VGND VGND VPWR VPWR clknet_5_3__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_24396_ net754 VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26135_ _09025_ _09374_ VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23347_ csr._csr_read_data_T_8\[26\] _07416_ csr.io_mret_vector\[26\] _07621_ _07773_
+ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__o221a_1
X_20559_ csr._csr_read_data_T_8\[16\] _05622_ _05698_ _05700_ _05702_ VGND VGND VPWR
+ VPWR _05703_ sky130_fd_sc_hd__a221o_2
XFILLER_0_46_1115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14080_ net2458 _10302_ _10305_ _10304_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__o211a_1
X_26066_ _08912_ _09330_ VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__nand2_1
X_23278_ fetch.bht.bhtTable_target_pc\[8\]\[22\] fetch.bht.bhtTable_target_pc\[9\]\[22\]
+ fetch.bht.bhtTable_target_pc\[10\]\[22\] fetch.bht.bhtTable_target_pc\[11\]\[22\]
+ _07708_ _07103_ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__mux4_1
XFILLER_0_104_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25017_ csr.mcycle\[8\] csr.mcycle\[10\] csr.mcycle\[9\] _08635_ VGND VGND VPWR VPWR
+ _08725_ sky130_fd_sc_hd__and4_1
XFILLER_0_219_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22229_ _06823_ _06628_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29825_ clknet_leaf_307_clock _02838_ VGND VGND VPWR VPWR decode.regfile.registers_18\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17770_ decode.regfile.registers_21\[24\] _12716_ _03148_ _03172_ _13164_ VGND VGND
+ VPWR VPWR _03173_ sky130_fd_sc_hd__o221a_1
X_14982_ _10964_ _10951_ VGND VGND VPWR VPWR _11000_ sky130_fd_sc_hd__nor2_1
X_26968_ net1995 _09866_ _09867_ _09865_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__o211a_1
X_29756_ clknet_leaf_310_clock _02769_ VGND VGND VPWR VPWR decode.regfile.registers_16\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16721_ _12685_ VGND VGND VPWR VPWR _12686_ sky130_fd_sc_hd__buf_2
X_28707_ clknet_leaf_131_clock _01720_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13933_ net2313 _10213_ _10218_ _10219_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25919_ _09128_ VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__clkbuf_4
X_29687_ clknet_leaf_282_clock _02700_ VGND VGND VPWR VPWR decode.regfile.registers_13\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26899_ net2513 _09822_ _09827_ _09825_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19440_ _10909_ _03636_ _09954_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__and3b_2
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28638_ clknet_leaf_176_clock _01651_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_16652_ _12522_ _12616_ _12547_ VGND VGND VPWR VPWR _12617_ sky130_fd_sc_hd__and3_2
XFILLER_0_199_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13864_ net2149 _10167_ _10178_ _10175_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_18_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15603_ _10651_ _10625_ _11054_ _11592_ VGND VGND VPWR VPWR _11593_ sky130_fd_sc_hd__o31a_1
XFILLER_0_92_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19371_ _04144_ _04642_ _04645_ _04660_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__a31oi_1
X_28569_ clknet_leaf_201_clock _01582_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16583_ _12547_ VGND VGND VPWR VPWR _12548_ sky130_fd_sc_hd__clkbuf_4
X_13795_ _10131_ VGND VGND VPWR VPWR _10132_ sky130_fd_sc_hd__clkbuf_4
X_18322_ _03626_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15534_ _11403_ _11523_ _11524_ _11525_ VGND VGND VPWR VPWR _11526_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18253_ net66 _10971_ _10757_ _10908_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__or4_1
X_15465_ decode.regfile.registers_1\[4\] _11115_ _11056_ _11108_ VGND VGND VPWR VPWR
+ _11458_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17204_ decode.regfile.registers_16\[10\] _12575_ _13140_ _13158_ VGND VGND VPWR
+ VPWR _13159_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14416_ net496 _10490_ _10498_ _10494_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18184_ decode.control.io_funct3\[2\] _10944_ _10941_ decode.control.io_funct7\[5\]
+ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15396_ decode.regfile.registers_20\[2\] _11102_ _11327_ _11390_ VGND VGND VPWR VPWR
+ _11391_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17135_ _13091_ _12706_ decode.regfile.registers_27\[8\] _13050_ VGND VGND VPWR VPWR
+ _13092_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14347_ net1297 _10447_ _10458_ _10453_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold607 fetch.bht.bhtTable_target_pc\[1\]\[17\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold618 fetch.bht.bhtTable_target_pc\[1\]\[21\] VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold629 fetch.bht.bhtTable_target_pc\[3\]\[17\] VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__dlygate4sd3_1
X_17066_ decode.regfile.registers_9\[7\] _12607_ _12599_ VGND VGND VPWR VPWR _13024_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14278_ _10418_ VGND VGND VPWR VPWR _10419_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16017_ _11191_ _11097_ _11375_ decode.regfile.registers_4\[18\] _11995_ VGND VGND
+ VPWR VPWR _11996_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_223_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_223_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 csr._csr_read_data_T_8\[7\] VGND VGND VPWR VPWR net2235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2019 fetch.bht.bhtTable_tag\[5\]\[18\] VGND VGND VPWR VPWR net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1307 fetch.bht.bhtTable_target_pc\[5\]\[6\] VGND VGND VPWR VPWR net1534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 decode.regfile.registers_14\[3\] VGND VGND VPWR VPWR net1545 sky130_fd_sc_hd__dlygate4sd3_1
X_17968_ _03364_ _03365_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__or2_1
Xhold1329 fetch.bht.bhtTable_tag\[3\]\[0\] VGND VGND VPWR VPWR net1556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19707_ _04944_ _04352_ _04983_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16919_ _12879_ VGND VGND VPWR VPWR _12880_ sky130_fd_sc_hd__buf_2
X_17899_ _12967_ _03296_ _03297_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__a31o_1
X_19638_ _04205_ _03918_ _04253_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19569_ _04056_ _04296_ _04301_ _04305_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__or4_1
XFILLER_0_177_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21600_ net1064 csr.minstret\[1\] _06323_ _06326_ _06327_ VGND VGND VPWR VPWR _01118_
+ sky130_fd_sc_hd__a311oi_1
XFILLER_0_34_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22580_ _06578_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_192_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_217_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21531_ _06285_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21462_ _06153_ net1403 _06241_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__mux2_1
X_24250_ _06217_ VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_170_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23201_ net76 _06887_ _07613_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__and3_1
X_20413_ _05571_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24181_ _08264_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__clkbuf_1
X_21393_ _06209_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23132_ execute.io_target_pc\[13\] _07346_ _07348_ _07571_ VGND VGND VPWR VPWR _07572_
+ sky130_fd_sc_hd__a211o_1
X_20344_ _05508_ _05509_ _05418_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23063_ fetch.bht.bhtTable_target_pc\[4\]\[10\] fetch.bht.bhtTable_target_pc\[5\]\[10\]
+ fetch.bht.bhtTable_target_pc\[6\]\[10\] fetch.bht.bhtTable_target_pc\[7\]\[10\]
+ _07108_ _07115_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__mux4_1
X_27940_ clknet_leaf_221_clock _00962_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20275_ _05412_ _05300_ _05457_ _03517_ _03551_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22014_ net2624 _06601_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__or2_1
X_27871_ clknet_leaf_326_clock _00900_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2520 decode.id_ex_rs1_data_reg\[17\] VGND VGND VPWR VPWR net2747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26822_ _09426_ _09776_ VGND VGND VPWR VPWR _09783_ sky130_fd_sc_hd__nand2_1
Xhold2531 decode.regfile.registers_14\[24\] VGND VGND VPWR VPWR net2758 sky130_fd_sc_hd__dlygate4sd3_1
X_29610_ clknet_leaf_276_clock _02623_ VGND VGND VPWR VPWR decode.regfile.registers_11\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2542 decode.io_id_pc\[8\] VGND VGND VPWR VPWR net2769 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2553 csr._minstret_T_3\[59\] VGND VGND VPWR VPWR net2780 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2564 decode.regfile.registers_30\[11\] VGND VGND VPWR VPWR net2791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1830 csr._mcycle_T_3\[38\] VGND VGND VPWR VPWR net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2575 decode.csr_read_reg VGND VGND VPWR VPWR net2802 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29541_ clknet_leaf_273_clock _02554_ VGND VGND VPWR VPWR decode.regfile.registers_9\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1841 fetch.bht.bhtTable_target_pc\[7\]\[7\] VGND VGND VPWR VPWR net2068 sky130_fd_sc_hd__dlygate4sd3_1
X_26753_ net2629 _09736_ _09742_ _09743_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_32_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1852 fetch.bht.bhtTable_tag\[7\]\[10\] VGND VGND VPWR VPWR net2079 sky130_fd_sc_hd__dlygate4sd3_1
X_23965_ _07959_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_32_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1863 fetch.bht.bhtTable_tag\[11\]\[2\] VGND VGND VPWR VPWR net2090 sky130_fd_sc_hd__dlygate4sd3_1
X_25704_ _08929_ _09122_ VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__nand2_1
Xhold1874 decode.regfile.registers_22\[18\] VGND VGND VPWR VPWR net2101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1885 fetch.bht.bhtTable_target_pc\[9\]\[2\] VGND VGND VPWR VPWR net2112 sky130_fd_sc_hd__dlygate4sd3_1
X_22916_ net186 _07366_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__and2_2
X_29472_ clknet_leaf_249_clock _02485_ VGND VGND VPWR VPWR decode.regfile.registers_7\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26684_ net2277 _09692_ _09703_ _09702_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__o211a_1
Xhold1896 decode.regfile.registers_5\[26\] VGND VGND VPWR VPWR net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23896_ _08117_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28423_ clknet_leaf_39_clock _01436_ VGND VGND VPWR VPWR decode.control.io_funct3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25635_ _08935_ _09079_ VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__nand2_1
X_22847_ _07319_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28354_ clknet_leaf_188_clock _01367_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_25566_ net1499 _09039_ _09045_ _09046_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__o211a_1
X_13580_ _09943_ memory.io_wb_readdata\[0\] _09944_ VGND VGND VPWR VPWR _09945_ sky130_fd_sc_hd__o21ai_2
X_22778_ _07282_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27305_ clknet_leaf_13_clock _00334_ VGND VGND VPWR VPWR decode.regfile.registers_31\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24517_ _08076_ net1511 _08439_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28285_ clknet_leaf_85_clock _01307_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[23\]
+ sky130_fd_sc_hd__dfxtp_2
X_21729_ _06425_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__clkbuf_1
X_25497_ net2738 _08995_ _09006_ _09004_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27236_ clknet_leaf_364_clock _00265_ VGND VGND VPWR VPWR decode.regfile.registers_29\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_15250_ net580 _11243_ _11246_ net505 VGND VGND VPWR VPWR _11247_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_62_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24448_ _08403_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14201_ _10373_ _10195_ _09933_ _10196_ VGND VGND VPWR VPWR _10374_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27167_ clknet_leaf_359_clock _00196_ VGND VGND VPWR VPWR decode.regfile.registers_27\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15181_ _10635_ VGND VGND VPWR VPWR _11178_ sky130_fd_sc_hd__clkbuf_4
X_24379_ _08366_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14132_ net522 _10332_ _10335_ _10328_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__o211a_1
X_26118_ _08964_ _09353_ VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27098_ clknet_leaf_349_clock _00127_ VGND VGND VPWR VPWR decode.regfile.registers_25\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14063_ net864 _10287_ _10295_ _10291_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__o211a_1
X_26049_ _08970_ _09285_ VGND VGND VPWR VPWR _09324_ sky130_fd_sc_hd__nand2_1
X_18940_ _04225_ _03705_ _03766_ _04238_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__o31a_1
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18871_ _04121_ _04169_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__or2_4
XFILLER_0_218_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29808_ clknet_leaf_295_clock _02821_ VGND VGND VPWR VPWR decode.regfile.registers_17\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_17822_ _02997_ _12767_ _12965_ decode.regfile.registers_29\[25\] _03223_ VGND VGND
+ VPWR VPWR _03224_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17753_ decode.regfile.registers_2\[24\] _12634_ _12628_ _03155_ VGND VGND VPWR VPWR
+ _03156_ sky130_fd_sc_hd__o211a_1
X_29739_ clknet_leaf_294_clock _02752_ VGND VGND VPWR VPWR decode.regfile.registers_15\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_14965_ _10989_ VGND VGND VPWR VPWR _10990_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16704_ _12668_ VGND VGND VPWR VPWR _12669_ sky130_fd_sc_hd__clkbuf_4
X_13916_ net1696 _10199_ _10209_ _10206_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17684_ decode.regfile.registers_11\[22\] _12594_ _12582_ _12550_ VGND VGND VPWR
+ VPWR _03089_ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14896_ _10932_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19423_ _04028_ _04485_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__nor2_1
X_16635_ _12599_ VGND VGND VPWR VPWR _12600_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13847_ _10036_ _10164_ VGND VGND VPWR VPWR _10169_ sky130_fd_sc_hd__nand2_1
X_16566_ _12530_ VGND VGND VPWR VPWR _12531_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19354_ _04129_ _04126_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__nand2b_2
X_13778_ _10116_ VGND VGND VPWR VPWR _10117_ sky130_fd_sc_hd__clkbuf_8
X_15517_ _11183_ VGND VGND VPWR VPWR _11509_ sky130_fd_sc_hd__clkbuf_4
X_18305_ decode.id_ex_rs2_data_reg\[18\] _03616_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__and2_1
X_19285_ _03594_ _04566_ _04578_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16497_ decode.regfile.registers_5\[31\] _11291_ _12461_ _12462_ VGND VGND VPWR VPWR
+ _12463_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_155_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18236_ csr._mcycle_T_3\[45\] csr._mcycle_T_3\[44\] csr._mcycle_T_3\[43\] csr._mcycle_T_3\[42\]
+ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__or4_1
XFILLER_0_217_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15448_ _11403_ _11438_ _11439_ _11441_ VGND VGND VPWR VPWR _11442_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_212_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18167_ _03511_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15379_ decode.regfile.registers_2\[2\] _11369_ _11297_ _11121_ _11373_ VGND VGND
+ VPWR VPWR _11374_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_128_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold404 decode.regfile.registers_27\[13\] VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__dlygate4sd3_1
X_17118_ decode.regfile.registers_17\[8\] _12580_ _12826_ _13074_ VGND VGND VPWR VPWR
+ _13075_ sky130_fd_sc_hd__o211a_1
X_18098_ _03475_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__clkbuf_1
Xhold415 decode.regfile.registers_30\[6\] VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold426 decode.regfile.registers_17\[10\] VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold437 decode.regfile.registers_28\[26\] VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold448 decode.regfile.registers_27\[28\] VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold459 decode.regfile.registers_3\[2\] VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__dlygate4sd3_1
X_17049_ net508 _12491_ _12706_ _10940_ VGND VGND VPWR VPWR _13008_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap189 _03795_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
X_20060_ decode.id_ex_imm_reg\[9\] _10706_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1104 fetch.bht.bhtTable_tag\[9\]\[8\] VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 fetch.bht.bhtTable_tag\[6\]\[4\] VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 fetch.bht.bhtTable_target_pc\[8\]\[7\] VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 fetch.bht.bhtTable_tag\[10\]\[7\] VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1148 fetch.bht.bhtTable_target_pc\[14\]\[12\] VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1159 fetch.bht.bhtTable_tag\[1\]\[17\] VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23750_ _08026_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_176_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ execute.io_reg_pc\[7\] _05915_ _05961_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22701_ net2736 _07235_ _07239_ _07234_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23681_ _07989_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ _05925_ _05921_ net63 VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25420_ net486 _08951_ _08957_ _08950_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__o211a_1
X_22632_ net2801 _07196_ net2780 VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_172_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25351_ net1525 _08906_ _08909_ _07247_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22563_ csr._minstret_T_3\[38\] _07147_ _07149_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24302_ _08064_ net2068 _08323_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__mux2_1
Xclkbuf_5_21__f_clock clknet_2_2_0_clock VGND VGND VPWR VPWR clknet_5_21__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_21514_ _06143_ net1940 _06274_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__mux2_1
X_28070_ clknet_leaf_216_clock _01092_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25282_ _08871_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1083 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22494_ _07088_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27021_ clknet_leaf_333_clock _00050_ VGND VGND VPWR VPWR decode.regfile.registers_22\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_24233_ _08291_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21445_ _06136_ net1444 _06230_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_359_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_359_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21376_ _06124_ net1718 _06199_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__mux2_1
X_24164_ _08057_ net1015 _08255_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23115_ _07098_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__clkbuf_8
X_20327_ _10864_ _10786_ decode.id_ex_pc_reg\[24\] _05482_ _10790_ VGND VGND VPWR
+ VPWR _05497_ sky130_fd_sc_hd__a41o_1
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28972_ clknet_leaf_109_clock _01985_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_24095_ net928 execute.io_target_pc\[3\] _06450_ VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__mux2_1
Xhold960 fetch.bht.bhtTable_target_pc\[8\]\[9\] VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold971 decode.regfile.registers_8\[15\] VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold982 decode.regfile.registers_21\[5\] VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__dlygate4sd3_1
X_23046_ fetch.bht.bhtTable_target_pc\[8\]\[9\] fetch.bht.bhtTable_target_pc\[9\]\[9\]
+ fetch.bht.bhtTable_target_pc\[10\]\[9\] fetch.bht.bhtTable_target_pc\[11\]\[9\]
+ _07407_ _07115_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__mux4_1
X_27923_ clknet_leaf_65_clock _00952_ VGND VGND VPWR VPWR csr.io_csr_write_enable
+ sky130_fd_sc_hd__dfxtp_1
X_20258_ _05444_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__clkbuf_1
Xhold993 decode.regfile.registers_25\[12\] VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27854_ clknet_leaf_325_clock _00883_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_129_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20189_ _05387_ _05388_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__xor2_1
XFILLER_0_215_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2350 decode.regfile.registers_17\[25\] VGND VGND VPWR VPWR net2577 sky130_fd_sc_hd__dlygate4sd3_1
X_26805_ net595 _09766_ _09773_ _09771_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__o211a_1
Xhold2361 decode.id_ex_rs1_data_reg\[5\] VGND VGND VPWR VPWR net2588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2372 decode.regfile.registers_4\[19\] VGND VGND VPWR VPWR net2599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27785_ clknet_leaf_334_clock _00814_ VGND VGND VPWR VPWR memory.io_wb_readdata\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_24997_ net1888 _08709_ _08711_ _06419_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__a211oi_1
Xhold2383 decode.regfile.registers_11\[14\] VGND VGND VPWR VPWR net2610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2394 decode.regfile.registers_10\[3\] VGND VGND VPWR VPWR net2621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1660 decode.regfile.registers_24\[15\] VGND VGND VPWR VPWR net1887 sky130_fd_sc_hd__dlygate4sd3_1
X_14750_ _10790_ _10791_ _10792_ VGND VGND VPWR VPWR _10793_ sky130_fd_sc_hd__or3_1
Xhold1671 csr._mcycle_T_3\[35\] VGND VGND VPWR VPWR net1898 sky130_fd_sc_hd__dlygate4sd3_1
X_26736_ _09412_ _09733_ VGND VGND VPWR VPWR _09734_ sky130_fd_sc_hd__nand2_1
X_29524_ clknet_leaf_265_clock _02537_ VGND VGND VPWR VPWR decode.regfile.registers_8\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_23948_ _08144_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__clkbuf_1
Xhold1682 csr.mcycle\[21\] VGND VGND VPWR VPWR net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1693 decode.regfile.registers_15\[23\] VGND VGND VPWR VPWR net1920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13701_ memory.csr_read_data_out_reg\[14\] _09989_ _10051_ VGND VGND VPWR VPWR _10052_
+ sky130_fd_sc_hd__o21bai_4
XFILLER_0_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29455_ clknet_leaf_261_clock _02468_ VGND VGND VPWR VPWR decode.regfile.registers_6\[21\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_196_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14681_ _10720_ execute.io_target_pc\[26\] _10722_ _10723_ VGND VGND VPWR VPWR _10724_
+ sky130_fd_sc_hd__o211a_1
X_26667_ _09422_ _09689_ VGND VGND VPWR VPWR _09694_ sky130_fd_sc_hd__nand2_1
X_23879_ execute.io_target_pc\[28\] VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__buf_2
X_16420_ _11371_ decode.regfile.registers_0\[29\] VGND VGND VPWR VPWR _12388_ sky130_fd_sc_hd__nand2_1
X_28406_ clknet_leaf_141_clock _01419_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_2
X_13632_ net957 _09989_ _09991_ VGND VGND VPWR VPWR _09992_ sky130_fd_sc_hd__o21ai_4
X_25618_ net847 _09068_ _09076_ _09074_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__o211a_1
X_29386_ clknet_leaf_259_clock _02399_ VGND VGND VPWR VPWR decode.regfile.registers_4\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26598_ _09428_ _09645_ VGND VGND VPWR VPWR _09654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28337_ clknet_leaf_237_clock _01350_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16351_ _12319_ _12065_ _12320_ VGND VGND VPWR VPWR _12321_ sky130_fd_sc_hd__a21oi_1
X_13563_ _09884_ _09914_ net289 net401 VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25549_ _08922_ _09036_ VGND VGND VPWR VPWR _09037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15302_ _11147_ VGND VGND VPWR VPWR _11298_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19070_ _04367_ _03704_ _04247_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__mux2_1
X_28268_ clknet_leaf_64_clock _01290_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16282_ decode.regfile.registers_11\[25\] _11180_ _12252_ _12253_ VGND VGND VPWR
+ VPWR _12254_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_229_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_217_Right_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18021_ _10609_ _12614_ _12629_ decode.regfile.registers_3\[31\] _03416_ VGND VGND
+ VPWR VPWR _03417_ sky130_fd_sc_hd__o221a_1
XFILLER_0_81_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15233_ decode.regfile.registers_21\[0\] _11061_ _11100_ _11224_ _11229_ VGND VGND
+ VPWR VPWR _11230_ sky130_fd_sc_hd__o311a_1
X_27219_ clknet_leaf_6_clock _00248_ VGND VGND VPWR VPWR decode.regfile.registers_29\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28199_ clknet_leaf_68_clock _01221_ VGND VGND VPWR VPWR csr.mscratch\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15164_ decode.regfile.registers_3\[0\] _11111_ _11142_ _11146_ _11160_ VGND VGND
+ VPWR VPWR _11161_ sky130_fd_sc_hd__a311o_1
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14115_ net2283 _10315_ _10324_ _10317_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19972_ net2741 _03599_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__nor2_1
X_15095_ _11091_ VGND VGND VPWR VPWR _11092_ sky130_fd_sc_hd__buf_4
X_14046_ _10147_ _10242_ VGND VGND VPWR VPWR _10284_ sky130_fd_sc_hd__nand2_1
X_18923_ _04220_ _04221_ _03790_ _03862_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18854_ _04149_ _04152_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17805_ decode.regfile.registers_15\[25\] _12585_ _12673_ VGND VGND VPWR VPWR _03207_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15997_ _10959_ decode.regfile.registers_26\[17\] _11349_ _10980_ _11347_ VGND VGND
+ VPWR VPWR _11977_ sky130_fd_sc_hd__o2111a_1
X_18785_ _03707_ decode.id_ex_imm_reg\[14\] VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17736_ _13407_ decode.regfile.registers_25\[23\] _13482_ _13294_ VGND VGND VPWR
+ VPWR _03140_ sky130_fd_sc_hd__or4_1
X_14948_ _10633_ VGND VGND VPWR VPWR _10976_ sky130_fd_sc_hd__clkbuf_4
X_14879_ _10912_ _10913_ _10916_ decode.immGen._imm_T_10\[2\] VGND VGND VPWR VPWR
+ _10919_ sky130_fd_sc_hd__and4bb_1
X_17667_ _12704_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__buf_2
XFILLER_0_202_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19406_ _04243_ _04433_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__or2_1
X_16618_ _12582_ VGND VGND VPWR VPWR _12583_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_214_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17598_ _03003_ _03004_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_214_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_1124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19337_ _04244_ _04273_ _04468_ _04628_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__a31o_1
X_16549_ _10595_ _11009_ _10925_ _12504_ VGND VGND VPWR VPWR _12514_ sky130_fd_sc_hd__or4_2
XFILLER_0_174_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19268_ _04050_ _04051_ _04516_ _04529_ _04400_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__o41ai_1
XFILLER_0_116_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18219_ csr.mcycle\[19\] VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__buf_2
XFILLER_0_54_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19199_ _03633_ decode.id_ex_aluop_reg\[3\] _03634_ _04299_ VGND VGND VPWR VPWR _04495_
+ sky130_fd_sc_hd__nor4_1
X_21230_ _06112_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold201 _10736_ VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 decode.regfile.registers_30\[14\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold223 decode.regfile.registers_30\[22\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold234 decode.id_ex_memtoreg_reg\[1\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
X_21161_ _06074_ _06070_ execute.csr_write_data_out_reg\[24\] VGND VGND VPWR VPWR
+ _06075_ sky130_fd_sc_hd__and3_1
Xhold245 decode.regfile.registers_14\[12\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold256 execute.csr_write_data_out_reg\[8\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold267 decode.regfile.registers_27\[3\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20112_ decode.id_ex_imm_reg\[13\] _10710_ _05310_ _05322_ VGND VGND VPWR VPWR _05323_
+ sky130_fd_sc_hd__o211ai_1
Xhold278 decode.regfile.registers_30\[0\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_TAPCELL_ROW_165_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21092_ _06034_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold289 decode.regfile.registers_18\[11\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20043_ _05249_ _05263_ _05255_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__nand3_1
X_24920_ net1087 _08659_ _08660_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_77_1203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24851_ _08613_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23802_ execute.io_target_pc\[3\] VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27570_ clknet_leaf_157_clock _00599_ VGND VGND VPWR VPWR csr.io_mem_pc\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_124_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24782_ _08577_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_124_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21994_ _06573_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_107 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_217_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26521_ _09426_ _09602_ VGND VGND VPWR VPWR _09610_ sky130_fd_sc_hd__nand2_1
X_23733_ net1402 csr.io_mem_pc\[29\] _08014_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__mux2_1
XANTENNA_118 _09128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_200_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_129 _10638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20945_ _05949_ _05945_ net58 VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29240_ clknet_leaf_170_clock _02253_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26452_ _09432_ _09558_ VGND VGND VPWR VPWR _09570_ sky130_fd_sc_hd__nand2_1
X_23664_ _07980_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_283_clock clknet_5_20__leaf_clock VGND VGND VPWR VPWR clknet_leaf_283_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20876_ _05916_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25403_ _10073_ VGND VGND VPWR VPWR _08945_ sky130_fd_sc_hd__clkbuf_8
X_29171_ clknet_leaf_188_clock _02184_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_22615_ net2156 _07185_ net2781 VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_27_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26383_ net2427 _09518_ _09529_ _09525_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_27_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23595_ _07943_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28122_ clknet_leaf_90_clock _01144_ VGND VGND VPWR VPWR csr.minstret\[27\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25334_ _08891_ net2622 VGND VGND VPWR VPWR _08898_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22546_ csr._minstret_T_3\[32\] _07136_ net2590 VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28053_ clknet_leaf_203_clock _01075_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_25265_ _08862_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_298_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_298_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22477_ _07071_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27004_ clknet_leaf_343_clock _00033_ VGND VGND VPWR VPWR decode.regfile.registers_22\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_24216_ _08282_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21428_ _06119_ net1595 _06219_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25196_ _10572_ net2669 _08826_ VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24147_ net850 execute.io_target_pc\[28\] _06427_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__mux2_1
X_21359_ _06107_ net2287 _06188_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_221_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_221_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_124_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24078_ _08211_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__clkbuf_1
X_28955_ clknet_leaf_172_clock _01968_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold790 fetch.bht.bhtTable_target_pc\[1\]\[29\] VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23029_ fetch.bht.bhtTable_target_pc\[12\]\[8\] fetch.bht.bhtTable_target_pc\[13\]\[8\]
+ fetch.bht.bhtTable_target_pc\[14\]\[8\] fetch.bht.bhtTable_target_pc\[15\]\[8\]
+ _07069_ _07111_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__mux4_1
X_27906_ clknet_leaf_18_clock _00935_ VGND VGND VPWR VPWR csr._mcycle_T_2\[27\] sky130_fd_sc_hd__dfxtp_2
X_15920_ decode.regfile.registers_20\[15\] _11452_ _11223_ _11901_ VGND VGND VPWR
+ VPWR _11902_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_53_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28886_ clknet_leaf_124_clock _01899_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15851_ _11252_ VGND VGND VPWR VPWR _11834_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_236_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_236_clock
+ sky130_fd_sc_hd__clkbuf_8
X_27837_ clknet_leaf_326_clock _00866_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2180 decode.regfile.registers_24\[28\] VGND VGND VPWR VPWR net2407 sky130_fd_sc_hd__dlygate4sd3_1
X_14802_ decode.id_ex_pc_reg\[15\] _10764_ _10809_ _10811_ _10844_ VGND VGND VPWR
+ VPWR _10845_ sky130_fd_sc_hd__o311a_1
Xhold2191 decode.regfile.registers_11\[17\] VGND VGND VPWR VPWR net2418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15782_ decode.regfile.registers_1\[12\] _11539_ _11766_ VGND VGND VPWR VPWR _11767_
+ sky130_fd_sc_hd__a21o_1
X_18570_ execute.csr_read_data_out_reg\[23\] _03661_ _03660_ VGND VGND VPWR VPWR _03869_
+ sky130_fd_sc_hd__or3_1
X_27768_ clknet_leaf_321_clock _00797_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1490 decode.regfile.registers_17\[21\] VGND VGND VPWR VPWR net1717 sky130_fd_sc_hd__dlygate4sd3_1
X_14733_ _10771_ _10775_ csr.io_mem_pc\[29\] VGND VGND VPWR VPWR _10776_ sky130_fd_sc_hd__a21oi_1
X_17521_ _11020_ _12490_ _12512_ decode.regfile.registers_12\[18\] _12591_ VGND VGND
+ VPWR VPWR _13468_ sky130_fd_sc_hd__o32a_1
X_29507_ clknet_leaf_252_clock _02520_ VGND VGND VPWR VPWR decode.regfile.registers_8\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_26719_ net537 _09723_ _09724_ _09717_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27699_ clknet_leaf_22_clock _00728_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17452_ decode.regfile.registers_19\[16\] _12679_ _12906_ _13400_ VGND VGND VPWR
+ VPWR _13401_ sky130_fd_sc_hd__o211a_1
X_14664_ _10706_ VGND VGND VPWR VPWR _10707_ sky130_fd_sc_hd__inv_2
X_29438_ clknet_leaf_248_clock _02451_ VGND VGND VPWR VPWR decode.regfile.registers_6\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16403_ decode.regfile.registers_22\[28\] _11096_ _12370_ _12371_ VGND VGND VPWR
+ VPWR _12372_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13615_ net670 _09938_ _09976_ _09957_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__o211a_1
X_17383_ _12494_ decode.regfile.registers_26\[14\] _13002_ _11010_ _11026_ VGND VGND
+ VPWR VPWR _13334_ sky130_fd_sc_hd__o2111a_1
X_29369_ clknet_leaf_246_clock _02382_ VGND VGND VPWR VPWR decode.regfile.registers_3\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14595_ _10637_ VGND VGND VPWR VPWR _10638_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19122_ _04280_ _04282_ _04324_ _04276_ _04418_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__o221a_1
X_16334_ _11260_ _12302_ _12303_ _12304_ VGND VGND VPWR VPWR _12305_ sky130_fd_sc_hd__a31o_1
X_13546_ _09879_ _09882_ VGND VGND VPWR VPWR _09917_ sky130_fd_sc_hd__nor2_4
XFILLER_0_82_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19053_ _03872_ _03844_ _03989_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__mux2_1
X_16265_ _11942_ net2782 _12095_ _12096_ _12097_ VGND VGND VPWR VPWR _12237_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_11_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18004_ _12712_ decode.regfile.registers_24\[30\] _12997_ _12998_ _11025_ VGND VGND
+ VPWR VPWR _03401_ sky130_fd_sc_hd__o2111a_1
X_15216_ decode.regfile.registers_18\[0\] _10955_ _11114_ _10989_ _10977_ VGND VGND
+ VPWR VPWR _11213_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_51_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16196_ _10959_ decode.regfile.registers_26\[23\] _11349_ _11348_ _10993_ VGND VGND
+ VPWR VPWR _12170_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_51_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15147_ _11091_ _11041_ _11143_ VGND VGND VPWR VPWR _11144_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19955_ net596 _03599_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__nor2_1
X_15078_ _11074_ VGND VGND VPWR VPWR _11075_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_207_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14029_ net2456 _10271_ _10274_ _10275_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__o211a_1
X_18906_ _03900_ _03914_ _03908_ decode.id_ex_rs1_data_reg\[19\] _03901_ VGND VGND
+ VPWR VPWR _04205_ sky130_fd_sc_hd__o221a_2
X_19886_ _04386_ _04776_ _05141_ _05155_ _04515_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_203_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18837_ _03816_ _04135_ net353 VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_117_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18768_ execute.io_reg_pc\[6\] _03776_ _03664_ net128 _04066_ VGND VGND VPWR VPWR
+ _04067_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17719_ decode.regfile.registers_6\[23\] _12735_ _12623_ _03122_ VGND VGND VPWR VPWR
+ _03123_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_136_1167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18699_ decode.id_ex_immsrc_reg decode.id_ex_imm_reg\[1\] VGND VGND VPWR VPWR _03998_
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_203_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20730_ _05804_ _00709_ _05834_ _05835_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__a31o_1
XFILLER_0_212_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20661_ csr.minstret\[31\] _05560_ _05622_ csr._csr_read_data_T_8\[31\] _05789_ VGND
+ VGND VPWR VPWR _05790_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22400_ fetch.bht.bhtTable_tag\[14\]\[21\] fetch.bht.bhtTable_tag\[15\]\[21\] _06616_
+ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23380_ _06795_ _07706_ _07707_ _07804_ _07705_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__o311a_2
X_20592_ csr._minstret_T_3\[53\] _05616_ _05618_ csr._csr_read_data_T_8\[21\] _05730_
+ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__a221o_1
X_22331_ _06925_ _06687_ _06640_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25050_ net1909 _08645_ _08746_ _06419_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_6_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22262_ _06730_ _06856_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24001_ net954 execute.io_target_pc\[21\] _08164_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21213_ _10820_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__buf_2
X_22193_ _06786_ _06787_ _06632_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21144_ _06065_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28740_ clknet_leaf_131_clock _01753_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25952_ _08948_ _09267_ VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__nand2_1
X_21075_ execute.csr_read_data_out_reg\[26\] _06014_ _03583_ VGND VGND VPWR VPWR _06024_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_126_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20026_ decode.id_ex_imm_reg\[4\] decode.id_ex_pc_reg\[4\] VGND VGND VPWR VPWR _05249_
+ sky130_fd_sc_hd__nand2_1
X_24903_ csr._mcycle_T_3\[35\] _08649_ _07179_ VGND VGND VPWR VPWR _08650_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_214_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28671_ clknet_leaf_176_clock _01684_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_25883_ _08956_ _09223_ VGND VGND VPWR VPWR _09229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_225_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27622_ clknet_leaf_147_clock _00651_ VGND VGND VPWR VPWR execute.io_target_pc\[31\]
+ sky130_fd_sc_hd__dfxtp_4
X_24834_ _08604_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27553_ clknet_leaf_42_clock _00582_ VGND VGND VPWR VPWR execute.io_mem_memtoreg\[1\]
+ sky130_fd_sc_hd__dfxtp_4
X_24765_ _08568_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__clkbuf_1
X_21977_ _06578_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer60 _09928_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer71 net302 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_1
X_26504_ _09408_ _09589_ VGND VGND VPWR VPWR _09600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23716_ net1349 csr.io_mem_pc\[21\] _08003_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__mux2_1
Xrebuffer82 _04038_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_166_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27484_ clknet_leaf_38_clock _00513_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dfxtp_2
X_20928_ _05944_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__clkbuf_1
X_24696_ _08057_ net1647 _08531_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__mux2_1
Xrebuffer93 net319 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29223_ clknet_leaf_106_clock _02236_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_26435_ _09415_ _09558_ VGND VGND VPWR VPWR _09560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23647_ _07971_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20859_ net116 _05903_ _05899_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29154_ clknet_leaf_165_clock _02167_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26366_ net2377 _09518_ _09520_ _09512_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__o211a_1
X_14380_ net722 _10477_ _10478_ _10468_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23578_ _06109_ net2119 _07930_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28105_ clknet_leaf_75_clock net607 VGND VGND VPWR VPWR csr.minstret\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_92_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25317_ _08880_ net2737 VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22529_ _07068_ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_187_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29085_ clknet_leaf_71_clock _02098_ VGND VGND VPWR VPWR csr._mcycle_T_3\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26297_ decode.regfile.registers_12\[24\] _09475_ _09480_ _09471_ VGND VGND VPWR
+ VPWR _02663_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28036_ clknet_leaf_188_clock _01058_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16050_ _11291_ _12026_ _12027_ VGND VGND VPWR VPWR _12028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_228_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25248_ _08087_ net2226 _08848_ VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_160_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_160_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15001_ _11012_ _11004_ _11006_ _11007_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25179_ net407 _08818_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_55_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19740_ _05014_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__inv_2
X_28938_ clknet_leaf_98_clock _01951_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16952_ _10927_ decode.regfile.registers_24\[4\] _10933_ _12759_ _12862_ VGND VGND
+ VPWR VPWR _12913_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_60_1070 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_175_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_175_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_217_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15903_ _11043_ decode.regfile.registers_4\[15\] _11503_ _10629_ _11462_ VGND VGND
+ VPWR VPWR _11885_ sky130_fd_sc_hd__a2111o_1
X_19671_ _04735_ _04245_ _04428_ _04949_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__a31o_1
XFILLER_0_216_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28869_ clknet_leaf_136_clock _01882_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16883_ _12841_ _12844_ VGND VGND VPWR VPWR _12845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_218_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18622_ _03785_ _10073_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__nand2_1
X_15834_ decode.regfile.registers_16\[13\] _11123_ _11799_ _11817_ VGND VGND VPWR
+ VPWR _11818_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_204_Left_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18553_ _03835_ _03838_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_194_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ decode.regfile.registers_23\[11\] _11232_ _11074_ _11750_ VGND VGND VPWR
+ VPWR _11751_ sky130_fd_sc_hd__a211o_1
XFILLER_0_220_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17504_ _10930_ VGND VGND VPWR VPWR _13451_ sky130_fd_sc_hd__clkbuf_4
X_14716_ csr.io_mem_pc\[27\] VGND VGND VPWR VPWR _10759_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_190_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15696_ _11646_ _11253_ _11064_ decode.regfile.registers_29\[9\] _11683_ VGND VGND
+ VPWR VPWR _11684_ sky130_fd_sc_hd__o221a_1
X_18484_ _03673_ _03740_ _03761_ _03742_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_190_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14647_ decode.id_ex_pc_reg\[4\] VGND VGND VPWR VPWR _10690_ sky130_fd_sc_hd__inv_2
X_17435_ _13382_ _12932_ _10615_ _12933_ _13383_ VGND VGND VPWR VPWR _13384_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_113_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_113_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _05059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_29 _08939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ _10612_ _10613_ decode.id_ex_ex_rd_reg\[4\] _10595_ _10620_ VGND VGND VPWR
+ VPWR _10621_ sky130_fd_sc_hd__a221o_1
X_17366_ _13311_ _13316_ _12735_ decode.regfile.registers_6\[14\] VGND VGND VPWR VPWR
+ _13317_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_126_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19105_ net314 _04320_ net317 _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__a31oi_1
X_13529_ _09905_ VGND VGND VPWR VPWR _09906_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_172_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16317_ decode.regfile.registers_8\[26\] _11285_ _11382_ _12287_ VGND VGND VPWR VPWR
+ _12288_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17297_ _10926_ VGND VGND VPWR VPWR _13250_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_213_Left_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16248_ decode.regfile.registers_13\[24\] _11047_ _11690_ _11198_ _12220_ VGND VGND
+ VPWR VPWR _12221_ sky130_fd_sc_hd__o311a_1
XFILLER_0_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19036_ _04160_ _04334_ _03989_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_209_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_128_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_128_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_209_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput103 net103 VGND VGND VPWR VPWR io_memory_address[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16179_ decode.regfile.registers_15\[22\] _11036_ _11205_ VGND VGND VPWR VPWR _12154_
+ sky130_fd_sc_hd__and3_1
Xoutput114 net114 VGND VGND VPWR VPWR io_memory_address[22] sky130_fd_sc_hd__clkbuf_4
Xoutput125 net125 VGND VGND VPWR VPWR io_memory_address[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput136 net136 VGND VGND VPWR VPWR io_memory_write_data[0] sky130_fd_sc_hd__clkbuf_4
Xoutput147 net147 VGND VGND VPWR VPWR io_memory_write_data[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput158 net158 VGND VGND VPWR VPWR io_memory_write_data[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19938_ _03581_ _05201_ net461 VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__and3b_1
XFILLER_0_103_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_9 _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_222_Left_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19869_ _04251_ _04252_ _05137_ _04304_ _05138_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__a311o_1
XFILLER_0_208_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21900_ csr.io_mret_vector\[19\] _10800_ _06539_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__mux2_1
X_22880_ net1453 _10760_ _07335_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21831_ _06479_ net590 _06396_ _06490_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24550_ _08456_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_156_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21762_ net1036 _10795_ _06439_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23501_ net1153 _07890_ _07887_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__or3b_1
XFILLER_0_93_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20713_ _05801_ _05808_ decode.id_ex_rs1_data_reg\[15\] _05825_ _00702_ VGND VGND
+ VPWR VPWR _00734_ sky130_fd_sc_hd__a32o_1
X_24481_ _08420_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__clkbuf_1
X_21693_ _03449_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__buf_6
XFILLER_0_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26220_ net2667 _09419_ _09433_ _09418_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23432_ _04459_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20644_ _05540_ csr.io_mret_vector\[29\] _05565_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_119_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26151_ _09998_ VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__buf_4
X_23363_ net86 _07706_ _07707_ _07788_ _07705_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__o311a_1
XFILLER_0_116_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20575_ _05439_ _05716_ _03449_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_115_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25102_ _08779_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22314_ fetch.bht.bhtTable_tag\[10\]\[0\] fetch.bht.bhtTable_tag\[11\]\[0\] _06644_
+ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26082_ _08929_ _09340_ VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__nand2_1
X_23294_ fetch.bht.bhtTable_target_pc\[12\]\[23\] fetch.bht.bhtTable_target_pc\[13\]\[23\]
+ fetch.bht.bhtTable_target_pc\[14\]\[23\] fetch.bht.bhtTable_target_pc\[15\]\[23\]
+ _07708_ _07710_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25033_ _10019_ _08734_ _08735_ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29910_ clknet_leaf_340_clock _02923_ VGND VGND VPWR VPWR decode.regfile.registers_20\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_22245_ fetch.bht.bhtTable_tag\[4\]\[19\] fetch.bht.bhtTable_tag\[5\]\[19\] _06706_
+ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_1092 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_92_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_92_clock
+ sky130_fd_sc_hd__clkbuf_8
X_29841_ clknet_leaf_299_clock _02854_ VGND VGND VPWR VPWR decode.regfile.registers_18\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_22176_ fetch.bht.bhtTable_tag\[4\]\[25\] fetch.bht.bhtTable_tag\[5\]\[25\] _06646_
+ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21127_ _06050_ _06046_ net1561 VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__and3_1
X_29772_ clknet_leaf_295_clock _02785_ VGND VGND VPWR VPWR decode.regfile.registers_16\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26984_ net2241 _09866_ _09875_ _09865_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_50_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28723_ clknet_leaf_140_clock _01736_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21058_ _06015_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__clkbuf_1
X_25935_ _08933_ _09253_ VGND VGND VPWR VPWR _09259_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_145_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20009_ decode.id_ex_imm_reg\[0\] decode.id_ex_pc_reg\[0\] decode.id_ex_pc_reg\[1\]
+ decode.id_ex_imm_reg\[1\] VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__a22o_1
X_28654_ clknet_leaf_112_clock _01667_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_13880_ _10117_ _10177_ VGND VGND VPWR VPWR _10187_ sky130_fd_sc_hd__nand2_1
X_25866_ _08939_ _09210_ VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24817_ _08595_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27605_ clknet_leaf_158_clock _00634_ VGND VGND VPWR VPWR execute.io_target_pc\[14\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_193_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28585_ clknet_leaf_101_clock _01598_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25797_ _09155_ VGND VGND VPWR VPWR _09179_ sky130_fd_sc_hd__buf_2
XFILLER_0_198_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15550_ decode.regfile.registers_0\[6\] _11539_ _11540_ VGND VGND VPWR VPWR _11541_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24748_ _08558_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__clkbuf_1
X_27536_ clknet_leaf_155_clock _00565_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_48_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_208 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clock clknet_5_3__leaf_clock VGND VGND VPWR VPWR clknet_leaf_30_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_219 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14501_ _10147_ _10505_ VGND VGND VPWR VPWR _10547_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _11472_ _11473_ VGND VGND VPWR VPWR _11474_ sky130_fd_sc_hd__and2_1
X_27467_ clknet_leaf_27_clock _00496_ VGND VGND VPWR VPWR csr.io_csr_address\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_96_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24679_ net1977 execute.io_target_pc\[28\] _07285_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29206_ clknet_leaf_240_clock _02219_ VGND VGND VPWR VPWR fetch.btb.btbTable\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17220_ _12695_ _13172_ _13173_ _13174_ VGND VGND VPWR VPWR _13175_ sky130_fd_sc_hd__a31o_1
X_14432_ _10426_ VGND VGND VPWR VPWR _10509_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_182_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26418_ net901 _09548_ _09550_ _09540_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__o211a_1
X_27398_ clknet_leaf_27_clock _00427_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_182_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17151_ _13105_ _12732_ _13106_ VGND VGND VPWR VPWR _13107_ sky130_fd_sc_hd__a21o_1
X_29137_ clknet_leaf_79_clock _02150_ VGND VGND VPWR VPWR csr.mcycle\[21\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_45_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_45_clock
+ sky130_fd_sc_hd__clkbuf_8
X_26349_ net2396 _09505_ _09510_ _09499_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14363_ _09975_ _10464_ VGND VGND VPWR VPWR _10469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput16 io_fetch_data[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xinput27 net373 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
X_16102_ _12078_ decode.regfile.registers_17\[20\] _11357_ VGND VGND VPWR VPWR _12079_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 io_memory_read_data[13] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
X_29068_ clknet_leaf_196_clock _02081_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput49 io_memory_read_data[23] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
X_17082_ decode.regfile.registers_22\[7\] _12527_ _13038_ _13039_ _12686_ VGND VGND
+ VPWR VPWR _13040_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14294_ _09999_ _10420_ VGND VGND VPWR VPWR _10429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16033_ _11251_ _11259_ decode.regfile.registers_27\[18\] _11984_ _12011_ VGND VGND
+ VPWR VPWR _12012_ sky130_fd_sc_hd__o32a_1
XFILLER_0_165_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28019_ clknet_leaf_239_clock _01041_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17984_ decode.regfile.registers_2\[30\] _12834_ _12639_ decode.regfile.registers_3\[30\]
+ _12837_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_100_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_200_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19723_ _03888_ _03893_ _04998_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_196_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16935_ decode.regfile.registers_12\[4\] _12591_ _12877_ _12895_ VGND VGND VPWR VPWR
+ _12896_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_196_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_221_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19654_ _04932_ _04192_ _04526_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__a21oi_1
X_16866_ decode.regfile.registers_13\[3\] _12533_ _12587_ _12662_ VGND VGND VPWR VPWR
+ _12828_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_192_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18605_ _03658_ execute.csr_read_data_out_reg\[17\] execute.io_reg_pc\[17\] _03776_
+ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__o22a_1
X_15817_ decode.regfile.registers_7\[13\] _11308_ _11169_ decode.regfile.registers_6\[13\]
+ _11165_ VGND VGND VPWR VPWR _11801_ sky130_fd_sc_hd__a221o_1
X_19585_ _04211_ _04197_ _04198_ _04866_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__or4_4
X_16797_ _12758_ _12760_ VGND VGND VPWR VPWR _12761_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18536_ decode.id_ex_rs1_data_reg\[25\] _03817_ _03698_ _03834_ VGND VGND VPWR VPWR
+ _03835_ sky130_fd_sc_hd__o31a_4
X_15748_ _11043_ decode.regfile.registers_4\[11\] _11503_ _10629_ _11083_ VGND VGND
+ VPWR VPWR _11734_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18467_ _03709_ decode.id_ex_imm_reg\[31\] _03729_ _03765_ VGND VGND VPWR VPWR _03766_
+ sky130_fd_sc_hd__a22oi_4
X_15679_ decode.regfile.registers_17\[9\] _10652_ _11112_ _11118_ _11666_ VGND VGND
+ VPWR VPWR _11667_ sky130_fd_sc_hd__a41o_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17418_ _13250_ decode.regfile.registers_24\[15\] _13170_ _13083_ _13367_ VGND VGND
+ VPWR VPWR _13368_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_151_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18398_ _03696_ _03678_ _03673_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__nand3_1
XFILLER_0_56_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17349_ _13099_ _13262_ _13182_ decode.regfile.registers_29\[13\] _13300_ VGND VGND
+ VPWR VPWR _13301_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20360_ csr.io_csr_address\[4\] csr.io_csr_address\[5\] csr.io_csr_address\[7\] csr.io_csr_address\[6\]
+ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__nor4_2
XFILLER_0_114_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19019_ decode.id_ex_imm_reg\[0\] _03728_ _03999_ _04002_ _04309_ VGND VGND VPWR
+ VPWR _04318_ sky130_fd_sc_hd__o221a_2
XFILLER_0_140_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20291_ _05417_ _05326_ _05469_ _05454_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_228_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_228_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22030_ fetch.bht.bhtTable_tag\[8\]\[22\] fetch.bht.bhtTable_tag\[9\]\[22\] fetch.bht.bhtTable_tag\[10\]\[22\]
+ fetch.bht.bhtTable_tag\[11\]\[22\] _06619_ _06624_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_149_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23981_ _08161_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25720_ _08943_ _09122_ VGND VGND VPWR VPWR _09135_ sky130_fd_sc_hd__nand2_1
X_22932_ execute.io_target_pc\[2\] _07346_ _07348_ _07382_ VGND VGND VPWR VPWR _07383_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_108_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25651_ _09067_ VGND VGND VPWR VPWR _09095_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_190_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22863_ net1760 csr.io_mem_pc\[18\] _07324_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24602_ _08483_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_179_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_119_Left_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28370_ clknet_leaf_209_clock _01383_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21814_ _06478_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25582_ net2196 _09052_ _09055_ _09046_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__o211a_1
X_22794_ net1127 _10812_ _07286_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27321_ clknet_leaf_31_clock _00350_ VGND VGND VPWR VPWR decode.id_ex_ex_rs1_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_24533_ _08093_ net2082 _08439_ VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__mux2_1
X_21745_ net903 csr.io_mem_pc\[12\] _06428_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27252_ clknet_leaf_31_clock _00281_ VGND VGND VPWR VPWR decode.regfile.registers_30\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_24464_ _08091_ net1644 _08411_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21676_ net2535 _06383_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26203_ _10091_ VGND VGND VPWR VPWR _09422_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23415_ _07070_ _07836_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20627_ csr._minstret_T_3\[58\] _05616_ _05618_ csr._csr_read_data_T_8\[26\] _05760_
+ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27183_ clknet_leaf_352_clock _00212_ VGND VGND VPWR VPWR decode.regfile.registers_28\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_24395_ net753 execute.io_target_pc\[20\] _08367_ VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26134_ _09372_ VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__clkbuf_4
X_23346_ _07089_ _07768_ _07769_ _07772_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20558_ csr._minstret_T_3\[48\] _05577_ _05578_ _05701_ VGND VGND VPWR VPWR _05702_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_225_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_128_Left_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26065_ net2065 _09329_ _09334_ _09333_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__o211a_1
X_23277_ _07098_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__buf_4
XFILLER_0_105_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20489_ csr.mtip _05604_ _05640_ _05641_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25016_ csr._mcycle_T_2\[10\] _08712_ _08722_ csr.mcycle\[9\] csr.mcycle\[10\] VGND
+ VGND VPWR VPWR _08724_ sky130_fd_sc_hd__a221oi_1
X_22228_ fetch.bht.bhtTable_tag\[0\]\[15\] fetch.bht.bhtTable_tag\[1\]\[15\] fetch.bht.bhtTable_tag\[2\]\[15\]
+ fetch.bht.bhtTable_tag\[3\]\[15\] _06617_ _06622_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__mux4_1
X_29824_ clknet_leaf_307_clock _02837_ VGND VGND VPWR VPWR decode.regfile.registers_18\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22159_ _06616_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29755_ clknet_leaf_310_clock _02768_ VGND VGND VPWR VPWR decode.regfile.registers_16\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_14981_ _10948_ _10954_ _10997_ net1121 _10999_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__o311a_1
X_26967_ net198 _09862_ VGND VGND VPWR VPWR _09867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28706_ clknet_leaf_135_clock _01719_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16720_ _12525_ _11009_ _10925_ _12523_ VGND VGND VPWR VPWR _12685_ sky130_fd_sc_hd__and4_1
X_13932_ _10131_ VGND VGND VPWR VPWR _10219_ sky130_fd_sc_hd__clkbuf_4
X_25918_ _08916_ _09243_ VGND VGND VPWR VPWR _09249_ sky130_fd_sc_hd__nand2_1
X_29686_ clknet_leaf_282_clock _02699_ VGND VGND VPWR VPWR decode.regfile.registers_13\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_26898_ _09426_ _09819_ VGND VGND VPWR VPWR _09827_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_137_Left_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28637_ clknet_leaf_177_clock _01650_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16651_ _10591_ VGND VGND VPWR VPWR _12616_ sky130_fd_sc_hd__clkbuf_4
X_13863_ _10074_ _10177_ VGND VGND VPWR VPWR _10178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25849_ net1337 _09199_ _09208_ _09209_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15602_ decode.regfile.registers_13\[7\] _10639_ _11187_ _11590_ _11591_ VGND VGND
+ VPWR VPWR _11592_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19370_ _04144_ _04645_ _04454_ _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__o211ai_1
X_28568_ clknet_leaf_199_clock _01581_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_13794_ _10130_ VGND VGND VPWR VPWR _10131_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16582_ _10607_ _10614_ VGND VGND VPWR VPWR _12547_ sky130_fd_sc_hd__nor2_1
X_18321_ decode.id_ex_rs2_data_reg\[26\] _03616_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27519_ clknet_leaf_47_clock _00548_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_4
X_15533_ _10960_ decode.regfile.registers_28\[5\] _11067_ _11038_ _11440_ VGND VGND
+ VPWR VPWR _11525_ sky130_fd_sc_hd__o2111a_1
X_28499_ clknet_leaf_184_clock _01512_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15464_ decode.regfile.registers_14\[4\] _11360_ _11273_ decode.regfile.registers_15\[4\]
+ _11361_ VGND VGND VPWR VPWR _11457_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18252_ decode.id_ex_funct3_reg\[1\] VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17203_ _12650_ _12772_ _12669_ decode.regfile.registers_14\[10\] _13157_ VGND VGND
+ VPWR VPWR _13158_ sky130_fd_sc_hd__o221a_1
X_14415_ _10117_ _10487_ VGND VGND VPWR VPWR _10498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18183_ decode.control.io_funct3\[2\] _10943_ decode.control.io_funct3\[0\] VGND
+ VGND VPWR VPWR _03521_ sky130_fd_sc_hd__nor3_1
X_15395_ decode.regfile.registers_19\[2\] _11354_ _11218_ _11389_ VGND VGND VPWR VPWR
+ _11390_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_146_Left_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_1228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17134_ _10939_ VGND VGND VPWR VPWR _13091_ sky130_fd_sc_hd__buf_2
X_14346_ _10136_ _10418_ VGND VGND VPWR VPWR _10458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold608 fetch.bht.bhtTable_tag\[8\]\[9\] VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17065_ decode.regfile.registers_8\[7\] _12892_ _12603_ _13022_ VGND VGND VPWR VPWR
+ _13023_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_204_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold619 fetch.bht.bhtTable_tag\[6\]\[8\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ _10417_ VGND VGND VPWR VPWR _10418_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16016_ _11993_ _11994_ VGND VGND VPWR VPWR _11995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_228_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_223_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_223_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2009 decode.io_id_pc\[21\] VGND VGND VPWR VPWR net2236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_1340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_209_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1308 fetch.bht.bhtTable_tag\[0\]\[5\] VGND VGND VPWR VPWR net1535 sky130_fd_sc_hd__dlygate4sd3_1
X_17967_ _12712_ decode.regfile.registers_24\[29\] _12997_ _12690_ _11025_ VGND VGND
+ VPWR VPWR _03365_ sky130_fd_sc_hd__o2111a_1
Xhold1319 fetch.bht.bhtTable_target_pc\[6\]\[23\] VGND VGND VPWR VPWR net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_155_Left_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19706_ _03888_ _04234_ _04277_ _04265_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__o211a_1
X_16918_ _10602_ _12508_ _12613_ VGND VGND VPWR VPWR _12879_ sky130_fd_sc_hd__or3_1
XFILLER_0_174_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17898_ _10929_ decode.regfile.registers_28\[27\] _02992_ VGND VGND VPWR VPWR _03298_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19637_ _04910_ _04916_ _04908_ _04667_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__o2bb2a_1
X_16849_ _12811_ VGND VGND VPWR VPWR _12812_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_177_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19568_ _04281_ _04283_ _04849_ _04850_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__o31a_1
XFILLER_0_215_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_215_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18519_ _03659_ execute.csr_read_data_out_reg\[27\] execute.io_reg_pc\[27\] _03777_
+ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19499_ _04186_ _04782_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_174_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21530_ _06101_ net1550 _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_164_Left_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21461_ _06246_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_170_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23200_ _06887_ _07613_ net76 VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20412_ csr.io_csr_address\[11\] _05526_ net218 _05520_ VGND VGND VPWR VPWR _05571_
+ sky130_fd_sc_hd__and4_1
X_24180_ _08074_ net1676 _08255_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__mux2_1
X_21392_ _06140_ net2044 _06199_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23131_ csr._csr_read_data_T_8\[13\] _06039_ csr.io_mret_vector\[13\] _06463_ _07570_
+ VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__a221o_1
X_20343_ _10854_ decode.id_ex_pc_reg\[28\] _05500_ _10697_ VGND VGND VPWR VPWR _05509_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_222_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23062_ _07391_ _07392_ _07503_ _07504_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_141_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20274_ _05455_ _05456_ _05411_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__a21oi_1
X_22013_ net2158 _06600_ _06611_ _06605_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27870_ clknet_leaf_326_clock _00899_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2510 decode.regfile.registers_0\[20\] VGND VGND VPWR VPWR net2737 sky130_fd_sc_hd__dlygate4sd3_1
X_26821_ net1748 _09779_ _09782_ _09771_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_4_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2521 execute.csr_write_data_out_reg\[22\] VGND VGND VPWR VPWR net2748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2532 decode.regfile.registers_4\[14\] VGND VGND VPWR VPWR net2759 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2543 csr._mcycle_T_2\[13\] VGND VGND VPWR VPWR net2770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2554 csr._minstret_T_3\[53\] VGND VGND VPWR VPWR net2781 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1820 fetch.bht.bhtTable_tag\[13\]\[8\] VGND VGND VPWR VPWR net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2565 net90 VGND VGND VPWR VPWR net2792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1831 fetch.bht.bhtTable_tag\[15\]\[10\] VGND VGND VPWR VPWR net2058 sky130_fd_sc_hd__dlygate4sd3_1
X_29540_ clknet_leaf_267_clock _02553_ VGND VGND VPWR VPWR decode.regfile.registers_9\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_23964_ _08152_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__clkbuf_1
Xhold2576 csr._mcycle_T_2\[31\] VGND VGND VPWR VPWR net2803 sky130_fd_sc_hd__dlygate4sd3_1
X_26752_ _09701_ VGND VGND VPWR VPWR _09743_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_32_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1842 decode.regfile.registers_26\[17\] VGND VGND VPWR VPWR net2069 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1853 decode.regfile.registers_8\[13\] VGND VGND VPWR VPWR net2080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1864 decode.regfile.registers_5\[30\] VGND VGND VPWR VPWR net2091 sky130_fd_sc_hd__dlygate4sd3_1
X_22915_ _06768_ _07359_ _07365_ _06896_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__and4_2
Xhold1875 fetch.bht.bhtTable_tag\[14\]\[5\] VGND VGND VPWR VPWR net2102 sky130_fd_sc_hd__dlygate4sd3_1
X_25703_ _09110_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__buf_2
Xhold1886 fetch.bht.bhtTable_tag\[7\]\[18\] VGND VGND VPWR VPWR net2113 sky130_fd_sc_hd__dlygate4sd3_1
X_26683_ _09436_ _09664_ VGND VGND VPWR VPWR _09703_ sky130_fd_sc_hd__nand2_1
X_29471_ clknet_leaf_250_clock _02484_ VGND VGND VPWR VPWR decode.regfile.registers_7\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_23895_ net1122 _08053_ _06179_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1897 fetch.bht.bhtTable_target_pc\[13\]\[2\] VGND VGND VPWR VPWR net2124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28422_ clknet_leaf_39_clock _01435_ VGND VGND VPWR VPWR decode.control.io_funct3\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_211_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22846_ net1413 _10878_ _09898_ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25634_ net1933 _09082_ _09085_ _09074_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28353_ clknet_leaf_186_clock _01366_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_25565_ _08990_ VGND VGND VPWR VPWR _09046_ sky130_fd_sc_hd__buf_2
X_22777_ _06151_ net2198 _07276_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24516_ _09901_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27304_ clknet_leaf_13_clock _00333_ VGND VGND VPWR VPWR decode.regfile.registers_31\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_21728_ _06422_ _09923_ _06025_ _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_82_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28284_ clknet_leaf_85_clock _01306_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_25496_ _08945_ _09005_ VGND VGND VPWR VPWR _09006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24447_ _08074_ net1601 _08400_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__mux2_1
X_27235_ clknet_leaf_364_clock _00264_ VGND VGND VPWR VPWR decode.regfile.registers_29\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21659_ csr._mcycle_T_2\[17\] _06325_ _06370_ csr.minstret\[17\] VGND VGND VPWR VPWR
+ _06371_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_62_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14200_ net331 VGND VGND VPWR VPWR _10373_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27166_ clknet_leaf_359_clock _00195_ VGND VGND VPWR VPWR decode.regfile.registers_27\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15180_ decode.regfile.registers_9\[0\] _10639_ _11134_ _11172_ _11176_ VGND VGND
+ VPWR VPWR _11177_ sky130_fd_sc_hd__a32o_1
X_24378_ net1339 execute.io_target_pc\[12\] _08356_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14131_ _09964_ _10333_ VGND VGND VPWR VPWR _10335_ sky130_fd_sc_hd__nand2_1
X_26117_ net2734 _09356_ _09363_ _09359_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23329_ _07075_ _07752_ _07754_ _07756_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27097_ clknet_leaf_357_clock _00126_ VGND VGND VPWR VPWR decode.regfile.registers_25\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14062_ _09984_ _10288_ VGND VGND VPWR VPWR _10295_ sky130_fd_sc_hd__nand2_1
X_26048_ net2655 _09313_ _09323_ _09318_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18870_ _04132_ _04144_ _04155_ _04168_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__nand4_1
XFILLER_0_98_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17821_ _12967_ _03220_ _03221_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__a31o_1
X_29807_ clknet_leaf_296_clock _02820_ VGND VGND VPWR VPWR decode.regfile.registers_17\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27999_ clknet_leaf_203_clock _01021_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17752_ decode.regfile.registers_0\[24\] _12932_ _12834_ _03154_ VGND VGND VPWR VPWR
+ _03155_ sky130_fd_sc_hd__a211o_1
X_29738_ clknet_leaf_285_clock _02751_ VGND VGND VPWR VPWR decode.regfile.registers_15\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_14964_ _10988_ VGND VGND VPWR VPWR _10989_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16703_ _11018_ _10617_ _12488_ _10603_ VGND VGND VPWR VPWR _12668_ sky130_fd_sc_hd__or4_1
X_13915_ _10008_ _10200_ VGND VGND VPWR VPWR _10209_ sky130_fd_sc_hd__nand2_1
X_29669_ clknet_leaf_281_clock _02682_ VGND VGND VPWR VPWR decode.regfile.registers_13\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_17683_ decode.regfile.registers_10\[22\] _12598_ _03086_ _03087_ VGND VGND VPWR
+ VPWR _03088_ sky130_fd_sc_hd__a22o_1
X_14895_ _10912_ _10913_ _10921_ _10931_ VGND VGND VPWR VPWR _10932_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_187_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19422_ _04471_ _04289_ _04056_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16634_ _12598_ VGND VGND VPWR VPWR _12599_ sky130_fd_sc_hd__clkbuf_4
X_13846_ net481 _10167_ _10168_ _10162_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19353_ _04635_ _04636_ _04446_ _04643_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16565_ _12529_ VGND VGND VPWR VPWR _12530_ sky130_fd_sc_hd__clkbuf_4
X_13777_ memory.csr_read_data_out_reg\[26\] _09987_ _10115_ VGND VGND VPWR VPWR _10116_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_174_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18304_ _03617_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__clkbuf_1
X_15516_ _11497_ _11506_ _11507_ VGND VGND VPWR VPWR _11508_ sky130_fd_sc_hd__o21ai_1
X_19284_ _04346_ _04569_ _04575_ _04577_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16496_ _11042_ decode.regfile.registers_4\[31\] _11190_ _10628_ _11083_ VGND VGND
+ VPWR VPWR _12462_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18235_ csr._mcycle_T_3\[57\] csr._mcycle_T_3\[56\] csr._mcycle_T_3\[55\] csr._mcycle_T_3\[54\]
+ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__or4_1
X_15447_ _10960_ decode.regfile.registers_28\[3\] _11067_ _11038_ _11440_ VGND VGND
+ VPWR VPWR _11441_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_212_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18166_ _03463_ _03464_ _10921_ decode.control.io_funct7\[2\] VGND VGND VPWR VPWR
+ _03511_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_5_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15378_ _11370_ _11372_ _11296_ VGND VGND VPWR VPWR _11373_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17117_ _13071_ _13072_ _13073_ VGND VGND VPWR VPWR _13074_ sky130_fd_sc_hd__a21o_1
X_14329_ _10092_ _10444_ VGND VGND VPWR VPWR _10449_ sky130_fd_sc_hd__nand2_1
Xhold405 decode.regfile.registers_13\[2\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__dlygate4sd3_1
X_18097_ _03469_ _03467_ _03474_ net2024 VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_106_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold416 decode.regfile.registers_21\[11\] VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_225_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold427 decode.regfile.registers_6\[8\] VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 decode.regfile.registers_30\[1\] VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold449 decode.regfile.registers_22\[28\] VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ _10931_ net2640 _12487_ VGND VGND VPWR VPWR _13007_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1105 decode.regfile.registers_14\[15\] VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__dlygate4sd3_1
X_18999_ decode.id_ex_rs2_data_reg\[4\] _03747_ _04030_ _03764_ VGND VGND VPWR VPWR
+ _04298_ sky130_fd_sc_hd__o22a_2
Xhold1116 fetch.bht.bhtTable_target_pc\[13\]\[26\] VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1127 fetch.bht.bhtTable_target_pc\[14\]\[24\] VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 fetch.bht.bhtTable_tag\[3\]\[12\] VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1149 fetch.bht.bhtTable_tag\[13\]\[22\] VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20961_ _05962_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_176_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22700_ csr._mcycle_T_2\[24\] _07236_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_176_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23680_ net861 csr.io_mem_pc\[31\] _07983_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_1343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20892_ _05857_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22631_ net1524 _07196_ _07197_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_172_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_172_Left_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25350_ _09964_ _08907_ VGND VGND VPWR VPWR _08909_ sky130_fd_sc_hd__nand2_1
X_22562_ csr._minstret_T_3\[38\] csr._minstret_T_3\[37\] csr._minstret_T_3\[36\] _07144_
+ _07148_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__a41o_1
XFILLER_0_158_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24301_ _08326_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__clkbuf_1
XINSDIODE1_380 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21513_ _06250_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25281_ _08869_ decode.regfile.registers_0\[2\] VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22493_ _10757_ _07087_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_135_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1095 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27020_ clknet_leaf_338_clock _00049_ VGND VGND VPWR VPWR decode.regfile.registers_22\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24232_ _08060_ net2061 _08289_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21444_ _06237_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24163_ _06250_ VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21375_ _06200_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23114_ net226 _07536_ _07537_ _07554_ _07535_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_9_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20326_ _10693_ _10725_ _05490_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24094_ _08219_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__clkbuf_1
X_28971_ clknet_leaf_94_clock _01984_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold950 fetch.bht.bhtTable_tag\[1\]\[13\] VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 fetch.bht.bhtTable_target_pc\[2\]\[15\] VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 fetch.bht.bhtTable_target_pc\[13\]\[5\] VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_181_Left_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23045_ fetch.bht.bhtTable_target_pc\[12\]\[9\] fetch.bht.bhtTable_target_pc\[13\]\[9\]
+ fetch.bht.bhtTable_target_pc\[14\]\[9\] fetch.bht.bhtTable_target_pc\[15\]\[9\]
+ _07407_ _07115_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__mux4_1
X_27922_ clknet_leaf_67_clock _00951_ VGND VGND VPWR VPWR csr.io_csr_write_address\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold983 fetch.bht.bhtTable_target_pc\[10\]\[16\] VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__dlygate4sd3_1
X_20257_ _05439_ _05443_ _05425_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_34_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold994 decode.regfile.registers_6\[15\] VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27853_ clknet_leaf_322_clock _00882_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20188_ _05374_ _05380_ _05381_ decode.id_ex_pc_reg\[26\] decode.id_ex_imm_reg\[26\]
+ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_129_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2340 decode.regfile.registers_1\[10\] VGND VGND VPWR VPWR net2567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2351 decode.regfile.registers_0\[9\] VGND VGND VPWR VPWR net2578 sky130_fd_sc_hd__dlygate4sd3_1
X_26804_ _09406_ _09763_ VGND VGND VPWR VPWR _09773_ sky130_fd_sc_hd__nand2_1
Xhold2362 decode.regfile.registers_3\[18\] VGND VGND VPWR VPWR net2589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27784_ clknet_leaf_334_clock _00813_ VGND VGND VPWR VPWR memory.io_wb_readdata\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2373 decode.regfile.registers_17\[31\] VGND VGND VPWR VPWR net2600 sky130_fd_sc_hd__dlygate4sd3_1
X_24996_ csr._mcycle_T_2\[3\] _08710_ _08709_ csr.mcycle\[3\] VGND VGND VPWR VPWR
+ _08711_ sky130_fd_sc_hd__a211oi_1
Xhold2384 decode.regfile.registers_27\[23\] VGND VGND VPWR VPWR net2611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1650 decode.regfile.registers_16\[21\] VGND VGND VPWR VPWR net1877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2395 decode.regfile.registers_0\[28\] VGND VGND VPWR VPWR net2622 sky130_fd_sc_hd__dlygate4sd3_1
X_29523_ clknet_leaf_265_clock _02536_ VGND VGND VPWR VPWR decode.regfile.registers_8\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1661 csr.mcycle\[3\] VGND VGND VPWR VPWR net1888 sky130_fd_sc_hd__dlygate4sd3_1
X_26735_ _09708_ VGND VGND VPWR VPWR _09733_ sky130_fd_sc_hd__buf_2
X_23947_ net987 _08105_ _06156_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1672 execute.csr_write_address_out_reg\[9\] VGND VGND VPWR VPWR net1899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1683 fetch.bht.bhtTable_tag\[6\]\[21\] VGND VGND VPWR VPWR net1910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1694 fetch.bht.bhtTable_target_pc\[0\]\[22\] VGND VGND VPWR VPWR net1921 sky130_fd_sc_hd__dlygate4sd3_1
X_13700_ _10021_ memory.io_wb_readdata\[14\] _10001_ memory.io_wb_reg_pc\[14\] _10050_
+ VGND VGND VPWR VPWR _10051_ sky130_fd_sc_hd__a221oi_2
X_14680_ execute.io_target_pc\[30\] _10684_ VGND VGND VPWR VPWR _10723_ sky130_fd_sc_hd__or2_1
X_29454_ clknet_leaf_261_clock _02467_ VGND VGND VPWR VPWR decode.regfile.registers_6\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_23878_ _08106_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26666_ net2338 _09692_ _09693_ _09688_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_190_Left_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28405_ clknet_leaf_141_clock _01418_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13631_ memory.io_wb_reg_pc\[5\] _09978_ _09977_ _09990_ VGND VGND VPWR VPWR _09991_
+ sky130_fd_sc_hd__a211o_1
X_22829_ _07310_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__clkbuf_1
X_25617_ _08916_ _09069_ VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__nand2_1
X_29385_ clknet_leaf_259_clock _02398_ VGND VGND VPWR VPWR decode.regfile.registers_4\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_26597_ net2248 _09649_ _09653_ _09648_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28336_ clknet_leaf_238_clock _01349_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13562_ csr.io_mem_pc\[4\] csr.io_mem_pc\[2\] csr.io_mem_pc\[3\] VGND VGND VPWR VPWR
+ _09928_ sky130_fd_sc_hd__and3_1
X_16350_ decode.regfile.registers_5\[27\] _11192_ _11138_ VGND VGND VPWR VPWR _12320_
+ sky130_fd_sc_hd__and3_1
X_25548_ _09023_ VGND VGND VPWR VPWR _09036_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_181_Right_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15301_ net346 VGND VGND VPWR VPWR _11297_ sky130_fd_sc_hd__buf_4
XFILLER_0_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16281_ decode.regfile.registers_10\[25\] _10637_ _11131_ _11315_ VGND VGND VPWR
+ VPWR _12253_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_229_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28267_ clknet_leaf_64_clock _01289_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_25479_ net1455 _08995_ _08996_ _08991_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_229_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18020_ _03414_ _03415_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15232_ _11228_ VGND VGND VPWR VPWR _11229_ sky130_fd_sc_hd__clkbuf_4
X_27218_ clknet_leaf_7_clock _00247_ VGND VGND VPWR VPWR decode.regfile.registers_29\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28198_ clknet_leaf_64_clock _01220_ VGND VGND VPWR VPWR csr.mscratch\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15163_ decode.regfile.registers_2\[0\] _10647_ _11149_ _11152_ _11159_ VGND VGND
+ VPWR VPWR _11160_ sky130_fd_sc_hd__o311a_1
XFILLER_0_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27149_ clknet_leaf_330_clock _00178_ VGND VGND VPWR VPWR decode.regfile.registers_26\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14114_ _10122_ _10312_ VGND VGND VPWR VPWR _10324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19971_ _05216_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15094_ decode.immGen._imm_T_24\[3\] decode.immGen._imm_T_24\[2\] VGND VGND VPWR
+ VPWR _11091_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14045_ net2207 _10244_ _10283_ _10275_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__o211a_1
X_18922_ _03781_ _03788_ _03795_ _03800_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__o22a_1
XFILLER_0_157_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18853_ _03707_ decode.id_ex_imm_reg\[11\] _04151_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17804_ decode.regfile.registers_14\[25\] _12670_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18784_ decode.id_ex_rs2_data_reg\[14\] _03746_ _04077_ _03764_ _04082_ VGND VGND
+ VPWR VPWR _04083_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_175_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15996_ _11076_ _11090_ decode.regfile.registers_25\[17\] _11945_ _11975_ VGND VGND
+ VPWR VPWR _11976_ sky130_fd_sc_hd__o32a_1
XFILLER_0_59_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17735_ _13339_ _03136_ _03137_ _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14947_ decode.control.io_opcode\[2\] decode.control.io_opcode\[1\] decode.control.io_opcode\[0\]
+ _10583_ _10952_ VGND VGND VPWR VPWR _10975_ sky130_fd_sc_hd__a41o_1
XFILLER_0_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17666_ _02997_ _13262_ _13182_ decode.regfile.registers_29\[21\] _03071_ VGND VGND
+ VPWR VPWR _03072_ sky130_fd_sc_hd__o221a_1
XFILLER_0_159_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14878_ _10918_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19405_ _03639_ _04165_ _04620_ _04303_ _04693_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__o32a_1
X_16617_ _12581_ VGND VGND VPWR VPWR _12582_ sky130_fd_sc_hd__clkbuf_4
X_13829_ net1301 _10153_ _10158_ _10132_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__o211a_1
X_17597_ decode.regfile.registers_4\[20\] _12548_ _13145_ decode.regfile.registers_5\[20\]
+ _12614_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_214_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19336_ _03972_ _03974_ _04007_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16548_ _10595_ _10606_ _11012_ _12512_ VGND VGND VPWR VPWR _12513_ sky130_fd_sc_hd__or4_2
XFILLER_0_58_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19267_ _04050_ _04051_ _04516_ _04529_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__o22a_1
X_16479_ _11260_ _12443_ _12444_ _12445_ VGND VGND VPWR VPWR _12446_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18218_ _03553_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19198_ _04009_ _04493_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18149_ _03495_ _03493_ _03500_ net2154 VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_142_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold202 decode.regfile.registers_31\[4\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold213 decode.regfile.registers_29\[17\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 decode.control.io_funct7\[2\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold235 _10677_ VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
X_21160_ _05866_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__clkbuf_2
Xhold246 decode.regfile.registers_6\[14\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold257 decode.regfile.registers_27\[9\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_165_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold268 fetch.bht.bhtTable_valid\[10\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
X_20111_ _05296_ _05305_ _05311_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__nand3_1
XFILLER_0_106_1153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_165_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold279 decode.regfile.registers_23\[14\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21091_ net2743 _09925_ _06031_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__and4bb_1
X_20042_ decode.id_ex_imm_reg\[3\] _10747_ _05250_ _05251_ VGND VGND VPWR VPWR _05263_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_77_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24850_ _06128_ net2115 _08607_ VGND VGND VPWR VPWR _08613_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23801_ _08054_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24781_ _08074_ net1375 _08574_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__mux2_1
X_21993_ _06571_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23732_ _08017_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__clkbuf_1
X_26520_ net2051 _09605_ _09609_ _09608_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__o211a_1
XANTENNA_108 net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20944_ _05953_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_119 _09128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23663_ net1596 csr.io_mem_pc\[23\] _07972_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__mux2_1
X_26451_ net2709 _09561_ _09569_ _09567_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20875_ net124 _05915_ _05911_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__and3_1
X_22614_ net1512 _07185_ _07186_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__o21a_1
X_25402_ net1761 _08928_ _08944_ _08927_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__o211a_1
X_29170_ clknet_leaf_184_clock _02183_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26382_ _09438_ _09490_ VGND VGND VPWR VPWR _09529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23594_ _06124_ net1565 _07941_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28121_ clknet_leaf_90_clock _01143_ VGND VGND VPWR VPWR csr.minstret\[26\] sky130_fd_sc_hd__dfxtp_1
X_25333_ _08897_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22545_ net2560 _07136_ _07137_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25264_ _08103_ net1668 _09906_ VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__mux2_1
X_28052_ clknet_leaf_213_clock _01074_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22476_ _07070_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24215_ _08109_ net1303 _06251_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27003_ clknet_leaf_343_clock _00032_ VGND VGND VPWR VPWR decode.regfile.registers_22\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_21427_ _06228_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25195_ net423 _08826_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24146_ _08246_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__clkbuf_1
X_21358_ _06191_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__clkbuf_1
X_20309_ _05340_ _10867_ _05473_ _10798_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_57_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28954_ clknet_leaf_128_clock _01967_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_24077_ net860 execute.io_target_pc\[26\] _07991_ VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold780 fetch.bht.bhtTable_target_pc\[2\]\[31\] VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__dlygate4sd3_1
X_21289_ _06152_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold791 fetch.bht.bhtTable_tag\[11\]\[18\] VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23028_ _07471_ _07472_ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__nor2_1
X_27905_ clknet_leaf_18_clock _00934_ VGND VGND VPWR VPWR csr._mcycle_T_2\[26\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_200_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28885_ clknet_leaf_116_clock _01898_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _11571_ net2787 _11722_ _11723_ _11724_ VGND VGND VPWR VPWR _11833_ sky130_fd_sc_hd__o2111a_1
X_27836_ clknet_leaf_325_clock _00865_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2170 decode.regfile.registers_2\[15\] VGND VGND VPWR VPWR net2397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14801_ decode.id_ex_pc_reg\[13\] _10810_ _10814_ _10689_ _10843_ VGND VGND VPWR
+ VPWR _10844_ sky130_fd_sc_hd__o221a_1
Xhold2181 decode.regfile.registers_1\[28\] VGND VGND VPWR VPWR net2408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2192 decode.regfile.registers_9\[26\] VGND VGND VPWR VPWR net2419 sky130_fd_sc_hd__dlygate4sd3_1
X_15781_ decode.regfile.registers_0\[12\] _11154_ _11190_ _11298_ VGND VGND VPWR VPWR
+ _11766_ sky130_fd_sc_hd__o2bb2ai_1
X_27767_ clknet_leaf_323_clock _00796_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_24979_ csr._mcycle_T_3\[62\] csr._mcycle_T_3\[61\] _08696_ VGND VGND VPWR VPWR _08699_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1480 fetch.bht.bhtTable_tag\[9\]\[24\] VGND VGND VPWR VPWR net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17520_ decode.regfile.registers_11\[18\] _12595_ _12583_ _12551_ _13466_ VGND VGND
+ VPWR VPWR _13467_ sky130_fd_sc_hd__a221o_1
X_29506_ clknet_leaf_252_clock _02519_ VGND VGND VPWR VPWR decode.regfile.registers_8\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1491 fetch.bht.bhtTable_tag\[7\]\[11\] VGND VGND VPWR VPWR net1718 sky130_fd_sc_hd__dlygate4sd3_1
X_14732_ _10772_ _10773_ _10774_ VGND VGND VPWR VPWR _10775_ sky130_fd_sc_hd__and3_1
X_26718_ _09396_ _09720_ VGND VGND VPWR VPWR _09724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27698_ clknet_leaf_22_clock _00727_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17451_ decode.regfile.registers_18\[16\] _12571_ _12561_ _13399_ VGND VGND VPWR
+ VPWR _13400_ sky130_fd_sc_hd__a211o_1
X_29437_ clknet_leaf_249_clock _02450_ VGND VGND VPWR VPWR decode.regfile.registers_6\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14663_ decode.id_ex_pc_reg\[9\] VGND VGND VPWR VPWR _10706_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26649_ net499 _09679_ _09683_ _09675_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16402_ _11263_ _11217_ _11085_ decode.regfile.registers_21\[28\] _11648_ VGND VGND
+ VPWR VPWR _12371_ sky130_fd_sc_hd__o32a_1
XFILLER_0_200_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13614_ _09975_ _09951_ VGND VGND VPWR VPWR _09976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29368_ clknet_leaf_246_clock _02381_ VGND VGND VPWR VPWR decode.regfile.registers_3\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_17382_ _10938_ decode.regfile.registers_25\[14\] _12505_ _12811_ VGND VGND VPWR
+ VPWR _13333_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14594_ _10636_ VGND VGND VPWR VPWR _10637_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19121_ _04297_ _04261_ _04263_ _04260_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__a211o_1
X_28319_ clknet_leaf_208_clock _01332_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_16333_ _10958_ decode.regfile.registers_26\[26\] _11676_ _11338_ _11564_ VGND VGND
+ VPWR VPWR _12304_ sky130_fd_sc_hd__o2111a_1
X_13545_ _09914_ _09892_ _09916_ net389 VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29299_ clknet_leaf_225_clock _02312_ VGND VGND VPWR VPWR decode.regfile.registers_1\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19052_ _03888_ _03944_ _04230_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16264_ _12133_ net478 _12202_ _12236_ _12132_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__o221a_1
XFILLER_0_125_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18003_ _11014_ _10936_ decode.regfile.registers_23\[30\] _12995_ VGND VGND VPWR
+ VPWR _03400_ sky130_fd_sc_hd__or4_1
X_15215_ decode.regfile.registers_17\[0\] _11094_ _11114_ _11119_ _11211_ VGND VGND
+ VPWR VPWR _11212_ sky130_fd_sc_hd__a41o_1
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16195_ _11942_ decode.regfile.registers_30\[23\] _12095_ _12096_ _12097_ VGND VGND
+ VPWR VPWR _12169_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_129_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15146_ decode.immGen._imm_T_24\[4\] decode.immGen._imm_T_24\[1\] VGND VGND VPWR
+ VPWR _11143_ sky130_fd_sc_hd__nor2_4
XFILLER_0_65_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19954_ _05211_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__clkbuf_1
X_15077_ _11073_ VGND VGND VPWR VPWR _11074_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_207_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_207_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14028_ _10131_ VGND VGND VPWR VPWR _10275_ sky130_fd_sc_hd__clkbuf_4
X_18905_ _04203_ _03902_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__nand2_2
X_19885_ _04589_ _05143_ _05152_ _05154_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_219_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_343_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_343_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_160_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18836_ net131 _03664_ _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_199_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_999 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18767_ execute.csr_read_data_out_reg\[6\] _03661_ _03660_ VGND VGND VPWR VPWR _04066_
+ sky130_fd_sc_hd__or3_1
X_15979_ _11951_ _11958_ _11135_ VGND VGND VPWR VPWR _11959_ sky130_fd_sc_hd__o21ai_1
X_17718_ _10610_ _12626_ _03117_ _03118_ _03121_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__o32a_1
XFILLER_0_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18698_ _03990_ _03991_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__nand3_4
Xclkbuf_leaf_358_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_358_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17649_ decode.regfile.registers_17\[21\] _12579_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20660_ csr._minstret_T_3\[63\] _05577_ _05578_ _05563_ csr._csr_read_data_T_9\[31\]
+ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19319_ _04075_ _04172_ _04585_ _04553_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_133_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20591_ csr.mcycle\[21\] _05587_ _05575_ csr.minstret\[21\] VGND VGND VPWR VPWR _05730_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22330_ fetch.bht.bhtTable_tag\[0\]\[8\] fetch.bht.bhtTable_tag\[1\]\[8\] fetch.bht.bhtTable_tag\[2\]\[8\]
+ fetch.bht.bhtTable_tag\[3\]\[8\] _06878_ _06621_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22261_ fetch.bht.bhtTable_tag\[12\]\[17\] fetch.bht.bhtTable_tag\[13\]\[17\] _06643_
+ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24000_ net1620 VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21212_ _06100_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__clkbuf_1
X_22192_ fetch.bht.bhtTable_tag\[4\]\[5\] fetch.bht.bhtTable_tag\[5\]\[5\] fetch.bht.bhtTable_tag\[6\]\[5\]
+ fetch.bht.bhtTable_tag\[7\]\[5\] _06700_ _06685_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21143_ _06062_ _06058_ net1691 VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21074_ _06023_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__clkbuf_1
X_25951_ net2322 _09256_ _09268_ _09264_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_126_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20025_ decode.id_ex_imm_reg\[4\] decode.id_ex_pc_reg\[4\] VGND VGND VPWR VPWR _05248_
+ sky130_fd_sc_hd__nor2_1
X_24902_ csr._mcycle_T_3\[34\] csr._mcycle_T_3\[33\] csr._mcycle_T_3\[32\] _08636_
+ VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__and4_1
X_28670_ clknet_leaf_173_clock _01683_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_25882_ net2602 _09226_ _09228_ _09222_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27621_ clknet_leaf_146_clock _00650_ VGND VGND VPWR VPWR execute.io_target_pc\[30\]
+ sky130_fd_sc_hd__dfxtp_4
X_24833_ _06111_ net1535 _08422_ VGND VGND VPWR VPWR _08604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27552_ clknet_leaf_42_clock _00581_ VGND VGND VPWR VPWR execute.io_mem_memtoreg\[0\]
+ sky130_fd_sc_hd__dfxtp_4
X_24764_ _08057_ net1820 _08563_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21976_ net1778 _06588_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer50 net276 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_29_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer61 _09928_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_1
X_26503_ net745 _09592_ _09599_ _09595_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__o211a_1
X_23715_ _08008_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer72 _06679_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20927_ _05937_ _05933_ net49 VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24695_ _06282_ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__clkbuf_8
X_27483_ clknet_leaf_72_clock _00512_ VGND VGND VPWR VPWR csr.mtip sky130_fd_sc_hd__dfxtp_1
Xrebuffer83 net309 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_1
Xrebuffer94 net320 VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_84_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29222_ clknet_leaf_87_clock _02235_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26434_ net2393 _09548_ _09559_ _09553_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__o211a_1
X_23646_ net823 _10807_ _07961_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20858_ _05906_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29153_ clknet_leaf_238_clock _02166_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23577_ _07933_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__clkbuf_1
X_26365_ _09422_ _09515_ VGND VGND VPWR VPWR _09520_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20789_ execute.io_mem_rd\[0\] _05867_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28104_ clknet_leaf_75_clock _01126_ VGND VGND VPWR VPWR csr.minstret\[9\] sky130_fd_sc_hd__dfxtp_1
X_22528_ _06633_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__buf_4
X_25316_ _08888_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__clkbuf_1
X_29084_ clknet_leaf_72_clock net1801 VGND VGND VPWR VPWR csr._mcycle_T_3\[32\] sky130_fd_sc_hd__dfxtp_1
X_26296_ _09428_ _09472_ VGND VGND VPWR VPWR _09480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28035_ clknet_leaf_190_clock _01057_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25247_ _08853_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__clkbuf_1
X_22459_ _06754_ fetch.btb.btbTable\[5\]\[1\] fetch.bht.bhtTable_valid\[5\] _06686_
+ _07053_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__a311o_1
XFILLER_0_84_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15000_ _10589_ VGND VGND VPWR VPWR _11012_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25178_ _09884_ _08808_ _09881_ VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24129_ net1130 execute.io_target_pc\[19\] _08232_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28937_ clknet_leaf_88_clock _01950_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16951_ _11015_ _10937_ decode.regfile.registers_23\[4\] _12520_ VGND VGND VPWR VPWR
+ _12912_ sky130_fd_sc_hd__or4_1
X_15902_ decode.regfile.registers_2\[15\] _11503_ _11148_ _11152_ _11883_ VGND VGND
+ VPWR VPWR _11884_ sky130_fd_sc_hd__o311a_1
XFILLER_0_60_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19670_ _04539_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_216_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28868_ clknet_leaf_131_clock _01881_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16882_ decode.regfile.registers_7\[3\] _12610_ _12737_ decode.regfile.registers_6\[3\]
+ _12843_ VGND VGND VPWR VPWR _12844_ sky130_fd_sc_hd__a221oi_1
X_18621_ _03797_ _03916_ _03889_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15833_ _11276_ _11815_ _11816_ VGND VGND VPWR VPWR _11817_ sky130_fd_sc_hd__o21a_1
X_27819_ clknet_leaf_321_clock _00848_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_28799_ clknet_leaf_179_clock _01812_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18552_ _03850_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_194_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ decode.regfile.registers_22\[11\] _11228_ _11262_ _11749_ VGND VGND VPWR
+ VPWR _11750_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_194_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17503_ _12708_ net411 _13415_ _13450_ _13219_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__o221a_1
XFILLER_0_213_1321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14715_ csr.io_trapped csr.io_mret _10757_ VGND VGND VPWR VPWR _10758_ sky130_fd_sc_hd__or3_2
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18483_ _10194_ _03755_ _03735_ _03736_ _03738_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_185_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15695_ _11403_ _11678_ _11680_ _11682_ VGND VGND VPWR VPWR _11683_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_190_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17434_ _12631_ decode.regfile.registers_0\[16\] VGND VGND VPWR VPWR _13383_ sky130_fd_sc_hd__nand2_1
X_14646_ decode.id_ex_pc_reg\[11\] VGND VGND VPWR VPWR _10689_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_170_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17365_ _13312_ _13314_ _13315_ VGND VGND VPWR VPWR _13316_ sky130_fd_sc_hd__o21ai_1
XANTENNA_19 _05488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14577_ _10619_ decode.id_ex_ex_rd_reg\[0\] VGND VGND VPWR VPWR _10620_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19104_ _04006_ _04228_ _04231_ _04401_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16316_ decode.regfile.registers_9\[26\] _11365_ _12278_ _12286_ VGND VGND VPWR VPWR
+ _12287_ sky130_fd_sc_hd__a2bb2oi_1
X_13528_ _09900_ _09880_ _09883_ _09890_ VGND VGND VPWR VPWR _09905_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17296_ _13081_ _13168_ decode.regfile.registers_23\[12\] _13041_ VGND VGND VPWR
+ VPWR _13249_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19035_ decode.id_ex_rs1_data_reg\[11\] _03689_ _04145_ _03701_ _04148_ VGND VGND
+ VPWR VPWR _04334_ sky130_fd_sc_hd__o221ai_4
X_16247_ _10639_ _11143_ _11036_ _12206_ _12219_ VGND VGND VPWR VPWR _12220_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_209_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput104 net104 VGND VGND VPWR VPWR io_memory_address[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput115 net115 VGND VGND VPWR VPWR io_memory_address[23] sky130_fd_sc_hd__clkbuf_4
X_16178_ decode.regfile.registers_13\[22\] _10642_ _11187_ _12151_ _12152_ VGND VGND
+ VPWR VPWR _12153_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput126 net126 VGND VGND VPWR VPWR io_memory_address[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput137 net137 VGND VGND VPWR VPWR io_memory_write_data[10] sky130_fd_sc_hd__clkbuf_4
X_15129_ _11058_ _10632_ _11047_ _11125_ VGND VGND VPWR VPWR _11126_ sky130_fd_sc_hd__or4_4
XFILLER_0_50_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput148 net148 VGND VGND VPWR VPWR io_memory_write_data[20] sky130_fd_sc_hd__clkbuf_4
Xoutput159 net159 VGND VGND VPWR VPWR io_memory_write_data[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_282_clock clknet_5_20__leaf_clock VGND VGND VPWR VPWR clknet_leaf_282_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19937_ _05202_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19868_ _04251_ _04252_ _05091_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18819_ _04115_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__inv_2
X_19799_ _04325_ _05034_ _05071_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_121_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_297_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_297_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21830_ _06480_ net662 _06316_ _06472_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_222_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21761_ _06443_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_220_clock clknet_5_31__leaf_clock VGND VGND VPWR VPWR clknet_leaf_220_clock
+ sky130_fd_sc_hd__clkbuf_8
X_23500_ _10670_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20712_ _05809_ decode.id_ex_rs1_data_reg\[15\] _05798_ VGND VGND VPWR VPWR _05825_
+ sky130_fd_sc_hd__a21oi_1
X_24480_ _08107_ net1654 _08411_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21692_ csr.minstret\[25\] _06381_ _06391_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23431_ _10965_ _07847_ _05206_ VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__or3b_1
XFILLER_0_176_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20643_ _05771_ _05774_ _05630_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_119_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26150_ net757 _09373_ _09384_ _09370_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__o211a_1
X_23362_ _07619_ _07573_ _07620_ _07787_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__a31o_1
XFILLER_0_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20574_ csr._csr_read_data_T_8\[18\] _05622_ _05712_ _05715_ VGND VGND VPWR VPWR
+ _05716_ sky130_fd_sc_hd__a211o_2
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25101_ _06117_ net1938 _08778_ VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__mux2_1
X_22313_ fetch.bht.bhtTable_tag\[12\]\[0\] fetch.bht.bhtTable_tag\[13\]\[0\] fetch.bht.bhtTable_tag\[14\]\[0\]
+ fetch.bht.bhtTable_tag\[15\]\[0\] _06617_ _06622_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_235_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_235_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26081_ _09328_ VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__buf_2
X_23293_ fetch.bht.bhtTable_target_pc\[0\]\[23\] fetch.bht.bhtTable_target_pc\[1\]\[23\]
+ fetch.bht.bhtTable_target_pc\[2\]\[23\] fetch.bht.bhtTable_target_pc\[3\]\[23\]
+ _07555_ _07710_ VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25032_ csr.mcycle\[15\] _08733_ VGND VGND VPWR VPWR _08735_ sky130_fd_sc_hd__nand2_1
X_22244_ fetch.bht.bhtTable_tag\[6\]\[19\] fetch.bht.bhtTable_tag\[7\]\[19\] _06707_
+ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29840_ clknet_leaf_298_clock _02853_ VGND VGND VPWR VPWR decode.regfile.registers_18\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_22175_ fetch.bht.bhtTable_tag\[6\]\[25\] fetch.bht.bhtTable_tag\[7\]\[25\] _06619_
+ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21126_ _06055_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__clkbuf_1
X_29771_ clknet_leaf_293_clock _02784_ VGND VGND VPWR VPWR decode.regfile.registers_16\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26983_ _10127_ _09838_ VGND VGND VPWR VPWR _09875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_1324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28722_ clknet_leaf_106_clock _01735_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25934_ net729 _09256_ _09258_ _09250_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__o211a_1
X_21057_ execute.csr_read_data_out_reg\[17\] _06014_ _06010_ VGND VGND VPWR VPWR _06015_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20008_ decode.id_ex_imm_reg\[2\] _10834_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__nor2_1
X_28653_ clknet_leaf_101_clock _01666_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25865_ net695 _09213_ _09218_ _09209_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27604_ clknet_leaf_158_clock _00633_ VGND VGND VPWR VPWR execute.io_target_pc\[13\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_92_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24816_ _08109_ net1864 _08585_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28584_ clknet_leaf_103_clock _01597_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25796_ net501 _09170_ _09178_ _09169_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27535_ clknet_leaf_318_clock _00564_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_2
X_24747_ _08109_ net1817 _06283_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_209 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21959_ csr._mcycle_T_2\[4\] _06572_ _06581_ _06579_ VGND VGND VPWR VPWR _01224_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_48_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ net634 _10507_ _10545_ _10546_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_104_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _11194_ decode.regfile.registers_12\[4\] decode.regfile.registers_13\[4\]
+ _11195_ _11198_ VGND VGND VPWR VPWR _11473_ sky130_fd_sc_hd__o221a_1
X_27466_ clknet_leaf_31_clock _00495_ VGND VGND VPWR VPWR csr.io_csr_address\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_104_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24678_ _08522_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_13_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29205_ clknet_leaf_163_clock _02218_ VGND VGND VPWR VPWR fetch.btb.btbTable\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26417_ _09398_ _09545_ VGND VGND VPWR VPWR _09550_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _09950_ _10507_ VGND VGND VPWR VPWR _10508_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23629_ _07962_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27397_ clknet_leaf_27_clock _00426_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_193_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29136_ clknet_leaf_80_clock _02149_ VGND VGND VPWR VPWR csr.mcycle\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17150_ decode.regfile.registers_4\[9\] _12618_ _12620_ decode.regfile.registers_5\[9\]
+ _12622_ VGND VGND VPWR VPWR _13106_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26348_ _09404_ _09502_ VGND VGND VPWR VPWR _09510_ sky130_fd_sc_hd__nand2_1
X_14362_ net604 _10463_ _10467_ _10468_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__o211a_1
Xinput17 io_fetch_data[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_0_141_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 net658 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
X_16101_ decode.regfile.registers_16\[20\] _11203_ _12076_ _12077_ VGND VGND VPWR
+ VPWR _12078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 io_memory_read_data[14] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_1
XFILLER_0_52_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29067_ clknet_leaf_212_clock _02080_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_17081_ decode.regfile.registers_21\[7\] _12682_ _12909_ VGND VGND VPWR VPWR _13039_
+ sky130_fd_sc_hd__o21a_1
X_14293_ net510 _10419_ _10428_ _10427_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26279_ _09410_ _09459_ VGND VGND VPWR VPWR _09470_ sky130_fd_sc_hd__nand2_1
X_28018_ clknet_leaf_220_clock _01040_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16032_ _11075_ _12009_ _12010_ _11486_ VGND VGND VPWR VPWR _12011_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_204_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17983_ decode.regfile.registers_13\[30\] _12927_ _12583_ VGND VGND VPWR VPWR _03380_
+ sky130_fd_sc_hd__and3_1
X_19722_ _04974_ _04977_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16934_ decode.regfile.registers_10\[4\] _12654_ _12878_ _12894_ VGND VGND VPWR VPWR
+ _12895_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_196_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19653_ _04866_ _04928_ _04931_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_221_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16865_ decode.regfile.registers_17\[3\] _11022_ _12567_ _12586_ _12570_ VGND VGND
+ VPWR VPWR _12827_ sky130_fd_sc_hd__a41o_1
X_18604_ _03898_ _03899_ _03902_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__or3_1
XFILLER_0_205_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15816_ net323 _11167_ decode.regfile.registers_10\[13\] _11381_ VGND VGND VPWR VPWR
+ _11800_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_137_1252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19584_ _04745_ _04828_ _04831_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a21boi_2
X_16796_ _12494_ decode.regfile.registers_26\[1\] _12759_ _11010_ _11026_ VGND VGND
+ VPWR VPWR _12760_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18535_ _03656_ _03832_ _03701_ _03833_ _03670_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15747_ _11729_ _11731_ _11732_ VGND VGND VPWR VPWR _11733_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_172_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18466_ decode.id_ex_rs2_data_reg\[31\] _03747_ _03690_ _03764_ VGND VGND VPWR VPWR
+ _03765_ sky130_fd_sc_hd__o22a_1
X_15678_ _11123_ decode.regfile.registers_16\[9\] _11126_ _11665_ VGND VGND VPWR VPWR
+ _11666_ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17417_ _12546_ VGND VGND VPWR VPWR _13367_ sky130_fd_sc_hd__buf_2
X_14629_ _10671_ VGND VGND VPWR VPWR _10672_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_151_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18397_ _03680_ _09929_ decode.io_wb_rd\[4\] _03652_ VGND VGND VPWR VPWR _03696_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_157_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17348_ _13221_ _13297_ _13298_ _13299_ VGND VGND VPWR VPWR _13300_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17279_ _12649_ _12615_ _13231_ VGND VGND VPWR VPWR _13232_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19018_ _04316_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20290_ _05467_ _05468_ _05420_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_228_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_228_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23980_ net785 execute.io_target_pc\[11\] _08153_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22931_ csr._csr_read_data_T_8\[2\] _06039_ csr.io_mret_vector\[2\] _06463_ _07381_
+ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_15__f_clock clknet_2_1_0_clock VGND VGND VPWR VPWR clknet_5_15__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_84_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25650_ net2599 _09082_ _09094_ _09087_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__o211a_1
X_22862_ _07327_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24601_ net899 execute.io_target_pc\[22\] _08473_ VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_179_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21813_ _06477_ _10019_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__and2_1
XFILLER_0_211_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22793_ _07291_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__clkbuf_1
X_25581_ _08956_ _09049_ VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_210_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27320_ clknet_leaf_31_clock _00349_ VGND VGND VPWR VPWR decode.id_ex_ex_rs1_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24532_ _08447_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__clkbuf_1
X_21744_ _06434_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27251_ clknet_leaf_31_clock _00280_ VGND VGND VPWR VPWR decode.regfile.registers_30\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_24463_ _08387_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__clkbuf_8
X_21675_ csr.minstret\[19\] csr.minstret\[20\] _06375_ VGND VGND VPWR VPWR _06383_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_136_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_174_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_174_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_190_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26202_ net2671 _09419_ _09421_ _09418_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__o211a_1
X_23414_ fetch.bht.bhtTable_target_pc\[4\]\[31\] fetch.bht.bhtTable_target_pc\[5\]\[31\]
+ _07066_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__mux2_1
X_20626_ csr.mcycle\[26\] _05587_ _05594_ csr.minstret\[26\] VGND VGND VPWR VPWR _05760_
+ sky130_fd_sc_hd__a22o_1
X_24394_ _08374_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__clkbuf_1
X_27182_ clknet_leaf_3_clock _00211_ VGND VGND VPWR VPWR decode.regfile.registers_27\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23345_ _07064_ _07770_ _07771_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26133_ _09372_ VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__clkbuf_4
X_20557_ csr.mcycle\[16\] _05587_ _05559_ csr.minstret\[16\] VGND VGND VPWR VPWR _05701_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23276_ _03500_ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__buf_2
XFILLER_0_132_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26064_ _08910_ _09330_ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__nand2_1
X_20488_ csr._minstret_T_3\[39\] _05555_ _05599_ csr.pie _05559_ VGND VGND VPWR VPWR
+ _05641_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_189_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_189_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22227_ _06785_ _06808_ _06820_ _06821_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__nand4b_2
X_25015_ net1155 _08722_ _08723_ _06419_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_218_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29823_ clknet_leaf_307_clock _02836_ VGND VGND VPWR VPWR decode.regfile.registers_18\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_22158_ _06740_ _06742_ _06746_ _06752_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21109_ _09955_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_112_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_112_clock
+ sky130_fd_sc_hd__clkbuf_8
X_29754_ clknet_leaf_310_clock _02767_ VGND VGND VPWR VPWR decode.regfile.registers_16\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_22089_ _00001_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__buf_4
X_14980_ _10948_ _10954_ _10997_ net433 _10999_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__o311a_1
X_26966_ _09838_ VGND VGND VPWR VPWR _09866_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28705_ clknet_leaf_173_clock _01718_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13931_ _10053_ _10210_ VGND VGND VPWR VPWR _10218_ sky130_fd_sc_hd__nand2_1
X_25917_ net2469 _09242_ _09248_ _09235_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__o211a_1
X_29685_ clknet_leaf_282_clock _02698_ VGND VGND VPWR VPWR decode.regfile.registers_13\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_26897_ net1953 _09822_ _09826_ _09825_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28636_ clknet_leaf_182_clock _01649_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_16650_ _12614_ VGND VGND VPWR VPWR _12615_ sky130_fd_sc_hd__buf_4
X_13862_ _10152_ VGND VGND VPWR VPWR _10177_ sky130_fd_sc_hd__buf_2
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25848_ _09128_ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_127_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_127_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_18_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15601_ _11046_ decode.regfile.registers_12\[7\] _10649_ _11052_ _10632_ VGND VGND
+ VPWR VPWR _11591_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_97_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28567_ clknet_leaf_193_clock _01580_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16581_ _11024_ VGND VGND VPWR VPWR _12546_ sky130_fd_sc_hd__clkbuf_4
X_25779_ net619 _09156_ _09168_ _09169_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__o211a_1
X_13793_ _09954_ VGND VGND VPWR VPWR _10130_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18320_ _03625_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15532_ _11250_ decode.regfile.registers_27\[5\] _11258_ VGND VGND VPWR VPWR _11524_
+ sky130_fd_sc_hd__or3_1
X_27518_ clknet_leaf_21_clock _00547_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28498_ clknet_leaf_168_clock _01511_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18251_ _03584_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__clkbuf_1
X_27449_ clknet_leaf_159_clock _00478_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15463_ _11271_ VGND VGND VPWR VPWR _11456_ sky130_fd_sc_hd__buf_2
XFILLER_0_56_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17202_ _12658_ _13154_ _13155_ _13156_ VGND VGND VPWR VPWR _13157_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14414_ net610 _10490_ _10497_ _10494_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__o211a_1
X_18182_ decode.immGen._imm_T_10\[3\] _03519_ _03520_ _10581_ _11004_ VGND VGND VPWR
+ VPWR _00508_ sky130_fd_sc_hd__o311a_1
XFILLER_0_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15394_ decode.regfile.registers_18\[2\] _11268_ _11271_ _11388_ VGND VGND VPWR VPWR
+ _11389_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29119_ clknet_leaf_68_clock net1889 VGND VGND VPWR VPWR csr.mcycle\[3\] sky130_fd_sc_hd__dfxtp_2
X_17133_ _12695_ _13085_ _13086_ _13089_ VGND VGND VPWR VPWR _13090_ sky130_fd_sc_hd__a31o_1
X_14345_ net836 _10447_ _10457_ _10453_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold609 decode.regfile.registers_29\[28\] VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__dlygate4sd3_1
X_17064_ _13018_ _13019_ _13021_ _12889_ VGND VGND VPWR VPWR _13022_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14276_ net332 _10195_ _09933_ _10240_ VGND VGND VPWR VPWR _10417_ sky130_fd_sc_hd__and4_1
XFILLER_0_204_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16015_ decode.regfile.registers_3\[18\] _11292_ _11367_ _10635_ VGND VGND VPWR VPWR
+ _11994_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17966_ decode.regfile.registers_23\[29\] _12714_ _03337_ _03363_ _12514_ VGND VGND
+ VPWR VPWR _03364_ sky130_fd_sc_hd__o221a_1
XFILLER_0_178_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1309 decode.regfile.registers_8\[0\] VGND VGND VPWR VPWR net1536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16917_ _12791_ VGND VGND VPWR VPWR _12878_ sky130_fd_sc_hd__buf_4
X_19705_ _03893_ _03888_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__and2b_1
XFILLER_0_205_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17897_ _02990_ _03068_ decode.regfile.registers_27\[27\] _13487_ VGND VGND VPWR
+ VPWR _03297_ sky130_fd_sc_hd__or4_1
XFILLER_0_192_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16848_ _12512_ VGND VGND VPWR VPWR _12811_ sky130_fd_sc_hd__clkbuf_2
X_19636_ _03633_ _03635_ _03634_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__nor4_1
XFILLER_0_215_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_195_Right_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19567_ _04281_ _04283_ _04734_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__o21ai_1
X_16779_ decode.regfile.registers_10\[1\] _12599_ _12741_ _12742_ VGND VGND VPWR VPWR
+ _12743_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18518_ _03816_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19498_ _04186_ _04782_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_91_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_91_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_174_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18449_ decode.id_ex_ex_use_rs2_reg execute.io_mem_regwrite VGND VGND VPWR VPWR _03748_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_185_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21460_ _06151_ net1515 _06241_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20411_ _05570_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21391_ _06208_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23130_ _07368_ _07566_ _05246_ _07569_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_77_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20342_ _10854_ decode.id_ex_pc_reg\[28\] _10697_ _05500_ VGND VGND VPWR VPWR _05508_
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_71_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23061_ net68 _06718_ _07472_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20273_ _10694_ _05452_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_73_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22012_ csr.mscratch\[28\] _06601_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2500 decode.regfile.registers_2\[22\] VGND VGND VPWR VPWR net2727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2511 decode.regfile.registers_2\[18\] VGND VGND VPWR VPWR net2738 sky130_fd_sc_hd__dlygate4sd3_1
X_26820_ _09424_ _09776_ VGND VGND VPWR VPWR _09782_ sky130_fd_sc_hd__nand2_1
Xhold2522 csr.minstret\[12\] VGND VGND VPWR VPWR net2749 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2533 fetch.btb.btbTable\[11\]\[1\] VGND VGND VPWR VPWR net2760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2544 decode.io_id_pc\[16\] VGND VGND VPWR VPWR net2771 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1810 decode.regfile.registers_17\[27\] VGND VGND VPWR VPWR net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2555 decode.regfile.registers_30\[25\] VGND VGND VPWR VPWR net2782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2566 net72 VGND VGND VPWR VPWR net2793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1821 decode.regfile.registers_1\[14\] VGND VGND VPWR VPWR net2048 sky130_fd_sc_hd__dlygate4sd3_1
X_26751_ _09430_ _09733_ VGND VGND VPWR VPWR _09742_ sky130_fd_sc_hd__nand2_1
Xhold1832 fetch.bht.bhtTable_target_pc\[7\]\[25\] VGND VGND VPWR VPWR net2059 sky130_fd_sc_hd__dlygate4sd3_1
X_23963_ net1143 execute.io_target_pc\[3\] _07983_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_44_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_44_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_32_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1843 decode.regfile.registers_18\[31\] VGND VGND VPWR VPWR net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1854 decode.regfile.registers_6\[23\] VGND VGND VPWR VPWR net2081 sky130_fd_sc_hd__dlygate4sd3_1
X_25702_ net804 _09111_ _09124_ _09115_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__o211a_1
Xhold1865 fetch.bht.bhtTable_target_pc\[10\]\[30\] VGND VGND VPWR VPWR net2092 sky130_fd_sc_hd__dlygate4sd3_1
X_22914_ _06888_ _07007_ _07363_ _07364_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__and4bb_1
X_29470_ clknet_leaf_250_clock _02483_ VGND VGND VPWR VPWR decode.regfile.registers_7\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1876 decode.io_id_pc\[26\] VGND VGND VPWR VPWR net2103 sky130_fd_sc_hd__dlygate4sd3_1
X_26682_ net2037 _09692_ _09700_ _09702_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__o211a_1
Xhold1887 fetch.bht.bhtTable_target_pc\[10\]\[24\] VGND VGND VPWR VPWR net2114 sky130_fd_sc_hd__dlygate4sd3_1
X_23894_ _08116_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__clkbuf_1
Xhold1898 fetch.bht.bhtTable_tag\[2\]\[20\] VGND VGND VPWR VPWR net2125 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28421_ clknet_leaf_39_clock _01434_ VGND VGND VPWR VPWR decode.immGen._imm_T_10\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25633_ _08933_ _09079_ VGND VGND VPWR VPWR _09085_ sky130_fd_sc_hd__nand2_1
X_22845_ _07318_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28352_ clknet_leaf_189_clock _01365_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_59_clock
+ sky130_fd_sc_hd__clkbuf_8
X_25564_ _08939_ _09036_ VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22776_ _07281_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27303_ clknet_leaf_13_clock _00332_ VGND VGND VPWR VPWR decode.regfile.registers_31\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24515_ _08438_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28283_ clknet_leaf_85_clock _01305_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_21727_ csr.mtie csr.ie csr.mtip _06423_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__a31o_1
X_25495_ _08978_ VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27234_ clknet_leaf_364_clock _00263_ VGND VGND VPWR VPWR decode.regfile.registers_29\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_24446_ _08402_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__clkbuf_1
X_21658_ _05691_ csr.minstret\[16\] csr.io_inst_retired _06363_ VGND VGND VPWR VPWR
+ _06370_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_62_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20609_ _05672_ _05741_ _05743_ _05745_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__a31o_1
X_27165_ clknet_leaf_359_clock _00194_ VGND VGND VPWR VPWR decode.regfile.registers_27\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_24377_ _08365_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__clkbuf_1
X_21589_ _10576_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14130_ net732 _10332_ _10334_ _10328_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__o211a_1
X_26116_ _08962_ _09353_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__nand2_1
X_23328_ _07755_ _07071_ _07080_ VGND VGND VPWR VPWR _07756_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27096_ clknet_leaf_354_clock _00125_ VGND VGND VPWR VPWR decode.regfile.registers_25\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14061_ net710 _10287_ _10294_ _10291_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__o211a_1
X_26047_ _08968_ _09285_ VGND VGND VPWR VPWR _09323_ sky130_fd_sc_hd__nand2_1
X_23259_ fetch.bht.bhtTable_target_pc\[0\]\[21\] fetch.bht.bhtTable_target_pc\[1\]\[21\]
+ fetch.bht.bhtTable_target_pc\[2\]\[21\] fetch.bht.bhtTable_target_pc\[3\]\[21\]
+ _07119_ _07071_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17820_ _10929_ decode.regfile.registers_28\[25\] _02992_ VGND VGND VPWR VPWR _03222_
+ sky130_fd_sc_hd__o21a_1
X_29806_ clknet_leaf_295_clock _02819_ VGND VGND VPWR VPWR decode.regfile.registers_17\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_27998_ clknet_leaf_204_clock _01020_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_17751_ decode.regfile.registers_1\[24\] net215 _12530_ VGND VGND VPWR VPWR _03154_
+ sky130_fd_sc_hd__and3_1
X_29737_ clknet_leaf_293_clock _02750_ VGND VGND VPWR VPWR decode.regfile.registers_15\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_26949_ net1663 _09853_ _09856_ _09852_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__o211a_1
X_14963_ _10651_ VGND VGND VPWR VPWR _10988_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16702_ _12666_ VGND VGND VPWR VPWR _12667_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13914_ net726 _10199_ _10208_ _10206_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29668_ clknet_leaf_277_clock _02681_ VGND VGND VPWR VPWR decode.regfile.registers_13\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_17682_ decode.regfile.registers_9\[22\] _11017_ _12502_ _12509_ _12652_ VGND VGND
+ VPWR VPWR _03087_ sky130_fd_sc_hd__o41a_1
XFILLER_0_215_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14894_ _10930_ VGND VGND VPWR VPWR _10931_ sky130_fd_sc_hd__buf_4
XFILLER_0_18_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19421_ _04359_ _04703_ _04391_ _04708_ _04392_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__a32o_1
XFILLER_0_226_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28619_ clknet_leaf_95_clock _01632_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16633_ _10609_ _12592_ _12597_ VGND VGND VPWR VPWR _12598_ sky130_fd_sc_hd__and3_2
X_13845_ _10031_ _10164_ VGND VGND VPWR VPWR _10168_ sky130_fd_sc_hd__nand2_1
X_29599_ clknet_leaf_270_clock _02612_ VGND VGND VPWR VPWR decode.regfile.registers_11\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1087 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19352_ _04638_ _04639_ _04641_ _04642_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__a22o_1
X_16564_ decode.immGen._imm_T_24\[16\] decode.immGen._imm_T_24\[15\] VGND VGND VPWR
+ VPWR _12529_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13776_ memory.io_wb_reg_pc\[26\] _09946_ _09947_ _10114_ VGND VGND VPWR VPWR _10115_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18303_ decode.id_ex_rs2_data_reg\[17\] _03616_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15515_ decode.regfile.registers_8\[5\] _11284_ _11287_ decode.regfile.registers_9\[5\]
+ _11131_ VGND VGND VPWR VPWR _11507_ sky130_fd_sc_hd__o221a_1
X_19283_ _04294_ _04571_ _04576_ _04514_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16495_ _12459_ _12460_ VGND VGND VPWR VPWR _12461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_216_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18234_ csr._mcycle_T_3\[53\] csr._mcycle_T_3\[52\] csr._mcycle_T_3\[51\] csr._mcycle_T_3\[50\]
+ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15446_ _11347_ VGND VGND VPWR VPWR _11440_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18165_ _03510_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15377_ decode.regfile.registers_1\[2\] _11371_ VGND VGND VPWR VPWR _11372_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17116_ _11021_ _12567_ _12586_ _12673_ decode.regfile.registers_16\[8\] VGND VGND
+ VPWR VPWR _13073_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14328_ net880 _10447_ _10448_ _10440_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__o211a_1
X_18096_ _10915_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__clkbuf_2
Xhold406 decode.regfile.registers_7\[9\] VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold417 decode.regfile.registers_17\[14\] VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold428 decode.regfile.registers_14\[7\] VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 decode.regfile.registers_28\[30\] VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17047_ decode.regfile.registers_29\[6\] _12965_ _12966_ _13005_ _12702_ VGND VGND
+ VPWR VPWR _13006_ sky130_fd_sc_hd__o221a_1
XFILLER_0_96_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14259_ _10107_ _10400_ VGND VGND VPWR VPWR _10408_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18998_ _03709_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__buf_4
Xhold1106 fetch.bht.bhtTable_tag\[9\]\[12\] VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 decode.regfile.registers_6\[1\] VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1128 fetch.bht.bhtTable_target_pc\[13\]\[31\] VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17949_ _12880_ _03346_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1139 decode.regfile.registers_25\[6\] VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20960_ execute.io_reg_pc\[6\] _05915_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__and3_1
XFILLER_0_224_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_176_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19619_ _04427_ _04879_ _04290_ _04541_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__and4b_1
X_20891_ _05924_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22630_ net2140 _07196_ _07179_ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_221_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22561_ _10576_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__buf_4
XFILLER_0_36_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_370 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24300_ _08062_ net2035 _08323_ VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__mux2_1
XINSDIODE1_381 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21512_ _06273_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22492_ _06720_ _06769_ _06822_ _07062_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__or4_4
X_25280_ _08870_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_135_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21443_ _06134_ net1568 _06230_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__mux2_1
X_24231_ _08290_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24162_ _08254_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_131_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21374_ _06122_ net2079 _06199_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23113_ _07347_ _07538_ _07553_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__or3_1
XFILLER_0_142_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20325_ _05420_ _05373_ _05495_ _05454_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_9_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28970_ clknet_leaf_98_clock _01983_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_24093_ net1174 execute.io_target_pc\[2\] _06450_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold940 decode.regfile.registers_13\[15\] VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 fetch.bht.bhtTable_tag\[3\]\[13\] VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold962 fetch.bht.bhtTable_target_pc\[8\]\[22\] VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__dlygate4sd3_1
X_23044_ csr._csr_read_data_T_8\[9\] _06039_ csr.io_mret_vector\[9\] _06463_ VGND
+ VGND VPWR VPWR _07488_ sky130_fd_sc_hd__a22o_1
X_27921_ clknet_leaf_70_clock _00950_ VGND VGND VPWR VPWR csr.io_csr_write_address\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold973 fetch.bht.bhtTable_tag\[8\]\[19\] VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__dlygate4sd3_1
X_20256_ _05441_ _05442_ _05277_ _05411_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__a22o_1
XFILLER_0_229_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold984 fetch.bht.bhtTable_target_pc\[15\]\[22\] VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 decode.regfile.registers_21\[17\] VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_30__f_clock clknet_2_3_0_clock VGND VGND VPWR VPWR clknet_5_30__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_27852_ clknet_leaf_321_clock _00881_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20187_ _05385_ _05386_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2330 decode.regfile.registers_27\[14\] VGND VGND VPWR VPWR net2557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2341 csr._csr_read_data_T_8\[10\] VGND VGND VPWR VPWR net2568 sky130_fd_sc_hd__dlygate4sd3_1
X_26803_ net2539 _09766_ _09772_ _09771_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__o211a_1
Xhold2352 decode.regfile.registers_6\[26\] VGND VGND VPWR VPWR net2579 sky130_fd_sc_hd__dlygate4sd3_1
X_27783_ clknet_leaf_324_clock _00812_ VGND VGND VPWR VPWR memory.io_wb_readdata\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24995_ _08703_ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__clkbuf_4
Xhold2363 csr._minstret_T_3\[33\] VGND VGND VPWR VPWR net2590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2374 decode.regfile.registers_2\[19\] VGND VGND VPWR VPWR net2601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1640 fetch.bht.bhtTable_target_pc\[6\]\[2\] VGND VGND VPWR VPWR net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2385 fetch.btb.btbTable\[8\]\[1\] VGND VGND VPWR VPWR net2612 sky130_fd_sc_hd__dlygate4sd3_1
X_29522_ clknet_leaf_265_clock _02535_ VGND VGND VPWR VPWR decode.regfile.registers_8\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1651 fetch.bht.bhtTable_tag\[7\]\[14\] VGND VGND VPWR VPWR net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2396 fetch.btb.btbTable\[6\]\[1\] VGND VGND VPWR VPWR net2623 sky130_fd_sc_hd__dlygate4sd3_1
X_26734_ net1767 _09723_ _09732_ _09730_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__o211a_1
X_23946_ _08143_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__clkbuf_1
Xhold1662 _02132_ VGND VGND VPWR VPWR net1889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1673 fetch.bht.bhtTable_tag\[14\]\[2\] VGND VGND VPWR VPWR net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1684 csr.mcycle\[25\] VGND VGND VPWR VPWR net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1695 fetch.bht.bhtTable_tag\[15\]\[6\] VGND VGND VPWR VPWR net1922 sky130_fd_sc_hd__dlygate4sd3_1
X_29453_ clknet_leaf_261_clock _02466_ VGND VGND VPWR VPWR decode.regfile.registers_6\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_26665_ _09420_ _09689_ VGND VGND VPWR VPWR _09693_ sky130_fd_sc_hd__nand2_1
X_23877_ _08105_ net1560 _07940_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__mux2_1
X_28404_ clknet_leaf_142_clock _01417_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13630_ _09943_ memory.io_wb_aluresult\[5\] _09980_ memory.io_wb_readdata\[5\] VGND
+ VGND VPWR VPWR _09990_ sky130_fd_sc_hd__a22o_1
X_25616_ net772 _09068_ _09075_ _09074_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__o211a_1
X_22828_ net1259 _10759_ _07308_ VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29384_ clknet_leaf_258_clock _02397_ VGND VGND VPWR VPWR decode.regfile.registers_4\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_26596_ _09426_ _09645_ VGND VGND VPWR VPWR _09653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28335_ clknet_leaf_222_clock _01348_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13561_ _09927_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
X_25547_ net1300 _09024_ _09035_ _09033_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__o211a_1
X_22759_ _07272_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15300_ _11295_ VGND VGND VPWR VPWR _11296_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28266_ clknet_leaf_61_clock _01288_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16280_ _11174_ _12249_ _12250_ _12251_ VGND VGND VPWR VPWR _12252_ sky130_fd_sc_hd__a31o_1
X_25478_ _08929_ _08992_ VGND VGND VPWR VPWR _08996_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_229_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15231_ _11227_ VGND VGND VPWR VPWR _11228_ sky130_fd_sc_hd__buf_2
X_27217_ clknet_leaf_329_clock _00246_ VGND VGND VPWR VPWR decode.regfile.registers_29\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24429_ _08393_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28197_ clknet_leaf_60_clock _01219_ VGND VGND VPWR VPWR csr.io_mret_vector\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15162_ _11154_ decode.regfile.registers_0\[0\] _11156_ _11158_ VGND VGND VPWR VPWR
+ _11159_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27148_ clknet_leaf_359_clock _00177_ VGND VGND VPWR VPWR decode.regfile.registers_26\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14113_ net2510 _10315_ _10323_ _10317_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__o211a_1
X_19970_ _10710_ _05214_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__and2_1
X_27079_ clknet_leaf_347_clock _00108_ VGND VGND VPWR VPWR decode.regfile.registers_24\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15093_ _11089_ VGND VGND VPWR VPWR _11090_ sky130_fd_sc_hd__clkbuf_4
X_14044_ _10142_ _10242_ VGND VGND VPWR VPWR _10283_ sky130_fd_sc_hd__nand2_1
X_18921_ _03795_ _03800_ _04218_ _04219_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__a211o_1
XFILLER_0_197_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18852_ decode.id_ex_rs2_data_reg\[11\] net199 _04145_ net259 _04150_ VGND VGND VPWR
+ VPWR _04151_ sky130_fd_sc_hd__o221a_1
XFILLER_0_197_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17803_ decode.regfile.registers_13\[25\] _12775_ _03203_ _03204_ _12664_ VGND VGND
+ VPWR VPWR _03205_ sky130_fd_sc_hd__a221oi_2
X_18783_ _03796_ _04079_ _03889_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__a21oi_1
X_15995_ decode.regfile.registers_23\[17\] _11262_ _11946_ _11974_ _11336_ VGND VGND
+ VPWR VPWR _11975_ sky130_fd_sc_hd__o221a_1
XFILLER_0_101_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17734_ _13250_ decode.regfile.registers_24\[23\] _12997_ _12998_ _13367_ VGND VGND
+ VPWR VPWR _03138_ sky130_fd_sc_hd__o2111a_1
X_14946_ _10963_ _10966_ _10974_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_216_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17665_ _13221_ _03067_ _03069_ _03070_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14877_ _10912_ _10913_ _10916_ decode.immGen._imm_T_10\[1\] VGND VGND VPWR VPWR
+ _10918_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_106_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_218_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1090 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19404_ _04291_ _04692_ _04646_ _04427_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__o2bb2a_1
X_16616_ _10593_ _10598_ decode.immGen._imm_T_24\[17\] VGND VGND VPWR VPWR _12581_
+ sky130_fd_sc_hd__and3_1
X_13828_ _09975_ _10154_ VGND VGND VPWR VPWR _10158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17596_ _12830_ _03001_ _03002_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_214_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19335_ _04469_ _04472_ net242 VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__mux2_2
X_16547_ _12511_ VGND VGND VPWR VPWR _12512_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13759_ memory.csr_read_data_out_reg\[23\] _09986_ _10099_ _10100_ VGND VGND VPWR
+ VPWR _10101_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_174_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19266_ _04052_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16478_ _10958_ decode.regfile.registers_26\[30\] _11676_ _11338_ _10992_ VGND VGND
+ VPWR VPWR _12445_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_72_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18217_ net2783 _10998_ _03552_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__and3_1
X_15429_ decode.regfile.registers_15\[3\] _11036_ _11204_ _11361_ VGND VGND VPWR VPWR
+ _11423_ sky130_fd_sc_hd__a31o_1
XFILLER_0_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19197_ _04022_ _04451_ _04448_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18148_ _03503_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold203 decode.regfile.registers_30\[13\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold214 decode.regfile.registers_31\[9\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_TAPCELL_ROW_169_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18079_ _10575_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__buf_2
XFILLER_0_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold225 decode.regfile.registers_25\[9\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold236 decode.regfile.registers_31\[26\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__buf_1
Xhold247 decode.exception_out_reg VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
X_20110_ _05319_ _05320_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__and2b_1
Xhold258 decode.regfile.registers_31\[23\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_165_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold269 decode.regfile.registers_30\[26\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__buf_1
X_21090_ _10576_ _06032_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_165_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20041_ _05260_ _05261_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_13_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23800_ _08053_ net1708 _07952_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24780_ _08576_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__clkbuf_1
X_21992_ csr._mcycle_T_2\[19\] _06587_ _06599_ _06592_ VGND VGND VPWR VPWR _01239_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_124_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23731_ net1340 _10771_ _08014_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__mux2_1
XANTENNA_109 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20943_ _05949_ _05945_ net57 VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_221_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26450_ _09430_ _09558_ VGND VGND VPWR VPWR _09569_ sky130_fd_sc_hd__nand2_1
X_23662_ _07979_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20874_ _05866_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__clkbuf_2
X_25401_ _08943_ _08923_ VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22613_ net2156 _07185_ _07179_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__a21oi_1
X_26381_ net1212 _09518_ _09528_ _09525_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__o211a_1
X_23593_ _07942_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28120_ clknet_leaf_89_clock _01142_ VGND VGND VPWR VPWR csr.minstret\[25\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_165_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25332_ _08891_ net2698 VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__and2_1
X_22544_ csr._minstret_T_3\[32\] csr.minstret\[31\] _06420_ _06422_ VGND VGND VPWR
+ VPWR _07137_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28051_ clknet_leaf_206_clock _01073_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25263_ _08861_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__clkbuf_1
X_22475_ _06661_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27002_ clknet_leaf_337_clock _00031_ VGND VGND VPWR VPWR decode.regfile.registers_22\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24214_ _08281_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__clkbuf_1
X_21426_ _06117_ net846 _06219_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__mux2_1
X_25194_ _09880_ _09883_ _08808_ VGND VGND VPWR VPWR _08826_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24145_ net810 execute.io_target_pc\[27\] _06427_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__mux2_1
X_21357_ _06105_ net2205 _06188_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20308_ _05340_ _10867_ _10798_ _05473_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_57_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28953_ clknet_leaf_128_clock _01966_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_24076_ _08210_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__clkbuf_1
X_21288_ net1881 _06151_ _06141_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold770 _08368_ VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold781 fetch.bht.bhtTable_target_pc\[12\]\[1\] VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 fetch.bht.bhtTable_tag\[11\]\[7\] VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27904_ clknet_leaf_81_clock _00933_ VGND VGND VPWR VPWR csr._mcycle_T_2\[25\] sky130_fd_sc_hd__dfxtp_1
X_23027_ net97 net96 net227 _07427_ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__and4_2
X_20239_ _05412_ _05253_ _05429_ _03517_ _03551_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_124_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28884_ clknet_leaf_118_clock _01897_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27835_ clknet_leaf_325_clock _00864_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2160 decode.regfile.registers_16\[10\] VGND VGND VPWR VPWR net2387 sky130_fd_sc_hd__dlygate4sd3_1
X_14800_ _10706_ net270 _10818_ _10819_ _10842_ VGND VGND VPWR VPWR _10843_ sky130_fd_sc_hd__o311a_1
Xhold2171 decode.regfile.registers_2\[3\] VGND VGND VPWR VPWR net2398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2182 decode.regfile.registers_17\[30\] VGND VGND VPWR VPWR net2409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15780_ decode.regfile.registers_10\[12\] _11382_ VGND VGND VPWR VPWR _11765_ sky130_fd_sc_hd__nor2_1
X_27766_ clknet_leaf_321_clock _00795_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_24978_ net2548 _08696_ net791 VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__a21oi_1
Xhold2193 decode.regfile.registers_27\[22\] VGND VGND VPWR VPWR net2420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1470 decode.regfile.registers_12\[17\] VGND VGND VPWR VPWR net1697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1481 fetch.bht.bhtTable_target_pc\[15\]\[2\] VGND VGND VPWR VPWR net1708 sky130_fd_sc_hd__dlygate4sd3_1
X_14731_ csr.io_mem_pc\[26\] csr.io_mem_pc\[27\] _10768_ VGND VGND VPWR VPWR _10774_
+ sky130_fd_sc_hd__and3_1
X_26717_ _09708_ VGND VGND VPWR VPWR _09723_ sky130_fd_sc_hd__clkbuf_4
X_29505_ clknet_leaf_250_clock _02518_ VGND VGND VPWR VPWR decode.regfile.registers_8\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_23929_ net1028 _08087_ _08130_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__mux2_1
Xhold1492 decode.regfile.registers_22\[17\] VGND VGND VPWR VPWR net1719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27697_ clknet_leaf_24_clock _00726_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17450_ decode.regfile.registers_17\[16\] _12579_ _13379_ _13398_ _12565_ VGND VGND
+ VPWR VPWR _13399_ sky130_fd_sc_hd__o221a_1
X_29436_ clknet_leaf_248_clock _02449_ VGND VGND VPWR VPWR decode.regfile.registers_6\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14662_ _10704_ VGND VGND VPWR VPWR _10705_ sky130_fd_sc_hd__inv_2
X_26648_ _09402_ _09676_ VGND VGND VPWR VPWR _09683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16401_ decode.regfile.registers_20\[28\] _11452_ _11223_ _12369_ VGND VGND VPWR
+ VPWR _12370_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_40_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13613_ net210 VGND VGND VPWR VPWR _09975_ sky130_fd_sc_hd__clkbuf_4
X_29367_ clknet_leaf_258_clock _02380_ VGND VGND VPWR VPWR decode.regfile.registers_3\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_17381_ decode.regfile.registers_24\[14\] _12691_ _13304_ _13331_ VGND VGND VPWR
+ VPWR _13332_ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14593_ _10635_ VGND VGND VPWR VPWR _10636_ sky130_fd_sc_hd__clkbuf_4
X_26579_ _09408_ _09632_ VGND VGND VPWR VPWR _09643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19120_ _04248_ _04257_ _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__o21ba_1
X_28318_ clknet_leaf_209_clock _01331_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_16332_ decode.regfile.registers_25\[26\] _11333_ _11336_ decode.regfile.registers_24\[26\]
+ VGND VGND VPWR VPWR _12303_ sky130_fd_sc_hd__o22a_1
XFILLER_0_229_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13544_ _09914_ _09890_ _09916_ net400 VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29298_ clknet_leaf_225_clock _02311_ VGND VGND VPWR VPWR decode.regfile.registers_1\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19051_ _04290_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__clkbuf_4
X_28249_ clknet_leaf_79_clock _01271_ VGND VGND VPWR VPWR csr._minstret_T_3\[49\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16263_ _11646_ _11834_ _11944_ decode.regfile.registers_29\[24\] _12235_ VGND VGND
+ VPWR VPWR _12236_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18002_ decode.regfile.registers_22\[30\] _13100_ _03398_ _13289_ VGND VGND VPWR
+ VPWR _03399_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15214_ _11124_ decode.regfile.registers_16\[0\] _11128_ _11210_ VGND VGND VPWR VPWR
+ _11211_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_11_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16194_ _12133_ net436 _12134_ _12168_ _12132_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__o221a_1
XFILLER_0_164_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15145_ _11141_ VGND VGND VPWR VPWR _11142_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19953_ decode.id_ex_pc_reg\[1\] _03627_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__and2_1
X_15076_ _10989_ _11072_ _11065_ VGND VGND VPWR VPWR _11073_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_207_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_207_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_207_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14027_ _10097_ _10268_ VGND VGND VPWR VPWR _10274_ sky130_fd_sc_hd__nand2_1
X_18904_ _03890_ decode.id_ex_imm_reg\[19\] _03898_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__a21oi_1
X_19884_ _03789_ _03790_ _05153_ _04465_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__o31a_1
XFILLER_0_219_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18835_ _03658_ execute.csr_read_data_out_reg\[9\] execute.io_reg_pc\[9\] _03662_
+ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_199_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15978_ _11367_ _11952_ _11953_ _11957_ VGND VGND VPWR VPWR _11958_ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18766_ _03708_ decode.id_ex_imm_reg\[7\] _04064_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_179_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17717_ decode.regfile.registers_2\[23\] _12634_ _12628_ _03120_ VGND VGND VPWR VPWR
+ _03121_ sky130_fd_sc_hd__o211a_1
X_14929_ _10957_ VGND VGND VPWR VPWR _10958_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18697_ net326 _03995_ net250 net359 decode.id_ex_immsrc_reg VGND VGND VPWR VPWR
+ _03996_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17648_ decode.regfile.registers_16\[21\] _13011_ _03033_ _03053_ VGND VGND VPWR
+ VPWR _03054_ sky130_fd_sc_hd__o22a_1
XFILLER_0_202_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17579_ _11026_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19318_ _04609_ _04345_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20590_ _05726_ _05729_ _05630_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__o21a_2
XFILLER_0_2_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19249_ _04337_ _04436_ _04329_ _04305_ _04543_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22260_ _06790_ _06850_ _06852_ _06854_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__o22a_1
XFILLER_0_171_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21211_ decode.id_ex_ex_rd_reg\[4\] _05214_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__and2_1
XFILLER_0_143_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22191_ fetch.bht.bhtTable_tag\[0\]\[5\] fetch.bht.bhtTable_tag\[1\]\[5\] fetch.bht.bhtTable_tag\[2\]\[5\]
+ fetch.bht.bhtTable_tag\[3\]\[5\] _06700_ _06685_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21142_ _06064_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4 _06313_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__buf_2
X_25950_ _08945_ _09267_ VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__nand2_1
X_21073_ execute.csr_read_data_out_reg\[25\] _06014_ _03583_ VGND VGND VPWR VPWR _06023_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20024_ _10575_ _05222_ _05246_ _10908_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__or4_4
X_24901_ net581 _08647_ _08648_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_126_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25881_ _08954_ _09223_ VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__nand2_1
X_27620_ clknet_leaf_147_clock _00649_ VGND VGND VPWR VPWR execute.io_target_pc\[29\]
+ sky130_fd_sc_hd__dfxtp_4
X_24832_ _08603_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27551_ clknet_leaf_38_clock _00580_ VGND VGND VPWR VPWR execute.io_mem_zero sky130_fd_sc_hd__dfxtp_1
X_24763_ _08567_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21975_ csr._mcycle_T_2\[11\] _06587_ _06590_ _06579_ VGND VGND VPWR VPWR _01231_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer40 net272 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26502_ _09406_ _09589_ VGND VGND VPWR VPWR _09599_ sky130_fd_sc_hd__nand2_1
Xrebuffer51 _04152_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__buf_1
XFILLER_0_222_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23714_ net932 _10795_ _08003_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__mux2_1
Xrebuffer62 net288 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer73 net302 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20926_ _05943_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__clkbuf_1
X_27482_ clknet_leaf_38_clock _00511_ VGND VGND VPWR VPWR decode.io_mret_out sky130_fd_sc_hd__dfxtp_1
X_24694_ _08530_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer84 net309 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_1
X_29221_ clknet_leaf_102_clock _02234_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer95 net321 VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26433_ _09412_ _09558_ VGND VGND VPWR VPWR _09559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23645_ _07970_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__clkbuf_1
X_20857_ net115 _05903_ _05899_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29152_ clknet_leaf_222_clock _02165_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26364_ net2307 _09518_ _09519_ _09512_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__o211a_1
X_23576_ _06107_ net1664 _07930_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20788_ _09955_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__clkbuf_4
X_28103_ clknet_leaf_74_clock net2437 VGND VGND VPWR VPWR csr.minstret\[8\] sky130_fd_sc_hd__dfxtp_1
X_25315_ _08880_ net2680 VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29083_ clknet_leaf_184_clock _02096_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_22527_ _07072_ _07120_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26295_ net2375 _09475_ _09479_ _09471_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28034_ clknet_leaf_168_clock _01056_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_25246_ _08085_ net1640 _08848_ VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22458_ _06616_ fetch.btb.btbTable\[4\]\[1\] fetch.bht.bhtTable_valid\[4\] VGND VGND
+ VPWR VPWR _07053_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_59_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21409_ _06218_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__clkbuf_8
X_25177_ _08817_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22389_ fetch.bht.bhtTable_tag\[8\]\[9\] fetch.bht.bhtTable_tag\[9\]\[9\] fetch.bht.bhtTable_tag\[10\]\[9\]
+ fetch.bht.bhtTable_tag\[11\]\[9\] _06754_ _06675_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_55_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24128_ net968 VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28936_ clknet_leaf_100_clock _01949_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24059_ net856 execute.io_target_pc\[17\] _08198_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__mux2_1
X_16950_ decode.regfile.registers_22\[4\] _12527_ _12908_ _12910_ _12686_ VGND VGND
+ VPWR VPWR _12911_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15901_ decode.regfile.registers_1\[15\] _11539_ _11882_ VGND VGND VPWR VPWR _11883_
+ sky130_fd_sc_hd__a21o_1
X_16881_ _12842_ VGND VGND VPWR VPWR _12843_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_218_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_216_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28867_ clknet_leaf_125_clock _01880_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_202_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15832_ decode.regfile.registers_13\[13\] _11046_ _11689_ _11318_ _11052_ VGND VGND
+ VPWR VPWR _11816_ sky130_fd_sc_hd__o32a_1
X_18620_ _03751_ net325 _03757_ net267 decode.id_ex_rs2_data_reg\[18\] VGND VGND VPWR
+ VPWR _03919_ sky130_fd_sc_hd__a311o_4
XFILLER_0_189_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27818_ clknet_leaf_321_clock _00847_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_28798_ clknet_leaf_176_clock _01811_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_194_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ decode.regfile.registers_21\[11\] _11222_ _11096_ _11748_ VGND VGND VPWR
+ VPWR _11749_ sky130_fd_sc_hd__a211o_1
X_18551_ _03848_ _03849_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__and2_1
XFILLER_0_220_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27749_ clknet_leaf_323_clock _00778_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_194_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _10756_ VGND VGND VPWR VPWR _10757_ sky130_fd_sc_hd__clkbuf_4
X_17502_ _13099_ _13262_ _13182_ decode.regfile.registers_29\[17\] _13449_ VGND VGND
+ VPWR VPWR _13450_ sky130_fd_sc_hd__o221a_1
XFILLER_0_197_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18482_ net194 _03772_ _03775_ _03780_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__a211oi_4
X_15694_ _10960_ decode.regfile.registers_28\[9\] _11067_ _11681_ _11440_ VGND VGND
+ VPWR VPWR _11682_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_190_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ decode.regfile.registers_1\[16\] VGND VGND VPWR VPWR _13382_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_190_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ execute.io_target_pc\[11\] VGND VGND VPWR VPWR _10688_ sky130_fd_sc_hd__inv_2
X_29419_ clknet_leaf_257_clock _02432_ VGND VGND VPWR VPWR decode.regfile.registers_5\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17364_ decode.regfile.registers_3\[14\] _12627_ _10608_ _12613_ VGND VGND VPWR VPWR
+ _13315_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_16_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14576_ _10618_ VGND VGND VPWR VPWR _10619_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19103_ decode.id_ex_aluop_reg\[1\] decode.id_ex_aluop_reg\[3\] decode.id_ex_aluop_reg\[2\]
+ _04299_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__or4_4
X_16315_ _11318_ _11085_ _12285_ VGND VGND VPWR VPWR _12286_ sky130_fd_sc_hd__o21ai_1
X_13527_ _09904_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17295_ decode.regfile.registers_22\[12\] _12528_ _13247_ _12687_ VGND VGND VPWR
+ VPWR _13248_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19034_ _04126_ _04137_ _04255_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__mux2_1
X_16246_ _11181_ _12217_ _12218_ VGND VGND VPWR VPWR _12219_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_209_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16177_ _11047_ decode.regfile.registers_12\[22\] _10650_ _11053_ _10632_ VGND VGND
+ VPWR VPWR _12152_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_24_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput105 net105 VGND VGND VPWR VPWR io_memory_address[14] sky130_fd_sc_hd__clkbuf_4
Xoutput116 net116 VGND VGND VPWR VPWR io_memory_address[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput127 net127 VGND VGND VPWR VPWR io_memory_address[5] sky130_fd_sc_hd__clkbuf_4
X_15128_ _11121_ VGND VGND VPWR VPWR _11125_ sky130_fd_sc_hd__buf_4
Xoutput138 net138 VGND VGND VPWR VPWR io_memory_write_data[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_220_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput149 net149 VGND VGND VPWR VPWR io_memory_write_data[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15059_ _11055_ VGND VGND VPWR VPWR _11056_ sky130_fd_sc_hd__buf_2
X_19936_ _03581_ _05201_ net466 VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__and3b_1
XFILLER_0_103_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19867_ net189 _04320_ net187 VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_207_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18818_ _04108_ _03914_ _03908_ decode.id_ex_rs1_data_reg\[12\] _04111_ VGND VGND
+ VPWR VPWR _04117_ sky130_fd_sc_hd__o221ai_4
X_19798_ _04297_ _04261_ _04263_ _05070_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_121_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18749_ _04042_ _04046_ _03746_ decode.id_ex_rs2_data_reg\[5\] _04047_ VGND VGND
+ VPWR VPWR _04048_ sky130_fd_sc_hd__o221a_1
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21760_ net815 _10800_ _06439_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20711_ _05801_ _05808_ decode.id_ex_rs1_data_reg\[14\] _05824_ _00701_ VGND VGND
+ VPWR VPWR _00733_ sky130_fd_sc_hd__a32o_1
XFILLER_0_187_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21691_ csr._mcycle_T_2\[26\] _06329_ csr.minstret\[26\] VGND VGND VPWR VPWR _06394_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23430_ _07849_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_1343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20642_ csr.mscratch\[28\] _05593_ _05625_ _05772_ _05773_ VGND VGND VPWR VPWR _05774_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23361_ csr._csr_read_data_T_8\[27\] _07416_ csr.io_mret_vector\[27\] _07621_ _07786_
+ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__o221a_1
X_20573_ csr.mscratch\[18\] _05592_ _05611_ _05713_ _05714_ VGND VGND VPWR VPWR _05715_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_116_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25100_ _08561_ VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__clkbuf_8
X_22312_ _06628_ _06900_ _06902_ _06906_ _06636_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_115_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26080_ net1607 _09329_ _09342_ _09333_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__o211a_1
X_23292_ fetch.bht.bhtTable_target_pc\[4\]\[23\] fetch.bht.bhtTable_target_pc\[5\]\[23\]
+ fetch.bht.bhtTable_target_pc\[6\]\[23\] fetch.bht.bhtTable_target_pc\[7\]\[23\]
+ _07708_ _07103_ VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25031_ csr._mcycle_T_2\[15\] _08712_ _08733_ csr.mcycle\[15\] VGND VGND VPWR VPWR
+ _08734_ sky130_fd_sc_hd__a211o_1
X_22243_ _06835_ _06678_ _06672_ _06837_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_48_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22174_ net68 _06739_ _06670_ net221 _06768_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_169_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21125_ _06050_ _06046_ net483 VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__and3_1
X_29770_ clknet_leaf_295_clock _02783_ VGND VGND VPWR VPWR decode.regfile.registers_16\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_26982_ net1993 _09866_ _09874_ _09865_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28721_ clknet_leaf_104_clock _01734_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_25933_ _08931_ _09253_ VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__nand2_1
X_21056_ _05864_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20007_ _04018_ _10711_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_214_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28652_ clknet_leaf_87_clock _01665_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25864_ _08937_ _09210_ VGND VGND VPWR VPWR _09218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_213_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_199_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24815_ _08594_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27603_ clknet_leaf_151_clock _00632_ VGND VGND VPWR VPWR execute.io_target_pc\[12\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_2_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28583_ clknet_leaf_111_clock _01596_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25795_ _08943_ _09166_ VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27534_ clknet_leaf_155_clock _00563_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_115_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24746_ _08557_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__clkbuf_1
X_21958_ net1569 _06574_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27465_ clknet_leaf_148_clock _00494_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[31\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_166_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20909_ _05934_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_1196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24677_ net1316 execute.io_target_pc\[27\] _07285_ VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ _06531_ _06519_ _06520_ _06532_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29204_ clknet_leaf_240_clock _02217_ VGND VGND VPWR VPWR fetch.btb.btbTable\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_26416_ net1265 _09548_ _09549_ _09540_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_13_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _10505_ VGND VGND VPWR VPWR _10507_ sky130_fd_sc_hd__clkbuf_4
X_23628_ net998 _10820_ _07961_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27396_ clknet_leaf_31_clock _00425_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29135_ clknet_leaf_78_clock _02148_ VGND VGND VPWR VPWR csr.mcycle\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26347_ net2131 _09505_ _09509_ _09499_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__o211a_1
X_14361_ _10426_ VGND VGND VPWR VPWR _10468_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_182_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23559_ net2122 _07918_ _07915_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__or3b_1
XFILLER_0_135_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_342_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_342_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 net386 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16100_ decode.regfile.registers_15\[20\] _11047_ _11199_ _11359_ VGND VGND VPWR
+ VPWR _12077_ sky130_fd_sc_hd__o31a_1
XFILLER_0_181_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29066_ clknet_leaf_208_clock _02079_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput29 net397 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
X_17080_ _12546_ _12554_ _12535_ _13037_ VGND VGND VPWR VPWR _13038_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26278_ net2615 _09462_ _09469_ _09458_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__o211a_1
X_14292_ _09993_ _10420_ VGND VGND VPWR VPWR _10428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28017_ clknet_leaf_234_clock _01039_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16031_ decode.regfile.registers_25\[18\] _11483_ _11484_ decode.regfile.registers_24\[18\]
+ VGND VGND VPWR VPWR _12010_ sky130_fd_sc_hd__o22a_1
X_25229_ _08068_ net914 _08837_ VGND VGND VPWR VPWR _08844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_357_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_357_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_176_Right_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17982_ decode.regfile.registers_14\[30\] _10619_ _12589_ _10612_ VGND VGND VPWR
+ VPWR _03379_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19721_ _04992_ _04993_ _04994_ _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__a31o_1
X_28919_ clknet_leaf_117_clock _01932_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_16933_ decode.regfile.registers_9\[4\] _12607_ _12891_ _12893_ _12600_ VGND VGND
+ VPWR VPWR _12894_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_196_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29899_ clknet_leaf_340_clock _02912_ VGND VGND VPWR VPWR decode.regfile.registers_20\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19652_ _03918_ _04200_ _04204_ _04930_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__a31o_1
X_16864_ _12564_ VGND VGND VPWR VPWR _12826_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_221_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18603_ _03900_ _03700_ _03688_ decode.id_ex_rs1_data_reg\[19\] _03901_ VGND VGND
+ VPWR VPWR _03902_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_189_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15815_ decode.regfile.registers_14\[13\] _11207_ _11273_ decode.regfile.registers_15\[13\]
+ _11361_ VGND VGND VPWR VPWR _11799_ sky130_fd_sc_hd__a221o_1
XFILLER_0_205_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16795_ _12690_ VGND VGND VPWR VPWR _12759_ sky130_fd_sc_hd__clkbuf_4
X_19583_ _04209_ _03933_ _04197_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15746_ decode.regfile.registers_3\[11\] _11614_ _11367_ _11178_ VGND VGND VPWR VPWR
+ _11732_ sky130_fd_sc_hd__o2bb2a_1
X_18534_ memory.csr_read_data_out_reg\[25\] _09987_ _10110_ VGND VGND VPWR VPWR _03833_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_220_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15677_ _11198_ _11662_ _11663_ _11664_ VGND VGND VPWR VPWR _11665_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18465_ _03763_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14628_ _10670_ decode.id_ex_memread_reg VGND VGND VPWR VPWR _10671_ sky130_fd_sc_hd__and2b_1
XFILLER_0_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17416_ _13081_ _13168_ decode.regfile.registers_23\[15\] _13041_ VGND VGND VPWR
+ VPWR _13366_ sky130_fd_sc_hd__or4_1
XFILLER_0_157_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18396_ _03681_ _03676_ _03694_ _03677_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_157_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17347_ _13215_ decode.regfile.registers_28\[13\] _13093_ VGND VGND VPWR VPWR _13299_
+ sky130_fd_sc_hd__o21a_1
X_14559_ _10601_ VGND VGND VPWR VPWR _10602_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17278_ decode.regfile.registers_6\[12\] _12735_ _13226_ _13230_ VGND VGND VPWR VPWR
+ _13231_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19017_ _03972_ _03974_ _04007_ net243 VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16229_ _11942_ decode.regfile.registers_30\[24\] _12095_ _12096_ _12097_ VGND VGND
+ VPWR VPWR _12202_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_228_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_228_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_181_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19919_ _05184_ _05186_ _04526_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_177_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22930_ _07368_ _07379_ _05246_ _07380_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_78_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22861_ net2074 _10803_ _07324_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24600_ _08482_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21812_ csr._mcycle_T_2\[7\] _06476_ _06460_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25580_ net2254 _09052_ _09054_ _09046_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22792_ net1096 _10878_ _07286_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24531_ _08091_ net1129 _08439_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21743_ net1821 _10812_ _06428_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27250_ clknet_leaf_32_clock _00279_ VGND VGND VPWR VPWR decode.regfile.registers_30\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_24462_ _08410_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21674_ csr._mcycle_T_2\[21\] _06320_ _06381_ csr.minstret\[21\] VGND VGND VPWR VPWR
+ _06382_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_43_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26201_ _09420_ _09413_ VGND VGND VPWR VPWR _09421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23413_ fetch.bht.bhtTable_target_pc\[0\]\[31\] fetch.bht.bhtTable_target_pc\[1\]\[31\]
+ fetch.bht.bhtTable_target_pc\[2\]\[31\] fetch.bht.bhtTable_target_pc\[3\]\[31\]
+ _07066_ _07070_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27181_ clknet_leaf_355_clock _00210_ VGND VGND VPWR VPWR decode.regfile.registers_27\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20625_ _05759_ _05671_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__nor2_1
X_24393_ net883 execute.io_target_pc\[19\] _08367_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26132_ _09371_ VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__buf_4
X_23344_ net220 net221 _07728_ net85 VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__a31o_1
XFILLER_0_172_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20556_ csr.minstret\[16\] _05573_ _05585_ csr.mcycle\[16\] _05699_ VGND VGND VPWR
+ VPWR _05700_ sky130_fd_sc_hd__a221o_1
XFILLER_0_225_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26063_ net2562 _09329_ _09332_ _09333_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23275_ _06248_ VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__buf_2
X_20487_ csr._csr_read_data_T_8\[7\] _05591_ _05516_ _05528_ _05639_ VGND VGND VPWR
+ VPWR _05640_ sky130_fd_sc_hd__a41o_1
XFILLER_0_85_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25014_ csr._mcycle_T_2\[9\] _08712_ _08635_ csr.mcycle\[8\] csr.mcycle\[9\] VGND
+ VGND VPWR VPWR _08723_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_123_1308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22226_ _06718_ _06717_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_225_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29822_ clknet_leaf_315_clock _02835_ VGND VGND VPWR VPWR decode.regfile.registers_18\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_22157_ _06632_ _06747_ _06749_ _06751_ _06642_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_121_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21108_ _06045_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29753_ clknet_leaf_311_clock _02766_ VGND VGND VPWR VPWR decode.regfile.registers_15\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_22088_ fetch.bht.bhtTable_tag\[6\]\[7\] fetch.bht.bhtTable_tag\[7\]\[7\] _06644_
+ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__mux2_1
X_26965_ net898 _09853_ _09864_ _09865_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__o211a_1
X_28704_ clknet_leaf_171_clock _01717_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_13930_ net1791 _10213_ _10217_ _10206_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25916_ _08914_ _09243_ VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__nand2_1
X_21039_ execute.csr_read_data_out_reg\[9\] _06002_ _05998_ VGND VGND VPWR VPWR _06005_
+ sky130_fd_sc_hd__and3_1
X_29684_ clknet_leaf_282_clock _02697_ VGND VGND VPWR VPWR decode.regfile.registers_13\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_26896_ _09424_ _09819_ VGND VGND VPWR VPWR _09826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28635_ clknet_leaf_173_clock _01648_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_13861_ net1927 _10167_ _10176_ _10175_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__o211a_1
X_25847_ _08920_ _09200_ VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15600_ _11588_ _11315_ _11589_ VGND VGND VPWR VPWR _11590_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16580_ _12544_ VGND VGND VPWR VPWR _12545_ sky130_fd_sc_hd__clkbuf_4
X_28566_ clknet_leaf_207_clock _01579_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13792_ _10128_ _09937_ VGND VGND VPWR VPWR _10129_ sky130_fd_sc_hd__nand2_1
X_25778_ _09128_ VGND VGND VPWR VPWR _09169_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15531_ decode.regfile.registers_26\[5\] _11081_ _11522_ _11235_ _11350_ VGND VGND
+ VPWR VPWR _11523_ sky130_fd_sc_hd__a221o_1
X_24729_ _08091_ net1576 _08542_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27517_ clknet_leaf_29_clock _00546_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dfxtp_1
X_28497_ clknet_leaf_188_clock _01510_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18250_ _03581_ _03583_ decode.id_ex_funct3_reg\[0\] VGND VGND VPWR VPWR _03584_
+ sky130_fd_sc_hd__and3b_1
X_27448_ clknet_leaf_149_clock _00477_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_15462_ _11269_ VGND VGND VPWR VPWR _11455_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_210_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_281_clock clknet_5_21__leaf_clock VGND VGND VPWR VPWR clknet_leaf_281_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17201_ decode.regfile.registers_13\[10\] _12533_ _12582_ _12662_ VGND VGND VPWR
+ VPWR _13156_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14413_ _10112_ _10487_ VGND VGND VPWR VPWR _10497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18181_ _10944_ _10941_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__or2b_1
XFILLER_0_155_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15393_ _11358_ _11387_ _11268_ VGND VGND VPWR VPWR _11388_ sky130_fd_sc_hd__a21oi_1
X_27379_ clknet_leaf_15_clock _00408_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[20\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_182_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17132_ _13087_ decode.regfile.registers_26\[8\] _12814_ _13047_ _13088_ VGND VGND
+ VPWR VPWR _13089_ sky130_fd_sc_hd__o2111a_1
X_29118_ clknet_leaf_69_clock _02131_ VGND VGND VPWR VPWR csr.mcycle\[2\] sky130_fd_sc_hd__dfxtp_1
X_14344_ _10128_ _10418_ VGND VGND VPWR VPWR _10457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_1232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29049_ clknet_leaf_127_clock _02062_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17063_ decode.regfile.registers_7\[7\] _10616_ _13020_ VGND VGND VPWR VPWR _13021_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_80_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_296_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_296_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14275_ net608 _10377_ _10416_ _10411_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16014_ _11296_ _11990_ _11991_ _11992_ _11614_ VGND VGND VPWR VPWR _11993_ sky130_fd_sc_hd__a311o_1
XFILLER_0_208_1287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_223_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_223_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ decode.regfile.registers_21\[29\] _12716_ _03338_ _03362_ _12909_ VGND VGND
+ VPWR VPWR _03363_ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19704_ _04446_ _04976_ _04979_ _04980_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__o31a_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16916_ decode.regfile.registers_11\[4\] _12595_ _12876_ _12551_ VGND VGND VPWR VPWR
+ _12877_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17896_ _12968_ _03293_ _03294_ _03295_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19635_ _04911_ _04913_ _04401_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__a211oi_2
Xclkbuf_leaf_234_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_234_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16847_ _12769_ _12808_ _12809_ VGND VGND VPWR VPWR _12810_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_178_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_215_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19566_ _04332_ _04790_ _04848_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_69_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16778_ decode.regfile.registers_9\[1\] _12497_ _12503_ _12510_ _12652_ VGND VGND
+ VPWR VPWR _12742_ sky130_fd_sc_hd__o41a_1
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18517_ net202 VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__buf_4
XFILLER_0_186_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15729_ _11435_ _11089_ decode.regfile.registers_23\[10\] _11087_ VGND VGND VPWR
+ VPWR _11716_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19497_ _04107_ _04757_ _04781_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_201_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_249_clock clknet_5_19__leaf_clock VGND VGND VPWR VPWR clknet_leaf_249_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_174_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18448_ _03746_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18379_ decode.io_wb_rd\[0\] decode.id_ex_ex_rs1_reg\[0\] VGND VGND VPWR VPWR _03678_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20410_ _05439_ _05569_ _05425_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_212_Right_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21390_ _06138_ net2113 _06199_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20341_ _05398_ _05412_ _03517_ _03551_ _05507_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23060_ _06718_ _07472_ net68 VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__a21oi_1
X_20272_ _10706_ decode.id_ex_pc_reg\[10\] _10689_ _05440_ _10694_ VGND VGND VPWR
+ VPWR _05455_ sky130_fd_sc_hd__a41o_1
XFILLER_0_4_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22011_ net1957 _06600_ _06610_ _06605_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2501 decode.regfile.registers_0\[8\] VGND VGND VPWR VPWR net2728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2512 execute.csr_read_data_out_reg\[1\] VGND VGND VPWR VPWR net2739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2523 fetch.btb.btbTable\[15\]\[1\] VGND VGND VPWR VPWR net2750 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2534 decode.regfile.registers_11\[9\] VGND VGND VPWR VPWR net2761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2545 decode.io_id_pc\[31\] VGND VGND VPWR VPWR net2772 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1800 decode.regfile.registers_21\[22\] VGND VGND VPWR VPWR net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1811 fetch.bht.bhtTable_tag\[14\]\[18\] VGND VGND VPWR VPWR net2038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2556 decode.control.io_funct7\[4\] VGND VGND VPWR VPWR net2783 sky130_fd_sc_hd__dlygate4sd3_1
X_26750_ net2410 _09736_ _09741_ _09730_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__o211a_1
X_23962_ _08151_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__clkbuf_1
Xhold1822 fetch.bht.bhtTable_tag\[14\]\[11\] VGND VGND VPWR VPWR net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2567 decode.regfile.registers_30\[19\] VGND VGND VPWR VPWR net2794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1833 fetch.bht.bhtTable_tag\[5\]\[21\] VGND VGND VPWR VPWR net2060 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1844 decode.regfile.registers_14\[13\] VGND VGND VPWR VPWR net2071 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25701_ _08925_ _09122_ VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__nand2_1
Xhold1855 fetch.bht.bhtTable_target_pc\[10\]\[21\] VGND VGND VPWR VPWR net2082 sky130_fd_sc_hd__dlygate4sd3_1
X_22913_ net69 _06794_ _06862_ net222 VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__o22a_1
Xhold1866 fetch.bht.bhtTable_tag\[4\]\[23\] VGND VGND VPWR VPWR net2093 sky130_fd_sc_hd__dlygate4sd3_1
X_26681_ _09701_ VGND VGND VPWR VPWR _09702_ sky130_fd_sc_hd__clkbuf_4
X_23893_ net1769 _08051_ _06179_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__mux2_1
Xhold1877 decode.regfile.registers_24\[17\] VGND VGND VPWR VPWR net2104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1888 fetch.bht.bhtTable_tag\[0\]\[13\] VGND VGND VPWR VPWR net2115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28420_ clknet_leaf_39_clock _01433_ VGND VGND VPWR VPWR decode.immGen._imm_T_10\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25632_ net1513 _09082_ _09084_ _09074_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__o211a_1
Xhold1899 decode.regfile.registers_30\[3\] VGND VGND VPWR VPWR net2126 sky130_fd_sc_hd__dlygate4sd3_1
X_22844_ net760 _10817_ _09898_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28351_ clknet_leaf_167_clock _01364_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25563_ net1981 _09039_ _09044_ _09033_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22775_ _06149_ net970 _07276_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27302_ clknet_leaf_14_clock _00331_ VGND VGND VPWR VPWR decode.regfile.registers_31\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_24514_ _08074_ net2139 _08428_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__mux2_1
X_28282_ clknet_leaf_85_clock _01304_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_21726_ csr.msie csr.msip csr.ie execute.exception_out_reg _06031_ VGND VGND VPWR
+ VPWR _06423_ sky130_fd_sc_hd__a311oi_1
X_25494_ net2545 _08995_ _09003_ _09004_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27233_ clknet_leaf_364_clock _00262_ VGND VGND VPWR VPWR decode.regfile.registers_29\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_24445_ _08072_ net1897 _08400_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21657_ _03580_ _06368_ _06369_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__nor3_1
XFILLER_0_19_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20608_ _05516_ _03755_ _05527_ _05744_ _05555_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__a41o_1
X_27164_ clknet_leaf_360_clock _00193_ VGND VGND VPWR VPWR decode.regfile.registers_27\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24376_ net955 execute.io_target_pc\[11\] _08356_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21588_ csr.io_csr_write_address\[11\] net352 _06314_ _06316_ VGND VGND VPWR VPWR
+ _06317_ sky130_fd_sc_hd__nand4_4
X_26115_ decode.regfile.registers_10\[24\] _09356_ _09362_ _09359_ VGND VGND VPWR
+ VPWR _02599_ sky130_fd_sc_hd__o211a_1
X_23327_ fetch.bht.bhtTable_target_pc\[6\]\[25\] fetch.bht.bhtTable_target_pc\[7\]\[25\]
+ _07106_ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20539_ csr.mcycle\[14\] _05588_ _05575_ csr.minstret\[14\] VGND VGND VPWR VPWR _05685_
+ sky130_fd_sc_hd__a22o_1
X_27095_ clknet_leaf_350_clock _00124_ VGND VGND VPWR VPWR decode.regfile.registers_25\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14060_ _09975_ _10288_ VGND VGND VPWR VPWR _10294_ sky130_fd_sc_hd__nand2_1
X_26046_ net2544 _09313_ _09322_ _09318_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__o211a_1
X_23258_ net80 net79 net224 _07636_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__nand4_1
XFILLER_0_132_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22209_ _06802_ _06803_ _06628_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__mux2_1
X_23189_ fetch.bht.bhtTable_target_pc\[0\]\[17\] fetch.bht.bhtTable_target_pc\[1\]\[17\]
+ fetch.bht.bhtTable_target_pc\[2\]\[17\] fetch.bht.bhtTable_target_pc\[3\]\[17\]
+ _07384_ _07113_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29805_ clknet_leaf_296_clock _02818_ VGND VGND VPWR VPWR decode.regfile.registers_17\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27997_ clknet_leaf_213_clock _01019_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17750_ decode.regfile.registers_3\[24\] _10616_ _12729_ _12838_ VGND VGND VPWR VPWR
+ _03153_ sky130_fd_sc_hd__a31o_1
X_14962_ _10987_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__clkbuf_1
X_29736_ clknet_leaf_285_clock _02749_ VGND VGND VPWR VPWR decode.regfile.registers_15\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_26948_ _10041_ _09849_ VGND VGND VPWR VPWR _09856_ sky130_fd_sc_hd__nand2_1
X_16701_ _12650_ VGND VGND VPWR VPWR _12666_ sky130_fd_sc_hd__clkbuf_4
X_13913_ _09999_ _10200_ VGND VGND VPWR VPWR _10208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29667_ clknet_leaf_287_clock _02680_ VGND VGND VPWR VPWR decode.regfile.registers_13\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_14893_ _10929_ VGND VGND VPWR VPWR _10930_ sky130_fd_sc_hd__clkbuf_4
X_17681_ _12888_ _03084_ _03085_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_528 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26879_ _09406_ _09806_ VGND VGND VPWR VPWR _09816_ sky130_fd_sc_hd__nand2_1
X_19420_ _04646_ _04463_ _04289_ _04707_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__a2bb2o_1
X_28618_ clknet_leaf_100_clock _01631_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_16632_ decode.immGen._imm_T_24\[19\] decode.immGen._imm_T_24\[15\] VGND VGND VPWR
+ VPWR _12597_ sky130_fd_sc_hd__nor2_4
X_13844_ _10152_ VGND VGND VPWR VPWR _10167_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29598_ clknet_leaf_270_clock _02611_ VGND VGND VPWR VPWR decode.regfile.registers_11\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19351_ _04130_ _04131_ _04612_ _04621_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__a2bb2o_1
X_28549_ clknet_leaf_174_clock _01562_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_16563_ _12527_ VGND VGND VPWR VPWR _12528_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13775_ _10060_ memory.io_wb_aluresult\[26\] _10004_ memory.io_wb_readdata\[26\]
+ _10005_ VGND VGND VPWR VPWR _10114_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18302_ _03595_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__buf_2
XFILLER_0_167_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15514_ _10648_ _10624_ _11084_ _11505_ VGND VGND VPWR VPWR _11506_ sky130_fd_sc_hd__o31a_1
XFILLER_0_169_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19282_ _04244_ _04510_ _04573_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__nand3_1
X_16494_ decode.regfile.registers_3\[31\] _11292_ _11293_ _10635_ VGND VGND VPWR VPWR
+ _12460_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_31_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18233_ csr._mcycle_T_3\[63\] csr._mcycle_T_3\[62\] csr._mcycle_T_3\[61\] csr._mcycle_T_3\[58\]
+ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__or4_1
X_15445_ _11250_ decode.regfile.registers_27\[3\] _11258_ VGND VGND VPWR VPWR _11439_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_154_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18164_ _03463_ _03464_ _10921_ decode.control.io_funct7\[1\] VGND VGND VPWR VPWR
+ _03510_ sky130_fd_sc_hd__and4bb_1
X_15376_ _11153_ VGND VGND VPWR VPWR _11371_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17115_ decode.regfile.registers_15\[8\] _12667_ _12773_ _13011_ VGND VGND VPWR VPWR
+ _13072_ sky130_fd_sc_hd__o31a_1
X_14327_ _10087_ _10444_ VGND VGND VPWR VPWR _10448_ sky130_fd_sc_hd__nand2_1
X_18095_ _03473_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold407 decode.regfile.registers_31\[30\] VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 csr._mcycle_T_3\[36\] VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17046_ decode.regfile.registers_27\[6\] _12507_ _12520_ _12967_ _13004_ VGND VGND
+ VPWR VPWR _13005_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_225_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold429 decode.regfile.registers_3\[5\] VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14258_ net1508 _10403_ _10407_ _10398_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14189_ _10122_ _10355_ VGND VGND VPWR VPWR _10367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_209_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18997_ _04255_ _03983_ _04248_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__or3_1
XFILLER_0_225_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1107 fetch.bht.bhtTable_tag\[0\]\[16\] VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_163_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 fetch.bht.bhtTable_target_pc\[3\]\[20\] VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ _12732_ _03341_ _03344_ _03345_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_173_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_173_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1129 fetch.bht.bhtTable_target_pc\[11\]\[19\] VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17879_ decode.regfile.registers_11\[27\] _12792_ _03267_ _03278_ VGND VGND VPWR
+ VPWR _03279_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_75_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19618_ _04199_ _03923_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_176_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20890_ _05858_ _05921_ net62 VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_188_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_188_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_177_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19549_ _04829_ _04831_ _04211_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_193_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22560_ csr._minstret_T_3\[37\] csr._minstret_T_3\[36\] _07144_ VGND VGND VPWR VPWR
+ _07147_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_360 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21511_ _06140_ net2086 _06263_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_371 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_382 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22491_ _07077_ _07083_ _07085_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_111_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_111_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_185_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24230_ _08057_ net2189 _08289_ VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__mux2_1
X_21442_ _06236_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24161_ _08055_ net1973 _06274_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21373_ _06187_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_20_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23112_ execute.io_target_pc\[12\] _07345_ _05864_ _07552_ VGND VGND VPWR VPWR _07553_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20324_ _05493_ _05494_ _05416_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_9_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_126_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_126_clock
+ sky130_fd_sc_hd__clkbuf_8
X_24092_ _08218_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold930 decode.regfile.registers_22\[6\] VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_222_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold941 fetch.bht.bhtTable_tag\[4\]\[4\] VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold952 fetch.bht.bhtTable_target_pc\[8\]\[2\] VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold963 fetch.bht.bhtTable_target_pc\[3\]\[23\] VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__dlygate4sd3_1
X_23043_ net97 _07343_ _07344_ _07487_ _06566_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__o311a_1
X_27920_ clknet_leaf_69_clock _00949_ VGND VGND VPWR VPWR csr.io_csr_write_address\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_20255_ _10678_ _10730_ _05430_ decode.id_ex_pc_reg\[8\] VGND VGND VPWR VPWR _05442_
+ sky130_fd_sc_hd__a31o_1
Xhold974 fetch.bht.bhtTable_target_pc\[1\]\[30\] VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 decode.regfile.registers_13\[28\] VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 fetch.bht.bhtTable_tag\[11\]\[22\] VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20186_ decode.id_ex_imm_reg\[27\] _10854_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__nand2_1
X_27851_ clknet_leaf_323_clock _00880_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2320 decode.regfile.registers_22\[21\] VGND VGND VPWR VPWR net2547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2331 decode.regfile.registers_0\[3\] VGND VGND VPWR VPWR net2558 sky130_fd_sc_hd__dlygate4sd3_1
X_26802_ _09404_ _09763_ VGND VGND VPWR VPWR _09772_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_95_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2342 csr._csr_read_data_T_8\[21\] VGND VGND VPWR VPWR net2569 sky130_fd_sc_hd__dlygate4sd3_1
X_24994_ _08633_ csr.mcycle\[1\] csr.mcycle\[2\] csr.mcycle\[0\] VGND VGND VPWR VPWR
+ _08709_ sky130_fd_sc_hd__and4_1
X_27782_ clknet_leaf_333_clock _00811_ VGND VGND VPWR VPWR memory.io_wb_readdata\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2353 decode.regfile.registers_5\[29\] VGND VGND VPWR VPWR net2580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2364 decode.regfile.registers_11\[16\] VGND VGND VPWR VPWR net2591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1630 fetch.bht.bhtTable_target_pc\[15\]\[5\] VGND VGND VPWR VPWR net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2375 decode.regfile.registers_7\[21\] VGND VGND VPWR VPWR net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1641 fetch.bht.bhtTable_target_pc\[12\]\[30\] VGND VGND VPWR VPWR net1868 sky130_fd_sc_hd__dlygate4sd3_1
X_29521_ clknet_leaf_266_clock _02534_ VGND VGND VPWR VPWR decode.regfile.registers_8\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_23945_ net1119 _08103_ _06156_ VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__mux2_1
Xhold2386 csr.msip VGND VGND VPWR VPWR net2613 sky130_fd_sc_hd__dlygate4sd3_1
X_26733_ _09410_ _09720_ VGND VGND VPWR VPWR _09732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2397 csr.mscratch\[29\] VGND VGND VPWR VPWR net2624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1652 fetch.bht.bhtTable_tag\[8\]\[6\] VGND VGND VPWR VPWR net1879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1663 decode.regfile.registers_6\[6\] VGND VGND VPWR VPWR net1890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1674 fetch.bht.bhtTable_target_pc\[6\]\[10\] VGND VGND VPWR VPWR net1901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1685 _02154_ VGND VGND VPWR VPWR net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1696 fetch.bht.bhtTable_target_pc\[2\]\[9\] VGND VGND VPWR VPWR net1923 sky130_fd_sc_hd__dlygate4sd3_1
X_26664_ _09664_ VGND VGND VPWR VPWR _09692_ sky130_fd_sc_hd__buf_2
X_29452_ clknet_leaf_261_clock _02465_ VGND VGND VPWR VPWR decode.regfile.registers_6\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_23876_ execute.io_target_pc\[27\] VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28403_ clknet_leaf_142_clock _01416_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_2
X_25615_ _08914_ _09069_ VGND VGND VPWR VPWR _09075_ sky130_fd_sc_hd__nand2_1
X_22827_ _07309_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__clkbuf_1
X_29383_ clknet_leaf_258_clock _02396_ VGND VGND VPWR VPWR decode.regfile.registers_4\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_26595_ decode.regfile.registers_16\[22\] _09649_ _09652_ _09648_ VGND VGND VPWR
+ VPWR _02789_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28334_ clknet_leaf_235_clock _01347_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13560_ _09926_ execute.io_mem_memwrite VGND VGND VPWR VPWR _09927_ sky130_fd_sc_hd__and2b_1
X_25546_ _08920_ _09026_ VGND VGND VPWR VPWR _09035_ sky130_fd_sc_hd__nand2_1
X_22758_ _06132_ net1362 _07265_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21709_ csr.minstret\[25\] _06407_ _06409_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28265_ clknet_leaf_64_clock net2646 VGND VGND VPWR VPWR csr._csr_read_data_T_8\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_192_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25477_ _08978_ VGND VGND VPWR VPWR _08995_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22689_ csr._mcycle_T_2\[20\] _07223_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_229_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15230_ _11226_ VGND VGND VPWR VPWR _11227_ sky130_fd_sc_hd__clkbuf_4
X_24428_ _08055_ net1777 _08389_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27216_ clknet_leaf_6_clock _00245_ VGND VGND VPWR VPWR decode.regfile.registers_29\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28196_ clknet_leaf_59_clock _01218_ VGND VGND VPWR VPWR csr.io_mret_vector\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15161_ decode.regfile.registers_1\[0\] _11116_ _11137_ _11157_ VGND VGND VPWR VPWR
+ _11158_ sky130_fd_sc_hd__and4_1
X_27147_ clknet_leaf_357_clock _00176_ VGND VGND VPWR VPWR decode.regfile.registers_26\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_24359_ _09910_ VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14112_ _10117_ _10312_ VGND VGND VPWR VPWR _10323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27078_ clknet_leaf_346_clock _00107_ VGND VGND VPWR VPWR decode.regfile.registers_24\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_15092_ _10657_ _10977_ _11060_ _10662_ VGND VGND VPWR VPWR _11089_ sky130_fd_sc_hd__or4b_4
XFILLER_0_120_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14043_ net2464 _10271_ _10282_ _10275_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__o211a_1
X_26029_ _09285_ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__clkbuf_4
X_18920_ _03811_ _03827_ _03826_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_90_clock clknet_5_8__leaf_clock VGND VGND VPWR VPWR clknet_leaf_90_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18851_ net308 _04147_ _03706_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17802_ _11020_ _12490_ _12512_ decode.regfile.registers_12\[25\] _12591_ VGND VGND
+ VPWR VPWR _03204_ sky130_fd_sc_hd__o32a_1
XFILLER_0_175_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18782_ decode.id_ex_rs1_data_reg\[14\] _03908_ net334 _03700_ _04080_ VGND VGND
+ VPWR VPWR _04081_ sky130_fd_sc_hd__o221ai_4
X_15994_ _11947_ _11973_ _11096_ VGND VGND VPWR VPWR _11974_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17733_ _11014_ _10936_ decode.regfile.registers_23\[23\] _12995_ VGND VGND VPWR
+ VPWR _03137_ sky130_fd_sc_hd__or4_1
X_29719_ clknet_leaf_284_clock _02732_ VGND VGND VPWR VPWR decode.regfile.registers_14\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14945_ _10667_ _10967_ _10952_ _10969_ _10973_ VGND VGND VPWR VPWR _10974_ sky130_fd_sc_hd__o41a_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17664_ _13215_ decode.regfile.registers_28\[21\] _02992_ VGND VGND VPWR VPWR _03070_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_218_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14876_ _10917_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_218_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19403_ _04691_ _04592_ _04269_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16615_ _12579_ VGND VGND VPWR VPWR _12580_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13827_ net2474 _10153_ _10157_ _10132_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__o211a_1
X_17595_ decode.regfile.registers_2\[20\] _12834_ _12639_ decode.regfile.registers_3\[20\]
+ _12838_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_106_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_214_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19334_ _04270_ _04463_ _04625_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_214_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16546_ _12510_ VGND VGND VPWR VPWR _12511_ sky130_fd_sc_hd__buf_4
X_13758_ _10003_ memory.io_wb_aluresult\[23\] _10001_ memory.io_wb_reg_pc\[23\] _09995_
+ VGND VGND VPWR VPWR _10100_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19265_ _04518_ _04039_ _04519_ _04558_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a31oi_4
X_16477_ decode.regfile.registers_25\[30\] _11333_ _11336_ decode.regfile.registers_24\[30\]
+ VGND VGND VPWR VPWR _12444_ sky130_fd_sc_hd__o22a_1
X_13689_ _10041_ VGND VGND VPWR VPWR _10042_ sky130_fd_sc_hd__buf_4
XFILLER_0_215_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18216_ _11149_ _03548_ _03549_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__nor3_1
XFILLER_0_155_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15428_ decode.regfile.registers_13\[3\] _11276_ _11407_ decode.regfile.registers_12\[3\]
+ _11421_ VGND VGND VPWR VPWR _11422_ sky130_fd_sc_hd__a221o_1
X_19196_ _03637_ _04306_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_clock clknet_5_7__leaf_clock VGND VGND VPWR VPWR clknet_leaf_43_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18147_ _03495_ _03493_ _03500_ net1984 VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__and4bb_1
X_15359_ _10662_ _10657_ _11048_ _11104_ VGND VGND VPWR VPWR _11354_ sky130_fd_sc_hd__or4_4
XFILLER_0_223_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold204 decode.regfile.registers_31\[14\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_TAPCELL_ROW_169_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold215 _11842_ VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18078_ _10997_ _10969_ _11034_ _03462_ _10999_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__o41a_1
Xhold226 decode.regfile.registers_27\[7\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 decode.regfile.registers_30\[11\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold248 csr._mcycle_T_3\[42\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 decode.regfile.registers_1\[22\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ _12674_ _12986_ _12987_ VGND VGND VPWR VPWR _12988_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_165_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_58_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20040_ decode.id_ex_imm_reg\[6\] decode.id_ex_pc_reg\[6\] VGND VGND VPWR VPWR _05261_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21991_ net1206 _06588_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23730_ _08016_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_124_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _05952_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23661_ net1264 _10787_ _07972_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20873_ _05914_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25400_ _10068_ VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22612_ _06377_ _07183_ _07185_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__nor3_1
XFILLER_0_7_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26380_ _09436_ _09490_ VGND VGND VPWR VPWR _09528_ sky130_fd_sc_hd__nand2_1
X_23592_ _06122_ net2058 _07941_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25331_ _08896_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22543_ csr.minstret\[30\] csr.minstret\[31\] _06417_ VGND VGND VPWR VPWR _07136_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_174_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_190 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28050_ clknet_leaf_221_clock _01072_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25262_ _08101_ net1447 _09906_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22474_ _07068_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27001_ clknet_leaf_338_clock _00030_ VGND VGND VPWR VPWR decode.regfile.registers_22\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_24213_ _08107_ net1507 _06251_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__mux2_1
X_21425_ _06227_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__clkbuf_1
X_25193_ _08825_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24144_ _08245_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21356_ _06190_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20307_ _05481_ _05219_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__nor2_1
X_28952_ clknet_leaf_120_clock _01965_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_24075_ net1749 execute.io_target_pc\[25\] _07991_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold760 fetch.bht.bhtTable_target_pc\[1\]\[27\] VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__dlygate4sd3_1
X_21287_ _10777_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold771 fetch.bht.bhtTable_tag\[2\]\[0\] VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold782 csr.minstret\[30\] VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27903_ clknet_leaf_89_clock _00932_ VGND VGND VPWR VPWR csr._mcycle_T_2\[24\] sky130_fd_sc_hd__dfxtp_2
X_23026_ net97 _07464_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20238_ _05427_ _05428_ _05415_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__o21a_1
Xhold793 decode.id_ex_isbranch_reg VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__dlygate4sd3_1
X_28883_ clknet_leaf_140_clock _01896_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27834_ clknet_leaf_324_clock _00863_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_20169_ decode.id_ex_imm_reg\[23\] _10786_ _05371_ _05365_ VGND VGND VPWR VPWR _05372_
+ sky130_fd_sc_hd__o22ai_2
Xhold2150 decode.regfile.registers_13\[21\] VGND VGND VPWR VPWR net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2161 decode.regfile.registers_14\[1\] VGND VGND VPWR VPWR net2388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2172 decode.regfile.registers_9\[0\] VGND VGND VPWR VPWR net2399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2183 decode.regfile.registers_18\[24\] VGND VGND VPWR VPWR net2410 sky130_fd_sc_hd__dlygate4sd3_1
X_27765_ clknet_leaf_323_clock _00794_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_24977_ net2548 _08696_ _08697_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__o21ba_1
Xhold2194 decode.regfile.registers_12\[11\] VGND VGND VPWR VPWR net2421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1460 fetch.bht.bhtTable_target_pc\[9\]\[20\] VGND VGND VPWR VPWR net1687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29504_ clknet_leaf_250_clock _02517_ VGND VGND VPWR VPWR decode.regfile.registers_8\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1471 fetch.bht.bhtTable_tag\[15\]\[20\] VGND VGND VPWR VPWR net1698 sky130_fd_sc_hd__dlygate4sd3_1
X_14730_ csr.io_mem_pc\[25\] VGND VGND VPWR VPWR _10773_ sky130_fd_sc_hd__buf_4
X_26716_ net1449 _09709_ _09722_ _09717_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__o211a_1
X_23928_ _08134_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__clkbuf_1
Xhold1482 decode.regfile.registers_26\[31\] VGND VGND VPWR VPWR net1709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1493 fetch.bht.bhtTable_target_pc\[13\]\[18\] VGND VGND VPWR VPWR net1720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27696_ clknet_leaf_21_clock _00725_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14661_ decode.id_ex_pc_reg\[5\] VGND VGND VPWR VPWR _10704_ sky130_fd_sc_hd__clkbuf_4
X_29435_ clknet_leaf_250_clock _02448_ VGND VGND VPWR VPWR decode.regfile.registers_6\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23859_ _08093_ net1855 _08079_ VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26647_ net711 _09679_ _09682_ _09675_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16400_ decode.regfile.registers_19\[28\] _11453_ _11219_ _12368_ VGND VGND VPWR
+ VPWR _12369_ sky130_fd_sc_hd__o211a_1
X_13612_ memory.csr_read_data_out_reg\[3\] _09941_ _09972_ _09973_ VGND VGND VPWR
+ VPWR _09974_ sky130_fd_sc_hd__o22ai_4
X_29366_ clknet_leaf_227_clock _02379_ VGND VGND VPWR VPWR decode.regfile.registers_3\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14592_ decode.immGen._imm_T_24\[11\] VGND VGND VPWR VPWR _10635_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ decode.regfile.registers_23\[14\] _12714_ _13305_ _13330_ _12515_ VGND VGND
+ VPWR VPWR _13331_ sky130_fd_sc_hd__o221a_1
X_26578_ net611 _09636_ _09642_ _09635_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28317_ clknet_leaf_211_clock _01330_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13543_ _09914_ _09887_ _09916_ net388 VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__a31o_1
X_16331_ _11232_ _12300_ _12301_ VGND VGND VPWR VPWR _12302_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25529_ _09949_ VGND VGND VPWR VPWR _09025_ sky130_fd_sc_hd__buf_4
X_29297_ clknet_leaf_224_clock _02310_ VGND VGND VPWR VPWR decode.regfile.registers_1\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19050_ _04240_ _04348_ _03588_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__a21oi_4
X_16262_ _11396_ _12232_ _12233_ _12234_ VGND VGND VPWR VPWR _12235_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28248_ clknet_leaf_78_clock _01270_ VGND VGND VPWR VPWR csr._minstret_T_3\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15213_ _11189_ _11200_ _11203_ _11209_ VGND VGND VPWR VPWR _11210_ sky130_fd_sc_hd__a211o_1
X_18001_ decode.regfile.registers_21\[30\] _12716_ _03376_ _03397_ _13164_ VGND VGND
+ VPWR VPWR _03398_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_11_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16193_ _11445_ _12166_ _12167_ _11246_ VGND VGND VPWR VPWR _12168_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28179_ clknet_leaf_57_clock _01201_ VGND VGND VPWR VPWR csr.io_mret_vector\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15144_ _11140_ VGND VGND VPWR VPWR _11141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19952_ _05210_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__clkbuf_1
X_15075_ _11071_ VGND VGND VPWR VPWR _11072_ sky130_fd_sc_hd__buf_4
XFILLER_0_205_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14026_ net2416 _10271_ _10273_ _10262_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__o211a_1
X_18903_ _04201_ _03938_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__nor2_1
XFILLER_0_226_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19883_ _04359_ _03788_ _04444_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__o21ai_1
X_18834_ memory.csr_read_data_out_reg\[9\] _10010_ _10022_ _10023_ VGND VGND VPWR
+ VPWR _04133_ sky130_fd_sc_hd__o22a_4
XFILLER_0_207_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18765_ decode.id_ex_rs2_data_reg\[7\] _03746_ _03764_ _04060_ _04063_ VGND VGND
+ VPWR VPWR _04064_ sky130_fd_sc_hd__o221a_1
XFILLER_0_222_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15977_ decode.regfile.registers_2\[17\] _11295_ net347 _11121_ _11956_ VGND VGND
+ VPWR VPWR _11957_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17716_ decode.regfile.registers_0\[23\] _12932_ _12834_ _03119_ VGND VGND VPWR VPWR
+ _03120_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14928_ _10956_ VGND VGND VPWR VPWR _10957_ sky130_fd_sc_hd__clkbuf_4
X_18696_ _03662_ execute.io_reg_pc\[1\] _03992_ _03994_ VGND VGND VPWR VPWR _03995_
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17647_ _12666_ _12773_ _12984_ decode.regfile.registers_14\[21\] _03052_ VGND VGND
+ VPWR VPWR _03053_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_63_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14859_ decode.id_ex_pc_reg\[20\] _10866_ _10870_ decode.id_ex_pc_reg\[18\] _10901_
+ VGND VGND VPWR VPWR _10902_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17578_ _12494_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__buf_2
XFILLER_0_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19317_ _04290_ _04273_ _04480_ _04608_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16529_ _10926_ VGND VGND VPWR VPWR _12494_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19248_ _04542_ _04409_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19179_ _04244_ _04474_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21210_ _10596_ _05671_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_93_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22190_ net91 _06784_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21141_ _06062_ _06058_ net2395 VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21072_ _06022_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20023_ _10758_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__clkbuf_4
X_24900_ net581 _08647_ _07179_ VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_126_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25880_ net2570 _09226_ _09227_ _09222_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24831_ _06109_ net1602 _08422_ VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24762_ _08055_ net1930 _08563_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27550_ clknet_leaf_42_clock _00579_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_2
X_21974_ net1936 _06588_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer30 _04310_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_1
Xrebuffer41 _10762_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23713_ _08007_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26501_ net2472 _09592_ _09598_ _09595_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27481_ clknet_leaf_52_clock _00510_ VGND VGND VPWR VPWR decode.io_wfi_out sky130_fd_sc_hd__dfxtp_1
X_20925_ _05937_ _05933_ net48 VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__and3_1
Xrebuffer52 _04152_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_1
X_24693_ _08055_ net1494 _06306_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer63 _03759_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__buf_1
Xrebuffer74 _06615_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer85 net309 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29220_ clknet_leaf_109_clock _02233_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_23644_ net1012 _10872_ _07961_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__mux2_1
X_26432_ _09533_ VGND VGND VPWR VPWR _09558_ sky130_fd_sc_hd__buf_2
Xrebuffer96 net321 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20856_ _05905_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29151_ clknet_leaf_235_clock _02164_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_26363_ _09420_ _09515_ VGND VGND VPWR VPWR _09519_ sky130_fd_sc_hd__nand2_1
X_23575_ _07932_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20787_ _05866_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25314_ _08887_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__clkbuf_1
X_28102_ clknet_leaf_68_clock _01124_ VGND VGND VPWR VPWR csr.minstret\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22526_ fetch.bht.bhtTable_target_pc\[4\]\[1\] fetch.bht.bhtTable_target_pc\[5\]\[1\]
+ _07119_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29082_ clknet_leaf_190_clock _02095_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26294_ _09426_ _09472_ VGND VGND VPWR VPWR _09479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25245_ _08852_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__clkbuf_1
X_28033_ clknet_leaf_195_clock _01055_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer120 net346 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22457_ _06645_ fetch.btb.btbTable\[9\]\[1\] fetch.bht.bhtTable_valid\[9\] _07051_
+ _06631_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__a311o_1
XFILLER_0_122_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_6__f_clock clknet_2_0_0_clock VGND VGND VPWR VPWR clknet_5_6__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21408_ _06217_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__clkbuf_8
X_25176_ _10573_ net2612 _08816_ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__mux2_1
X_22388_ _06673_ _06982_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24127_ net967 execute.io_target_pc\[18\] _08232_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21339_ _06180_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24058_ _08201_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__clkbuf_1
X_28935_ clknet_leaf_113_clock _01948_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold590 decode.regfile.registers_20\[12\] VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23009_ fetch.bht.bhtTable_target_pc\[4\]\[7\] fetch.bht.bhtTable_target_pc\[5\]\[7\]
+ fetch.bht.bhtTable_target_pc\[6\]\[7\] fetch.bht.bhtTable_target_pc\[7\]\[7\] _07407_
+ _07072_ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__mux4_1
X_15900_ decode.regfile.registers_0\[15\] _11300_ _11129_ _11298_ VGND VGND VPWR VPWR
+ _11882_ sky130_fd_sc_hd__o2bb2ai_1
X_28866_ clknet_leaf_134_clock _01879_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16880_ _12592_ _12616_ _12547_ VGND VGND VPWR VPWR _12842_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_202_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15831_ decode.regfile.registers_12\[13\] _11689_ _11278_ _11814_ VGND VGND VPWR
+ VPWR _11815_ sky130_fd_sc_hd__o22a_1
X_27817_ clknet_leaf_323_clock _00846_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_28797_ clknet_leaf_179_clock _01810_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18550_ _03844_ _03847_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__nand2_1
X_15762_ decode.regfile.registers_20\[11\] _11219_ _11726_ _11747_ _11648_ VGND VGND
+ VPWR VPWR _11748_ sky130_fd_sc_hd__o221a_1
X_27748_ clknet_leaf_35_clock _00777_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_194_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1290 fetch.bht.bhtTable_tag\[8\]\[17\] VGND VGND VPWR VPWR net1517 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _13221_ _13446_ _13447_ _13448_ VGND VGND VPWR VPWR _13449_ sky130_fd_sc_hd__a31o_1
X_14713_ _10676_ _10686_ _10701_ _10755_ _09900_ VGND VGND VPWR VPWR _10756_ sky130_fd_sc_hd__a41oi_4
X_18481_ _03656_ _03779_ decode.id_ex_rs1_data_reg\[29\] _03689_ VGND VGND VPWR VPWR
+ _03780_ sky130_fd_sc_hd__o22ai_4
X_15693_ _11037_ VGND VGND VPWR VPWR _11681_ sky130_fd_sc_hd__clkbuf_4
X_27679_ clknet_leaf_28_clock _00708_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[21\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_213_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17432_ decode.regfile.registers_3\[16\] _12639_ _10609_ _12625_ VGND VGND VPWR VPWR
+ _13381_ sky130_fd_sc_hd__o2bb2a_1
X_29418_ clknet_leaf_257_clock _02431_ VGND VGND VPWR VPWR decode.regfile.registers_5\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14644_ execute.io_target_pc\[27\] VGND VGND VPWR VPWR _10687_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17363_ decode.regfile.registers_1\[14\] _12630_ _12829_ _10614_ _13313_ VGND VGND
+ VPWR VPWR _13314_ sky130_fd_sc_hd__o221a_1
X_29349_ clknet_leaf_228_clock _02362_ VGND VGND VPWR VPWR decode.regfile.registers_3\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14575_ _10617_ VGND VGND VPWR VPWR _10618_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_200_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19102_ _03637_ decode.id_ex_aluop_reg\[1\] decode.id_ex_aluop_reg\[3\] decode.id_ex_aluop_reg\[2\]
+ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__nor4_2
XFILLER_0_184_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16314_ decode.regfile.registers_5\[26\] _11192_ _11139_ _12283_ _12284_ VGND VGND
+ VPWR VPWR _12285_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13526_ net495 _09903_ VGND VGND VPWR VPWR _09904_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_153_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17294_ decode.regfile.registers_21\[12\] _12716_ _13222_ _13246_ _12806_ VGND VGND
+ VPWR VPWR _13247_ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19033_ _04248_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__buf_4
XFILLER_0_180_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16245_ decode.regfile.registers_11\[24\] _11180_ _11689_ _11280_ VGND VGND VPWR
+ VPWR _12218_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_70_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16176_ decode.regfile.registers_11\[22\] _11072_ _11204_ _11407_ _12150_ VGND VGND
+ VPWR VPWR _12151_ sky130_fd_sc_hd__a311o_1
XFILLER_0_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput106 net106 VGND VGND VPWR VPWR io_memory_address[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput117 net117 VGND VGND VPWR VPWR io_memory_address[25] sky130_fd_sc_hd__clkbuf_4
Xoutput128 net128 VGND VGND VPWR VPWR io_memory_address[6] sky130_fd_sc_hd__clkbuf_4
X_15127_ _11123_ VGND VGND VPWR VPWR _11124_ sky130_fd_sc_hd__clkbuf_4
Xoutput139 net139 VGND VGND VPWR VPWR io_memory_write_data[12] sky130_fd_sc_hd__clkbuf_4
X_15058_ decode.immGen._imm_T_24\[4\] VGND VGND VPWR VPWR _11055_ sky130_fd_sc_hd__inv_2
X_19935_ _09955_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14009_ _10053_ _10255_ VGND VGND VPWR VPWR _10264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19866_ _04243_ _04966_ _05135_ _04436_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_208_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18817_ _04115_ _04112_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__nor2_1
X_19797_ _03835_ _03812_ _04274_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18748_ _03715_ _03725_ _04041_ _03726_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__o31a_1
XFILLER_0_76_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18679_ _09945_ _09948_ memory.csr_read_data_out_reg\[0\] _09942_ VGND VGND VPWR
+ VPWR _03978_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20710_ _05809_ decode.id_ex_rs1_data_reg\[14\] _05798_ VGND VGND VPWR VPWR _05824_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21690_ net746 _06392_ _06393_ _06352_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_37_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20641_ _05627_ csr.io_mret_vector\[28\] _05603_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23360_ _07089_ _07780_ _07781_ _07785_ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__a211o_1
XFILLER_0_117_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20572_ _05541_ csr.io_mret_vector\[18\] _05602_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22311_ _06903_ _06678_ _06631_ _06905_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__a211o_1
XFILLER_0_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23291_ net223 _07706_ _07707_ _07721_ _07705_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__o311a_1
XFILLER_0_85_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25030_ _06331_ _08732_ _08733_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__nor3_1
XFILLER_0_147_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22242_ _06684_ _06836_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_200_Left_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22173_ net88 _06753_ _06767_ net224 VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21124_ _06054_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26981_ net195 _09862_ VGND VGND VPWR VPWR _09874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28720_ clknet_leaf_121_clock _01733_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[4\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25932_ net691 _09256_ _09257_ _09250_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__o211a_1
X_21055_ _06013_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20006_ _00549_ _05228_ _05230_ _05231_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__o22a_1
X_28651_ clknet_leaf_89_clock _01664_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_25863_ net488 _09213_ _09217_ _09209_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27602_ clknet_leaf_152_clock _00631_ VGND VGND VPWR VPWR execute.io_target_pc\[11\]
+ sky130_fd_sc_hd__dfxtp_4
X_24814_ _08107_ net1488 _08585_ VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__mux2_1
X_28582_ clknet_leaf_97_clock _01595_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25794_ net800 _09170_ _09177_ _09169_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27533_ clknet_leaf_156_clock _00562_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_97_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24745_ _08107_ net1541 _06283_ VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__mux2_1
X_21957_ net590 _06572_ _06580_ _06579_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_226_Right_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _05925_ _05933_ net39 VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__and3_1
X_24676_ _08521_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27464_ clknet_leaf_147_clock _00493_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[30\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21888_ csr._mcycle_T_2\[15\] _06521_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_867 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29203_ clknet_leaf_163_clock _02216_ VGND VGND VPWR VPWR fetch.btb.btbTable\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23627_ _07960_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__buf_4
XFILLER_0_166_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26415_ _09396_ _09545_ VGND VGND VPWR VPWR _09549_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20839_ net106 _05891_ _05887_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_13_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27395_ clknet_leaf_26_clock _00424_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29134_ clknet_leaf_76_clock _02147_ VGND VGND VPWR VPWR csr.mcycle\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14360_ _09970_ _10464_ VGND VGND VPWR VPWR _10467_ sky130_fd_sc_hd__nand2_1
X_23558_ net2779 _07917_ _07923_ _05805_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__o211a_1
X_26346_ _09402_ _09502_ VGND VGND VPWR VPWR _09509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22509_ _07100_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__buf_4
Xinput19 net378 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
X_29065_ clknet_leaf_220_clock _02078_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26277_ _09408_ _09459_ VGND VGND VPWR VPWR _09469_ sky130_fd_sc_hd__nand2_1
X_14291_ net2110 _10419_ _10425_ _10427_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__o211a_1
X_23489_ net22 _07875_ _07883_ _07879_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28016_ clknet_leaf_223_clock _01038_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16030_ decode.regfile.registers_23\[18\] _11088_ _11985_ _12008_ VGND VGND VPWR
+ VPWR _12009_ sky130_fd_sc_hd__o22a_1
X_25228_ _08843_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25159_ _08807_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17981_ _11022_ _12567_ _12586_ _12673_ decode.regfile.registers_16\[30\] VGND VGND
+ VPWR VPWR _03378_ sky130_fd_sc_hd__a32o_1
XFILLER_0_229_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19720_ _04995_ _04994_ _04454_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__o21ai_1
X_28918_ clknet_leaf_123_clock _01931_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_16932_ _11019_ _12504_ _12511_ decode.regfile.registers_8\[4\] _12892_ VGND VGND
+ VPWR VPWR _12893_ sky130_fd_sc_hd__o32a_1
XFILLER_0_229_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29898_ clknet_leaf_340_clock _02911_ VGND VGND VPWR VPWR decode.regfile.registers_20\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19651_ _04202_ _04207_ _04885_ _04206_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__o31ai_1
X_28849_ clknet_leaf_105_clock _01862_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_16863_ decode.regfile.registers_20\[3\] _11024_ _12553_ _12823_ _12824_ VGND VGND
+ VPWR VPWR _12825_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_221_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18602_ _03768_ _03769_ _03770_ _03896_ _03669_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__o41a_2
XFILLER_0_189_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15814_ decode.regfile.registers_18\[13\] _11225_ _11113_ _10988_ _10976_ VGND VGND
+ VPWR VPWR _11798_ sky130_fd_sc_hd__o2111a_1
X_19582_ _04209_ _03933_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16794_ _12513_ decode.regfile.registers_25\[1\] _12713_ _12757_ _12694_ VGND VGND
+ VPWR VPWR _12758_ sky130_fd_sc_hd__o221a_1
XFILLER_0_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18533_ execute.io_mem_memtoreg\[1\] execute.io_mem_memtoreg\[0\] execute.io_reg_pc\[25\]
+ _03831_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__o31a_1
X_15745_ _11154_ decode.regfile.registers_0\[11\] _11156_ _11730_ VGND VGND VPWR VPWR
+ _11731_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_38_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18464_ _03759_ net260 _03760_ _03762_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_155_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ decode.regfile.registers_14\[9\] _11207_ _11273_ decode.regfile.registers_15\[9\]
+ _11201_ VGND VGND VPWR VPWR _11664_ sky130_fd_sc_hd__a221o_1
XFILLER_0_213_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17415_ decode.regfile.registers_22\[15\] _13100_ _13364_ _13289_ VGND VGND VPWR
+ VPWR _13365_ sky130_fd_sc_hd__a211o_1
XFILLER_0_184_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14627_ _10587_ _10590_ _10600_ _10622_ _10669_ VGND VGND VPWR VPWR _10670_ sky130_fd_sc_hd__o41a_4
XFILLER_0_74_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18395_ decode.id_ex_ex_rs1_reg\[3\] _10194_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__or2b_4
XFILLER_0_172_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _13091_ _13176_ decode.regfile.registers_27\[13\] _13050_ VGND VGND VPWR
+ VPWR _13298_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14558_ decode.immGen._imm_T_24\[16\] VGND VGND VPWR VPWR _10601_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13509_ _09889_ VGND VGND VPWR VPWR _09890_ sky130_fd_sc_hd__buf_2
XFILLER_0_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17277_ _10610_ _12626_ _12629_ decode.regfile.registers_3\[12\] _13229_ VGND VGND
+ VPWR VPWR _13230_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14489_ net509 _10533_ _10540_ _10535_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19016_ _04296_ _04303_ _04305_ _04306_ _04314_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__o311a_1
X_16228_ _12133_ net485 _12169_ _12201_ _12132_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_228_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_228_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16159_ _11942_ decode.regfile.registers_30\[22\] _12095_ _12096_ _12097_ VGND VGND
+ VPWR VPWR _12134_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_110_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19918_ _05185_ _04215_ _05158_ _05159_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_177_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19849_ _03772_ net191 _03775_ _03794_ _03800_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_138_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22860_ _07326_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21811_ _06461_ csr.ie csr.pie _06032_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__o22a_1
XFILLER_0_223_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22791_ _07290_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_179_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24530_ _08446_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21742_ _06433_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_1271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24461_ _08089_ net1814 _08400_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21673_ _06377_ _06379_ _06381_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_43_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23412_ _07832_ _07833_ _07080_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__mux2_1
X_26200_ net198 VGND VGND VPWR VPWR _09420_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_43_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20624_ _05754_ _05756_ _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__a21oi_4
X_27180_ clknet_leaf_362_clock _00209_ VGND VGND VPWR VPWR decode.regfile.registers_27\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_24392_ net1510 VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26131_ _09930_ _10194_ _10150_ _08902_ VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__and4b_1
X_23343_ net85 net220 net221 _07728_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__nand4_1
Xclkbuf_5_24__f_clock clknet_2_3_0_clock VGND VGND VPWR VPWR clknet_5_24__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_20555_ _05541_ csr.io_mret_vector\[16\] _05602_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26062_ _09263_ VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__clkbuf_4
X_23274_ net80 _07536_ _07537_ _07704_ _07705_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__o311a_1
XFILLER_0_162_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20486_ csr.io_mret_vector\[7\] _05580_ _05581_ csr.mscratch\[7\] _05638_ VGND VGND
+ VPWR VPWR _05639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25013_ _08703_ _08716_ csr.mcycle\[7\] csr.mcycle\[8\] VGND VGND VPWR VPWR _08722_
+ sky130_fd_sc_hd__and4bb_1
X_22225_ _06740_ _06811_ _06815_ _06819_ net85 VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__a311o_1
XFILLER_0_131_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29821_ clknet_leaf_315_clock _02834_ VGND VGND VPWR VPWR decode.regfile.registers_18\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_22156_ _06750_ _06652_ _06629_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__a21o_1
XFILLER_0_219_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21107_ _05949_ _05945_ net2301 VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29752_ clknet_leaf_311_clock _02765_ VGND VGND VPWR VPWR decode.regfile.registers_15\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22087_ _06678_ _06681_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26964_ _09956_ VGND VGND VPWR VPWR _09865_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28703_ clknet_leaf_176_clock _01716_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21038_ _06004_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__clkbuf_1
X_25915_ net2413 _09242_ _09247_ _09235_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__o211a_1
X_29683_ clknet_leaf_283_clock _02696_ VGND VGND VPWR VPWR decode.regfile.registers_13\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26895_ net2267 _09822_ _09824_ _09825_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28634_ clknet_leaf_177_clock _01647_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_13860_ _10069_ _10164_ VGND VGND VPWR VPWR _10176_ sky130_fd_sc_hd__nand2_1
X_25846_ net2430 _09199_ _09207_ _09194_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28565_ clknet_leaf_205_clock _01578_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_22989_ fetch.bht.bhtTable_target_pc\[6\]\[6\] fetch.bht.bhtTable_target_pc\[7\]\[6\]
+ _07069_ VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__mux2_1
X_13791_ _10127_ VGND VGND VPWR VPWR _10128_ sky130_fd_sc_hd__clkbuf_8
X_25777_ _08925_ _09166_ VGND VGND VPWR VPWR _09168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15530_ _11050_ _11089_ decode.regfile.registers_25\[5\] _11494_ _11521_ VGND VGND
+ VPWR VPWR _11522_ sky130_fd_sc_hd__o32a_1
X_27516_ clknet_leaf_29_clock _00545_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dfxtp_1
X_24728_ _08548_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28496_ clknet_leaf_185_clock _01509_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27447_ clknet_leaf_149_clock _00476_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_15461_ _11219_ VGND VGND VPWR VPWR _11454_ sky130_fd_sc_hd__clkbuf_4
X_24659_ net1106 execute.io_target_pc\[18\] _08508_ VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17200_ decode.regfile.registers_12\[10\] _12489_ _11018_ _12540_ VGND VGND VPWR
+ VPWR _13155_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14412_ net543 _10490_ _10496_ _10494_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18180_ decode.immGen._imm_T_10\[4\] decode.immGen._imm_T_10\[2\] decode.immGen._imm_T_10\[1\]
+ decode.immGen._imm_T_10\[0\] VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15392_ decode.regfile.registers_16\[2\] _11359_ _11362_ _11386_ _11126_ VGND VGND
+ VPWR VPWR _11387_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27378_ clknet_leaf_10_clock _00407_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[19\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_189_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29117_ clknet_leaf_70_clock _02130_ VGND VGND VPWR VPWR csr.mcycle\[1\] sky130_fd_sc_hd__dfxtp_1
X_17131_ _11026_ VGND VGND VPWR VPWR _13088_ sky130_fd_sc_hd__clkbuf_4
X_26329_ net889 _09491_ _09498_ _09499_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__o211a_1
X_14343_ net891 _10447_ _10456_ _10453_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29048_ clknet_leaf_122_clock _02061_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14274_ _10147_ _10375_ VGND VGND VPWR VPWR _10416_ sky130_fd_sc_hd__nand2_1
X_17062_ _12522_ _12616_ _10608_ VGND VGND VPWR VPWR _13020_ sky130_fd_sc_hd__and3_2
XFILLER_0_208_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16013_ decode.regfile.registers_2\[18\] _11295_ VGND VGND VPWR VPWR _11992_ sky130_fd_sc_hd__nor2_1
XFILLER_0_208_1299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_115_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1085 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_223_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _12561_ _03360_ _03361_ _12906_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19703_ _04503_ _03888_ _04189_ _04505_ _03894_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__a2111o_1
X_16915_ _12583_ VGND VGND VPWR VPWR _12876_ sky130_fd_sc_hd__clkbuf_4
X_17895_ _02986_ decode.regfile.registers_26\[27\] _13002_ _13484_ _02987_ VGND VGND
+ VPWR VPWR _03295_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19634_ _03924_ _04889_ _04207_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__and3_1
X_16846_ _12494_ decode.regfile.registers_24\[2\] _12691_ VGND VGND VPWR VPWR _12809_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19565_ _04847_ _04252_ _04251_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16777_ _12726_ _12739_ _12740_ VGND VGND VPWR VPWR _12741_ sky130_fd_sc_hd__a21o_1
XFILLER_0_215_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13989_ net2333 _10243_ _10252_ _10249_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_124_Left_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18516_ _03768_ _03769_ _03770_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__nor3_2
X_15728_ decode.regfile.registers_22\[10\] _11096_ _11713_ _11714_ _11232_ VGND VGND
+ VPWR VPWR _11715_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19496_ _04117_ _04115_ _04107_ _04103_ _04100_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__o32a_1
XFILLER_0_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18447_ net315 VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_174_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15659_ _11493_ decode.regfile.registers_24\[9\] VGND VGND VPWR VPWR _11647_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18378_ decode.io_wb_rd\[1\] decode.id_ex_ex_rs1_reg\[1\] VGND VGND VPWR VPWR _03677_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_111_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17329_ decode.regfile.registers_14\[13\] _10604_ _10618_ _12772_ VGND VGND VPWR
+ VPWR _13281_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20340_ _05505_ _05506_ _05418_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Left_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20271_ _05417_ _05294_ _05453_ _05454_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_73_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22010_ csr.mscratch\[27\] _06601_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2502 decode.regfile.registers_9\[30\] VGND VGND VPWR VPWR net2729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2513 decode.regfile.registers_7\[28\] VGND VGND VPWR VPWR net2740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2524 fetch.btb.btbTable\[0\]\[1\] VGND VGND VPWR VPWR net2751 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2535 csr._minstret_T_3\[63\] VGND VGND VPWR VPWR net2762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2546 net86 VGND VGND VPWR VPWR net2773 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1801 execute.io_mem_rd\[4\] VGND VGND VPWR VPWR net2028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1812 fetch.bht.bhtTable_tag\[7\]\[17\] VGND VGND VPWR VPWR net2039 sky130_fd_sc_hd__dlygate4sd3_1
X_23961_ net1501 execute.io_target_pc\[2\] _07983_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__mux2_1
Xhold2557 decode.regfile.registers_30\[21\] VGND VGND VPWR VPWR net2784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 fetch.bht.bhtTable_target_pc\[15\]\[23\] VGND VGND VPWR VPWR net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 csr._minstret_T_3\[55\] VGND VGND VPWR VPWR net2795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1834 fetch.bht.bhtTable_target_pc\[6\]\[5\] VGND VGND VPWR VPWR net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_341_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_341_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_32_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1845 decode.regfile.registers_2\[13\] VGND VGND VPWR VPWR net2072 sky130_fd_sc_hd__dlygate4sd3_1
X_25700_ net1263 _09111_ _09123_ _09115_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__o211a_1
X_22912_ net225 _06698_ _06916_ _06894_ _07362_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_32_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23892_ _08115_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__clkbuf_1
Xhold1856 fetch.bht.bhtTable_tag\[13\]\[1\] VGND VGND VPWR VPWR net2083 sky130_fd_sc_hd__dlygate4sd3_1
X_26680_ _10130_ VGND VGND VPWR VPWR _09701_ sky130_fd_sc_hd__buf_2
Xhold1867 fetch.bht.bhtTable_tag\[0\]\[20\] VGND VGND VPWR VPWR net2094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1878 decode.regfile.registers_7\[27\] VGND VGND VPWR VPWR net2105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_142_Left_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1889 decode.regfile.registers_21\[9\] VGND VGND VPWR VPWR net2116 sky130_fd_sc_hd__dlygate4sd3_1
X_22843_ _07317_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__clkbuf_1
X_25631_ _08931_ _09079_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28350_ clknet_leaf_195_clock _01363_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22774_ _07280_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__clkbuf_1
X_25562_ _08937_ _09036_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_356_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_356_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_211_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27301_ clknet_leaf_13_clock _00330_ VGND VGND VPWR VPWR decode.regfile.registers_31\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_24513_ _08437_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21725_ _10576_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28281_ clknet_leaf_85_clock _01303_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_25493_ _08990_ VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27232_ clknet_leaf_2_clock _00261_ VGND VGND VPWR VPWR decode.regfile.registers_29\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_24444_ _08401_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__clkbuf_1
X_21656_ _05691_ csr.minstret\[16\] _06366_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20607_ _03737_ _03718_ csr._csr_read_data_T_8\[23\] VGND VGND VPWR VPWR _05744_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_19_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24375_ _08364_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27163_ clknet_leaf_360_clock _00192_ VGND VGND VPWR VPWR decode.regfile.registers_27\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_21587_ csr.io_csr_write_address\[0\] _06315_ csr.io_csr_write_address\[1\] VGND
+ VGND VPWR VPWR _06316_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_105_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_151_Left_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23326_ _07110_ _07753_ VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__and2b_1
X_26114_ _08960_ _09353_ VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__nand2_1
X_20538_ _05681_ _05684_ _05414_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27094_ clknet_leaf_329_clock _00123_ VGND VGND VPWR VPWR decode.regfile.registers_25\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23257_ net79 net224 _07636_ net80 VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__a31o_1
X_26045_ _08966_ _09310_ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__nand2_1
X_20469_ csr._minstret_T_3\[37\] _05616_ _05622_ csr._csr_read_data_T_8\[5\] _05623_
+ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22208_ fetch.bht.bhtTable_tag\[8\]\[24\] fetch.bht.bhtTable_tag\[9\]\[24\] fetch.bht.bhtTable_tag\[10\]\[24\]
+ fetch.bht.bhtTable_tag\[11\]\[24\] _06645_ _06651_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__mux4_1
X_23188_ fetch.bht.bhtTable_target_pc\[4\]\[17\] fetch.bht.bhtTable_target_pc\[5\]\[17\]
+ fetch.bht.bhtTable_target_pc\[6\]\[17\] fetch.bht.bhtTable_target_pc\[7\]\[17\]
+ _07384_ _07386_ VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29804_ clknet_leaf_295_clock _02817_ VGND VGND VPWR VPWR decode.regfile.registers_17\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_22139_ fetch.bht.bhtTable_tag\[2\]\[4\] fetch.bht.bhtTable_tag\[3\]\[4\] _06706_
+ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__mux2_1
X_27996_ clknet_leaf_206_clock _01018_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_29735_ clknet_leaf_285_clock _02748_ VGND VGND VPWR VPWR decode.regfile.registers_15\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14961_ _10974_ _10986_ VGND VGND VPWR VPWR _10987_ sky130_fd_sc_hd__and2_1
X_26947_ net643 _09853_ _09855_ _09852_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_309_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_309_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_215_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_160_Left_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16700_ decode.regfile.registers_13\[0\] _12586_ _12589_ _12660_ _12664_ VGND VGND
+ VPWR VPWR _12665_ sky130_fd_sc_hd__a311o_1
XFILLER_0_57_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13912_ net962 _10199_ _10207_ _10206_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__o211a_1
X_29666_ clknet_leaf_287_clock _02679_ VGND VGND VPWR VPWR decode.regfile.registers_13\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_17680_ decode.regfile.registers_8\[22\] _12843_ _12606_ VGND VGND VPWR VPWR _03085_
+ sky130_fd_sc_hd__a21oi_1
X_14892_ _10928_ VGND VGND VPWR VPWR _10929_ sky130_fd_sc_hd__clkbuf_4
X_26878_ net2120 _09809_ _09815_ _09812_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28617_ clknet_leaf_88_clock _01630_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16631_ decode.regfile.registers_11\[0\] _12595_ _12583_ _12551_ VGND VGND VPWR VPWR
+ _12596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13843_ net492 _10153_ _10166_ _10162_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__o211a_1
X_25829_ _10373_ _10150_ _08902_ _09935_ VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__and4_1
X_29597_ clknet_leaf_270_clock _02610_ VGND VGND VPWR VPWR decode.regfile.registers_11\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19350_ _04130_ _04131_ _04640_ _04454_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__o31a_1
X_28548_ clknet_leaf_188_clock _01561_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_16562_ _12526_ VGND VGND VPWR VPWR _12527_ sky130_fd_sc_hd__buf_2
X_13774_ net2417 _10083_ _10113_ _10077_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18301_ _03615_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__clkbuf_1
X_15513_ decode.regfile.registers_5\[5\] _11192_ _11139_ _11502_ _11504_ VGND VGND
+ VPWR VPWR _11505_ sky130_fd_sc_hd__a32o_1
XFILLER_0_214_1281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19281_ _04294_ _04571_ _04574_ _04360_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28479_ clknet_leaf_238_clock _01492_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16493_ decode.regfile.registers_2\[31\] _11296_ _11297_ _11121_ _12458_ VGND VGND
+ VPWR VPWR _12459_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_216_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_216_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18232_ csr.mcycle\[29\] _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__nand2_1
X_15444_ _11236_ _11433_ _11434_ _11437_ VGND VGND VPWR VPWR _11438_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_807 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18163_ _03509_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_212_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15375_ _11117_ _11137_ _11157_ decode.regfile.registers_0\[2\] VGND VGND VPWR VPWR
+ _11370_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17114_ decode.regfile.registers_14\[8\] _12664_ _13069_ _13070_ _12585_ VGND VGND
+ VPWR VPWR _13071_ sky130_fd_sc_hd__a221o_1
XFILLER_0_170_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14326_ _10418_ VGND VGND VPWR VPWR _10447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18094_ _03469_ _03467_ _03465_ net2195 VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold408 decode.regfile.registers_30\[28\] VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 _08651_ VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__dlygate4sd3_1
X_17045_ _12968_ _13000_ _13001_ _13003_ VGND VGND VPWR VPWR _13004_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_225_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14257_ _10102_ _10400_ VGND VGND VPWR VPWR _10407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14188_ net1862 _10359_ _10366_ _10357_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18996_ _04294_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1108 fetch.bht.bhtTable_target_pc\[0\]\[8\] VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__dlygate4sd3_1
X_17947_ decode.regfile.registers_3\[29\] _12639_ _10609_ _12625_ VGND VGND VPWR VPWR
+ _03345_ sky130_fd_sc_hd__o2bb2a_1
Xhold1119 _08205_ VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_163_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17878_ _12602_ decode.regfile.registers_9\[27\] _12652_ _03277_ VGND VGND VPWR VPWR
+ _03278_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19617_ _04791_ _04897_ _04272_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__mux2_1
X_16829_ _12791_ VGND VGND VPWR VPWR _12792_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_176_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19548_ _04827_ _04781_ _04811_ _04830_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19479_ _04103_ _04100_ _04359_ _04504_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__a211o_1
XINSDIODE1_350 _03580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21510_ _06272_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_361 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_372 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_383 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22490_ _07084_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21441_ _06132_ net1150 _06230_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24160_ _08253_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21372_ _06198_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_131_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23111_ net280 _07548_ _07551_ _03592_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__o211ai_1
X_20323_ _10864_ _10786_ decode.id_ex_pc_reg\[24\] _05482_ VGND VGND VPWR VPWR _05494_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_4_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24091_ net913 execute.io_target_pc\[1\] _06450_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__mux2_1
Xhold920 fetch.bht.bhtTable_tag\[12\]\[23\] VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold931 csr._mcycle_T_2\[31\] VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_9_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23042_ _06025_ _07484_ _07345_ _07486_ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__a31o_1
Xhold942 decode.regfile.registers_7\[1\] VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_222_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold953 fetch.bht.bhtTable_target_pc\[1\]\[19\] VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__dlygate4sd3_1
X_20254_ decode.id_ex_rdsel_reg _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__nor2_1
Xhold964 fetch.bht.bhtTable_tag\[13\]\[20\] VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold975 fetch.bht.bhtTable_target_pc\[12\]\[13\] VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold986 fetch.bht.bhtTable_target_pc\[8\]\[14\] VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold997 fetch.bht.bhtTable_target_pc\[8\]\[10\] VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27850_ clknet_leaf_323_clock _00879_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20185_ decode.id_ex_imm_reg\[27\] _10854_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__or2_1
Xhold2310 decode.regfile.registers_12\[18\] VGND VGND VPWR VPWR net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2321 csr._mcycle_T_3\[61\] VGND VGND VPWR VPWR net2548 sky130_fd_sc_hd__dlygate4sd3_1
X_26801_ net894 _09766_ _09770_ _09771_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_280_clock clknet_5_21__leaf_clock VGND VGND VPWR VPWR clknet_leaf_280_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2332 decode.regfile.registers_26\[19\] VGND VGND VPWR VPWR net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_27781_ clknet_leaf_334_clock _00810_ VGND VGND VPWR VPWR memory.io_wb_readdata\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2343 decode.regfile.registers_7\[20\] VGND VGND VPWR VPWR net2570 sky130_fd_sc_hd__dlygate4sd3_1
X_24993_ _08701_ _03557_ _06327_ _08708_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_192_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2354 csr._mcycle_T_2\[2\] VGND VGND VPWR VPWR net2581 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1620 execute.csr_write_address_out_reg\[6\] VGND VGND VPWR VPWR net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2365 decode.regfile.registers_24\[23\] VGND VGND VPWR VPWR net2592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29520_ clknet_leaf_265_clock _02533_ VGND VGND VPWR VPWR decode.regfile.registers_8\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1631 fetch.bht.bhtTable_tag\[6\]\[22\] VGND VGND VPWR VPWR net1858 sky130_fd_sc_hd__dlygate4sd3_1
X_26732_ net715 _09723_ _09731_ _09730_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__o211a_1
Xhold2376 decode.regfile.registers_8\[31\] VGND VGND VPWR VPWR net2603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2387 fetch.bht.bhtTable_target_pc\[15\]\[6\] VGND VGND VPWR VPWR net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1642 fetch.bht.bhtTable_tag\[10\]\[18\] VGND VGND VPWR VPWR net1869 sky130_fd_sc_hd__dlygate4sd3_1
X_23944_ _08142_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__clkbuf_1
Xhold1653 fetch.bht.bhtTable_target_pc\[14\]\[17\] VGND VGND VPWR VPWR net1880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2398 _01249_ VGND VGND VPWR VPWR net2625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1664 decode.regfile.registers_22\[0\] VGND VGND VPWR VPWR net1891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1675 fetch.bht.bhtTable_tag\[14\]\[12\] VGND VGND VPWR VPWR net1902 sky130_fd_sc_hd__dlygate4sd3_1
X_29451_ clknet_leaf_254_clock _02464_ VGND VGND VPWR VPWR decode.regfile.registers_6\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1686 csr.mscratch\[2\] VGND VGND VPWR VPWR net1913 sky130_fd_sc_hd__dlygate4sd3_1
X_26663_ net793 _09679_ _09691_ _09688_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23875_ _08104_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__clkbuf_1
Xhold1697 decode.regfile.registers_16\[13\] VGND VGND VPWR VPWR net1924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_295_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_295_clock
+ sky130_fd_sc_hd__clkbuf_8
X_28402_ clknet_leaf_142_clock _01415_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_4
X_25614_ net811 _09068_ _09073_ _09074_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__o211a_1
X_22826_ net1003 _10760_ _07308_ VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29382_ clknet_leaf_257_clock _02395_ VGND VGND VPWR VPWR decode.regfile.registers_4\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26594_ _09424_ _09645_ VGND VGND VPWR VPWR _09652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28333_ clknet_leaf_222_clock _01346_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25545_ net622 _09024_ _09034_ _09033_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__o211a_1
X_22757_ _07271_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21708_ csr.minstret\[19\] csr.minstret\[26\] csr.io_inst_retired _06408_ VGND VGND
+ VPWR VPWR _06409_ sky130_fd_sc_hd__and4_1
X_28264_ clknet_leaf_64_clock _01286_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22688_ net2604 _07222_ _07231_ _07221_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25476_ net946 _08979_ _08994_ _08991_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27215_ clknet_leaf_352_clock _00244_ VGND VGND VPWR VPWR decode.regfile.registers_29\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_229_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24427_ _08392_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21639_ csr._mcycle_T_2\[12\] _06325_ _06338_ _06355_ csr.minstret\[12\] VGND VGND
+ VPWR VPWR _06356_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_212_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28195_ clknet_leaf_85_clock _01217_ VGND VGND VPWR VPWR csr.io_mret_vector\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_229_Left_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15160_ _11108_ VGND VGND VPWR VPWR _11157_ sky130_fd_sc_hd__clkbuf_4
X_27146_ clknet_leaf_358_clock _00175_ VGND VGND VPWR VPWR decode.regfile.registers_26\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_24358_ _08355_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_233_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_233_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14111_ net2651 _10315_ _10322_ _10317_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__o211a_1
X_23309_ _07734_ _07735_ _07736_ _07737_ _07371_ _07127_ VGND VGND VPWR VPWR _07738_
+ sky130_fd_sc_hd__mux4_2
X_15091_ _11087_ VGND VGND VPWR VPWR _11088_ sky130_fd_sc_hd__clkbuf_4
X_24289_ _08051_ net2296 _06210_ VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27077_ clknet_leaf_347_clock _00106_ VGND VGND VPWR VPWR decode.regfile.registers_24\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14042_ _10136_ _10242_ VGND VGND VPWR VPWR _10282_ sky130_fd_sc_hd__nand2_1
X_26028_ net2052 _09300_ _09312_ _09305_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18850_ _04145_ net355 _03687_ decode.id_ex_rs1_data_reg\[11\] _04148_ VGND VGND
+ VPWR VPWR _04149_ sky130_fd_sc_hd__o221a_2
XFILLER_0_140_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_248_clock clknet_5_19__leaf_clock VGND VGND VPWR VPWR clknet_leaf_248_clock
+ sky130_fd_sc_hd__clkbuf_8
X_17801_ _12595_ _03201_ _03202_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__o21ai_1
X_18781_ _03817_ _04079_ _03774_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__a21oi_2
X_27979_ clknet_leaf_200_clock _01001_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_15993_ _11060_ _11098_ _11454_ decode.regfile.registers_20\[17\] _11972_ VGND VGND
+ VPWR VPWR _11973_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_175_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17732_ decode.regfile.registers_22\[23\] _13100_ _03135_ _13289_ VGND VGND VPWR
+ VPWR _03136_ sky130_fd_sc_hd__a211o_1
X_29718_ clknet_leaf_283_clock _02731_ VGND VGND VPWR VPWR decode.regfile.registers_14\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14944_ net66 _10972_ VGND VGND VPWR VPWR _10973_ sky130_fd_sc_hd__nor2_8
XFILLER_0_215_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17663_ _02990_ _03068_ decode.regfile.registers_27\[21\] _13487_ VGND VGND VPWR
+ VPWR _03069_ sky130_fd_sc_hd__or4_1
X_29649_ clknet_leaf_279_clock _02662_ VGND VGND VPWR VPWR decode.regfile.registers_12\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14875_ _10912_ _10913_ _10916_ decode.immGen._imm_T_10\[0\] VGND VGND VPWR VPWR
+ _10917_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_218_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19402_ _04647_ _04690_ _04324_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_218_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16614_ _12578_ VGND VGND VPWR VPWR _12579_ sky130_fd_sc_hd__clkbuf_4
X_13826_ _09970_ _10154_ VGND VGND VPWR VPWR _10157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17594_ decode.regfile.registers_1\[20\] decode.regfile.registers_0\[20\] _12631_
+ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19333_ _04623_ _04486_ _04249_ _04624_ _04541_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__o221a_1
XFILLER_0_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16545_ _12509_ VGND VGND VPWR VPWR _12510_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_214_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13757_ _10003_ _10021_ memory.io_wb_readdata\[23\] VGND VGND VPWR VPWR _10099_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_171_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19264_ _04034_ _04056_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16476_ _10992_ _11244_ _11261_ _12442_ VGND VGND VPWR VPWR _12443_ sky130_fd_sc_hd__a31o_1
X_13688_ memory.csr_read_data_out_reg\[12\] _09989_ _10039_ _10040_ VGND VGND VPWR
+ VPWR _10041_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_31_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18215_ _10577_ _03546_ _03550_ _03551_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__nor4_1
XFILLER_0_26_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15427_ _11419_ _11420_ _11186_ VGND VGND VPWR VPWR _11421_ sky130_fd_sc_hd__a21oi_1
X_19195_ _04490_ _04346_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_208_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18146_ _03502_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15358_ _10956_ decode.regfile.registers_22\[2\] _11093_ _11264_ _10989_ VGND VGND
+ VPWR VPWR _11353_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_41_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold205 _10716_ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
Xwire180 net181 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14309_ net671 _10434_ _10437_ _10427_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_169_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18077_ _10944_ _10941_ _10581_ _10946_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_895 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold216 decode.regfile.registers_31\[19\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ _11284_ VGND VGND VPWR VPWR _11285_ sky130_fd_sc_hd__buf_4
Xhold227 decode.regfile.registers_30\[19\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 net113 VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17028_ decode.regfile.registers_16\[6\] _12673_ _12901_ VGND VGND VPWR VPWR _12987_
+ sky130_fd_sc_hd__a21oi_1
Xhold249 decode.regfile.registers_30\[29\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18979_ _04275_ _04276_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21990_ csr._mcycle_T_2\[18\] _06587_ _06598_ _06592_ VGND VGND VPWR VPWR _01238_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_68_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20941_ _05949_ _05945_ net55 VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_124_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23660_ _07978_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__clkbuf_1
X_20872_ net123 _05903_ _05911_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22611_ _07184_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23591_ _07940_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22542_ _03580_ _07135_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__nor2_1
X_25330_ _08891_ net2693 VGND VGND VPWR VPWR _08896_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_27_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_180 execute.io_reg_pc\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_191 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25261_ _08860_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__clkbuf_1
X_22473_ _07067_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__buf_6
XFILLER_0_161_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27000_ clknet_leaf_337_clock _00029_ VGND VGND VPWR VPWR decode.regfile.registers_22\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24212_ _08280_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__clkbuf_1
X_21424_ _06115_ net1683 _06219_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25192_ _10572_ fetch.btb.btbTable\[4\]\[1\] _08824_ VGND VGND VPWR VPWR _08825_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24143_ net863 execute.io_target_pc\[26\] _06427_ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__mux2_1
X_21355_ _06103_ net1242 _06188_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20306_ _05411_ _05349_ _05479_ _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_114_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24074_ _08209_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__clkbuf_1
X_28951_ clknet_leaf_124_clock _01964_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold750 fetch.bht.bhtTable_target_pc\[12\]\[26\] VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21286_ _06150_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_1320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold761 fetch.bht.bhtTable_target_pc\[8\]\[26\] VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold772 fetch.bht.bhtTable_target_pc\[3\]\[5\] VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__dlygate4sd3_1
X_27902_ clknet_leaf_81_clock _00931_ VGND VGND VPWR VPWR csr._mcycle_T_2\[23\] sky130_fd_sc_hd__dfxtp_1
X_23025_ net96 _07343_ _07344_ _07470_ _06566_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_57_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold783 fetch.bht.bhtTable_tag\[0\]\[3\] VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__dlygate4sd3_1
X_20237_ _10834_ _10747_ decode.id_ex_pc_reg\[4\] VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_229_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28882_ clknet_leaf_108_clock _01895_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold794 fetch.bht.bhtTable_tag\[0\]\[19\] VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27833_ clknet_leaf_324_clock _00862_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20168_ decode.id_ex_imm_reg\[22\] _10864_ _10786_ decode.id_ex_imm_reg\[23\] VGND
+ VGND VPWR VPWR _05371_ sky130_fd_sc_hd__a22o_1
Xhold2140 decode.regfile.registers_18\[26\] VGND VGND VPWR VPWR net2367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2151 decode.regfile.registers_10\[23\] VGND VGND VPWR VPWR net2378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2162 decode.regfile.registers_8\[26\] VGND VGND VPWR VPWR net2389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2173 decode.regfile.registers_11\[21\] VGND VGND VPWR VPWR net2400 sky130_fd_sc_hd__dlygate4sd3_1
X_27764_ clknet_leaf_317_clock _00793_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_20099_ _05296_ _05305_ _05311_ _05302_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__a31o_1
X_24976_ csr._mcycle_T_3\[61\] csr._mcycle_T_3\[60\] csr._mcycle_T_3\[59\] _08693_
+ _03579_ VGND VGND VPWR VPWR _08697_ sky130_fd_sc_hd__a41o_1
Xhold2184 decode.regfile.registers_25\[23\] VGND VGND VPWR VPWR net2411 sky130_fd_sc_hd__dlygate4sd3_1
X_29503_ clknet_leaf_252_clock _02516_ VGND VGND VPWR VPWR decode.regfile.registers_8\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2195 decode.regfile.registers_7\[2\] VGND VGND VPWR VPWR net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1450 decode.regfile.registers_4\[6\] VGND VGND VPWR VPWR net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 fetch.bht.bhtTable_tag\[9\]\[9\] VGND VGND VPWR VPWR net1688 sky130_fd_sc_hd__dlygate4sd3_1
X_26715_ _09392_ _09720_ VGND VGND VPWR VPWR _09722_ sky130_fd_sc_hd__nand2_1
X_23927_ net834 _08085_ _08130_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__mux2_1
Xhold1472 decode.regfile.registers_15\[16\] VGND VGND VPWR VPWR net1699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27695_ clknet_leaf_23_clock _00724_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1483 decode.regfile.registers_5\[3\] VGND VGND VPWR VPWR net1710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1494 fetch.bht.bhtTable_target_pc\[7\]\[17\] VGND VGND VPWR VPWR net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29434_ clknet_leaf_255_clock _02447_ VGND VGND VPWR VPWR decode.regfile.registers_6\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14660_ execute.io_target_pc\[0\] VGND VGND VPWR VPWR _10703_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26646_ _09400_ _09676_ VGND VGND VPWR VPWR _09682_ sky130_fd_sc_hd__nand2_1
X_23858_ execute.io_target_pc\[21\] VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__buf_2
XFILLER_0_197_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13611_ _09939_ memory.io_wb_aluresult\[3\] _09961_ memory.io_wb_reg_pc\[3\] _09960_
+ VGND VGND VPWR VPWR _09973_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22809_ net887 csr.io_mem_pc\[18\] _07297_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__mux2_1
X_29365_ clknet_leaf_227_clock _02378_ VGND VGND VPWR VPWR decode.regfile.registers_3\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26577_ _09406_ _09632_ VGND VGND VPWR VPWR _09642_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14591_ _10633_ decode.id_ex_ex_rd_reg\[1\] VGND VGND VPWR VPWR _10634_ sky130_fd_sc_hd__nand2_1
X_23789_ _06151_ net1707 _08041_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28316_ clknet_leaf_203_clock _01329_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16330_ decode.regfile.registers_23\[26\] _11232_ _11074_ VGND VGND VPWR VPWR _12301_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13542_ _09914_ _09894_ _09916_ net396 VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__a31o_1
X_25528_ _09023_ VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29296_ clknet_leaf_224_clock _02309_ VGND VGND VPWR VPWR decode.regfile.registers_1\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28247_ clknet_leaf_78_clock _01269_ VGND VGND VPWR VPWR csr._minstret_T_3\[47\]
+ sky130_fd_sc_hd__dfxtp_2
X_16261_ _11756_ decode.regfile.registers_28\[24\] _11871_ _11681_ _11448_ VGND VGND
+ VPWR VPWR _12234_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_129_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25459_ net1434 _08979_ _08984_ _08972_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18000_ decode.regfile.registers_19\[30\] _12678_ _03377_ _03396_ _12906_ VGND VGND
+ VPWR VPWR _03397_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_172_clock clknet_5_24__leaf_clock VGND VGND VPWR VPWR clknet_leaf_172_clock
+ sky130_fd_sc_hd__clkbuf_8
X_15212_ decode.regfile.registers_15\[0\] _11036_ _11205_ _11208_ decode.regfile.registers_14\[0\]
+ VGND VGND VPWR VPWR _11209_ sky130_fd_sc_hd__a32o_1
XFILLER_0_168_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28178_ clknet_leaf_60_clock _01200_ VGND VGND VPWR VPWR csr.io_mret_vector\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16192_ _11489_ decode.regfile.registers_28\[22\] decode.regfile.registers_29\[22\]
+ _11255_ VGND VGND VPWR VPWR _12167_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15143_ _11055_ _10627_ decode.immGen._imm_T_24\[11\] VGND VGND VPWR VPWR _11140_
+ sky130_fd_sc_hd__and3_1
X_27129_ clknet_leaf_356_clock _00158_ VGND VGND VPWR VPWR decode.regfile.registers_26\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19951_ decode.id_ex_pc_reg\[0\] _03627_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15074_ _11070_ VGND VGND VPWR VPWR _11071_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_187_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_187_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_207_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14025_ _10092_ _10268_ VGND VGND VPWR VPWR _10273_ sky130_fd_sc_hd__nand2_1
X_18902_ _04199_ _04200_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_207_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19882_ _05145_ _05148_ _05151_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_208_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18833_ _04130_ _04131_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_110_clock clknet_5_11__leaf_clock VGND VGND VPWR VPWR clknet_leaf_110_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_199_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18764_ _03715_ _03725_ _04059_ _03727_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__o31a_1
X_15976_ _11129_ _11147_ _11954_ _11955_ VGND VGND VPWR VPWR _11956_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_101_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17715_ decode.regfile.registers_1\[23\] net215 _12530_ VGND VGND VPWR VPWR _03119_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14927_ _10955_ VGND VGND VPWR VPWR _10956_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18695_ _03993_ _03657_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_222_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17646_ _12659_ _03049_ _03050_ _03051_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_63_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14858_ decode.id_ex_pc_reg\[18\] _10870_ _10874_ _10900_ VGND VGND VPWR VPWR _10901_
+ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_63_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_125_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_125_clock
+ sky130_fd_sc_hd__clkbuf_8
X_13809_ net2308 _09951_ _10143_ _10132_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__o211a_1
XFILLER_0_212_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17577_ _13407_ decode.regfile.registers_25\[19\] _13482_ _13294_ VGND VGND VPWR
+ VPWR _02985_ sky130_fd_sc_hd__or4_1
X_14789_ decode.id_ex_pc_reg\[1\] csr.io_mem_pc\[1\] VGND VGND VPWR VPWR _10832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19316_ _04330_ _04482_ _04607_ _04243_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16528_ _12492_ VGND VGND VPWR VPWR _12493_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19247_ _04259_ _04342_ _04541_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16459_ _11043_ decode.regfile.registers_4\[30\] _11503_ _10629_ _11083_ VGND VGND
+ VPWR VPWR _12426_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_186_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19178_ _04472_ _04473_ net242 VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18129_ _03492_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21140_ _06063_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21071_ execute.csr_read_data_out_reg\[24\] _06014_ _03583_ VGND VGND VPWR VPWR _06022_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_111_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20022_ _05245_ _05239_ _00551_ _05227_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_207_Right_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24830_ _08602_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24761_ _08566_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21973_ csr._mcycle_T_2\[10\] _06587_ _06589_ _06579_ VGND VGND VPWR VPWR _01230_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_87_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer20 net246 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__buf_1
XFILLER_0_193_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26500_ _09404_ _09589_ VGND VGND VPWR VPWR _09598_ sky130_fd_sc_hd__nand2_1
Xrebuffer31 _03763_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_1
X_23712_ net1178 _10800_ _08003_ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__mux2_1
Xrebuffer42 _10762_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
X_27480_ clknet_leaf_52_clock _00509_ VGND VGND VPWR VPWR decode.exception_out_reg
+ sky130_fd_sc_hd__dfxtp_1
X_20924_ _05942_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer53 _03724_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd1_1
X_24692_ _08529_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer64 net290 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer75 _00568_ VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dlymetal6s4s_1
XFILLER_0_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer86 net309 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_1
X_26431_ net2186 _09548_ _09557_ _09553_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23643_ _07969_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__clkbuf_1
X_20855_ net114 _05903_ _05899_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__and3_1
Xrebuffer97 _11069_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29150_ clknet_leaf_223_clock _02163_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26362_ _09490_ VGND VGND VPWR VPWR _09518_ sky130_fd_sc_hd__buf_2
XFILLER_0_193_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23574_ _06105_ net2017 _07930_ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20786_ _03590_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28101_ clknet_leaf_74_clock net2677 VGND VGND VPWR VPWR csr.minstret\[6\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_46_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25313_ _08880_ decode.regfile.registers_0\[18\] VGND VGND VPWR VPWR _08887_ sky130_fd_sc_hd__and2_1
X_22525_ _07067_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__clkbuf_8
X_29081_ clknet_leaf_169_clock _02094_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26293_ net2647 _09475_ _09478_ _09471_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28032_ clknet_leaf_187_clock _01054_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer110 net336 VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25244_ _08083_ net2111 _08848_ VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__mux2_1
Xrebuffer121 net346 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22456_ _06754_ fetch.btb.btbTable\[8\]\[1\] fetch.bht.bhtTable_valid\[8\] VGND VGND
+ VPWR VPWR _07051_ sky130_fd_sc_hd__and3b_1
XFILLER_0_150_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21407_ _09900_ _10556_ _10557_ _09916_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__or4bb_4
X_22387_ fetch.bht.bhtTable_tag\[0\]\[9\] fetch.bht.bhtTable_tag\[1\]\[9\] fetch.bht.bhtTable_tag\[2\]\[9\]
+ fetch.bht.bhtTable_tag\[3\]\[9\] _06754_ _06622_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__mux4_1
X_25175_ net416 _08816_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24126_ net1437 VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__clkbuf_1
X_21338_ net808 _10760_ _06179_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1091 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21269_ net1052 _06138_ _06120_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__mux2_1
X_24057_ net1322 execute.io_target_pc\[16\] _08198_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__mux2_1
X_28934_ clknet_leaf_97_clock _01947_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold580 _01234_ VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold591 decode.regfile.registers_1\[21\] VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd3_1
X_23008_ fetch.bht.bhtTable_target_pc\[0\]\[7\] fetch.bht.bhtTable_target_pc\[1\]\[7\]
+ fetch.bht.bhtTable_target_pc\[2\]\[7\] fetch.bht.bhtTable_target_pc\[3\]\[7\] _07407_
+ _07072_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__mux4_1
X_28865_ clknet_leaf_175_clock _01878_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_202_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ decode.regfile.registers_11\[13\] _11070_ _11470_ _11800_ _11813_ VGND VGND
+ VPWR VPWR _11814_ sky130_fd_sc_hd__a32o_1
X_27816_ clknet_leaf_323_clock _00845_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_202_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28796_ clknet_leaf_181_clock _01809_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_204_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15761_ decode.regfile.registers_18\[11\] _11059_ _11149_ _11406_ _11746_ VGND VGND
+ VPWR VPWR _11747_ sky130_fd_sc_hd__o311a_1
X_27747_ clknet_leaf_35_clock _00776_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24959_ csr._mcycle_T_3\[55\] csr._mcycle_T_3\[54\] csr._mcycle_T_3\[53\] _08682_
+ _03579_ VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__a41o_1
Xclkbuf_leaf_42_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_42_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold1280 fetch.bht.bhtTable_target_pc\[5\]\[28\] VGND VGND VPWR VPWR net1507 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17500_ _13215_ decode.regfile.registers_28\[17\] _13093_ VGND VGND VPWR VPWR _13448_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_194_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1291 fetch.bht.bhtTable_target_pc\[3\]\[7\] VGND VGND VPWR VPWR net1518 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ _10702_ execute.io_target_pc\[14\] _10715_ _10740_ _10754_ VGND VGND VPWR
+ VPWR _10755_ sky130_fd_sc_hd__a2111oi_2
X_18480_ execute.io_reg_pc\[29\] _03777_ _03666_ net121 _03778_ VGND VGND VPWR VPWR
+ _03779_ sky130_fd_sc_hd__o221a_1
X_15692_ _11679_ decode.regfile.registers_27\[9\] _11258_ VGND VGND VPWR VPWR _11680_
+ sky130_fd_sc_hd__or3_1
X_27678_ clknet_leaf_21_clock _00707_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17431_ decode.regfile.registers_9\[16\] _12776_ _12592_ _12532_ _12598_ VGND VGND
+ VPWR VPWR _13380_ sky130_fd_sc_hd__a41o_1
X_29417_ clknet_leaf_257_clock _02430_ VGND VGND VPWR VPWR decode.regfile.registers_5\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14643_ execute.io_target_pc\[22\] _10677_ _10679_ _10683_ _10685_ VGND VGND VPWR
+ VPWR _10686_ sky130_fd_sc_hd__o2111a_1
X_26629_ _09383_ _09666_ VGND VGND VPWR VPWR _09672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_213_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17362_ _12530_ _10591_ _12557_ decode.regfile.registers_0\[14\] VGND VGND VPWR VPWR
+ _13313_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29348_ clknet_leaf_228_clock _02361_ VGND VGND VPWR VPWR decode.regfile.registers_3\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_57_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_57_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14574_ _10616_ VGND VGND VPWR VPWR _10617_ sky130_fd_sc_hd__clkbuf_4
X_19101_ _03670_ net261 _04320_ net317 VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16313_ _11313_ decode.regfile.registers_4\[26\] _10647_ _10629_ _11462_ VGND VGND
+ VPWR VPWR _12284_ sky130_fd_sc_hd__a2111o_1
X_13525_ _09902_ VGND VGND VPWR VPWR _09903_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_153_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29279_ clknet_leaf_241_clock _02292_ VGND VGND VPWR VPWR decode.regfile.registers_1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_17293_ decode.regfile.registers_19\[12\] _12679_ _12906_ _13245_ VGND VGND VPWR
+ VPWR _13246_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19032_ _04317_ _04319_ _04323_ _04329_ _04330_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16244_ decode.regfile.registers_10\[24\] _11183_ _12215_ _12216_ VGND VGND VPWR
+ VPWR _12217_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16175_ _11382_ decode.regfile.registers_10\[22\] _11364_ _12149_ VGND VGND VPWR
+ VPWR _12150_ sky130_fd_sc_hd__o211a_1
Xoutput107 net107 VGND VGND VPWR VPWR io_memory_address[16] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15126_ _11122_ VGND VGND VPWR VPWR _11123_ sky130_fd_sc_hd__clkbuf_4
Xoutput118 net118 VGND VGND VPWR VPWR io_memory_address[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput129 net129 VGND VGND VPWR VPWR io_memory_address[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15057_ _11053_ VGND VGND VPWR VPWR _11054_ sky130_fd_sc_hd__clkbuf_8
X_19934_ _03588_ _04238_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14008_ net768 _10258_ _10263_ _10262_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_183_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19865_ _04338_ _05006_ _05062_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18816_ _03706_ decode.id_ex_imm_reg\[12\] _04113_ _04114_ VGND VGND VPWR VPWR _04115_
+ sky130_fd_sc_hd__a22oi_4
X_19796_ _03772_ net196 _03775_ _03806_ _03809_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_208_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15959_ _11489_ decode.regfile.registers_28\[16\] decode.regfile.registers_29\[16\]
+ _11255_ VGND VGND VPWR VPWR _11940_ sky130_fd_sc_hd__o22a_1
X_18747_ net207 net206 net203 VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__o21ai_4
X_18678_ _03675_ _03685_ decode.id_ex_rs1_data_reg\[0\] _03655_ VGND VGND VPWR VPWR
+ _03977_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_37_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17629_ decode.regfile.registers_0\[21\] _12631_ _12508_ _12933_ VGND VGND VPWR VPWR
+ _03035_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_82_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20640_ csr.minstret\[28\] _05573_ _05585_ csr.mcycle\[28\] VGND VGND VPWR VPWR _05772_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20571_ csr.minstret\[18\] _05573_ _05585_ csr.mcycle\[18\] VGND VGND VPWR VPWR _05713_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22310_ _06684_ _06904_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23290_ _07619_ _07573_ _07620_ _07720_ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__a31o_1
XFILLER_0_160_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22241_ fetch.bht.bhtTable_tag\[0\]\[19\] fetch.bht.bhtTable_tag\[1\]\[19\] _06706_
+ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22172_ _06636_ _06760_ _06766_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_30_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21123_ _06050_ _06046_ net877 VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26980_ net2653 _09866_ _09873_ _09865_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25931_ _08929_ _09253_ VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__nand2_1
X_21054_ execute.csr_read_data_out_reg\[16\] _06002_ _06010_ VGND VGND VPWR VPWR _06013_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20005_ _05222_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__clkbuf_4
X_28650_ clknet_leaf_97_clock _01663_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_25862_ _08935_ _09210_ VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_226_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27601_ clknet_leaf_152_clock _00630_ VGND VGND VPWR VPWR execute.io_target_pc\[10\]
+ sky130_fd_sc_hd__dfxtp_4
X_24813_ _08593_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28581_ clknet_leaf_139_clock _01594_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25793_ _08941_ _09166_ VGND VGND VPWR VPWR _09177_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27532_ clknet_leaf_156_clock _00561_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_55_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24744_ _08556_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_190_Right_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21956_ net2042 _06574_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27463_ clknet_leaf_149_clock _00492_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _09955_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24675_ net977 execute.io_target_pc\[26\] _07285_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21887_ csr.io_mret_vector\[15\] _10807_ _06515_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29202_ clknet_leaf_240_clock _02215_ VGND VGND VPWR VPWR fetch.btb.btbTable\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26414_ _09533_ VGND VGND VPWR VPWR _09548_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_104_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23626_ _07959_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _05895_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__clkbuf_1
X_27394_ clknet_leaf_33_clock _00423_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_194_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29133_ clknet_leaf_81_clock _02146_ VGND VGND VPWR VPWR csr.mcycle\[17\] sky130_fd_sc_hd__dfxtp_1
X_26345_ net819 _09505_ _09508_ _09499_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__o211a_1
X_23557_ net2103 _07918_ _07915_ VGND VGND VPWR VPWR _07923_ sky130_fd_sc_hd__or3b_1
XFILLER_0_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20769_ _05853_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22508_ fetch.bht.bhtTable_target_pc\[12\]\[1\] fetch.bht.bhtTable_target_pc\[13\]\[1\]
+ fetch.bht.bhtTable_target_pc\[14\]\[1\] fetch.bht.bhtTable_target_pc\[15\]\[1\]
+ _07099_ _07101_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__mux4_1
X_29064_ clknet_leaf_166_clock _02077_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_26276_ net1945 _09462_ _09468_ _09458_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__o211a_1
X_14290_ _10426_ VGND VGND VPWR VPWR _10427_ sky130_fd_sc_hd__clkbuf_4
X_23488_ decode.control.io_funct7\[4\] _07876_ _07873_ VGND VGND VPWR VPWR _07883_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_150_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28015_ clknet_leaf_217_clock _01037_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25227_ _08066_ net2238 _08837_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__mux2_1
X_22439_ _06636_ _07024_ _07033_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_150_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25158_ _10573_ net2564 _08806_ VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_969 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24109_ _08227_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17980_ decode.regfile.registers_18\[30\] _10925_ _12569_ _11023_ _11008_ VGND VGND
+ VPWR VPWR _03377_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_204_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25089_ _08772_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_179_Left_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16931_ _12726_ VGND VGND VPWR VPWR _12892_ sky130_fd_sc_hd__clkbuf_4
X_28917_ clknet_leaf_116_clock _01930_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_29897_ clknet_leaf_301_clock _02910_ VGND VGND VPWR VPWR decode.regfile.registers_20\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_196_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16862_ _12536_ VGND VGND VPWR VPWR _12824_ sky130_fd_sc_hd__clkbuf_4
X_19650_ _04829_ _04831_ _04928_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__a21oi_2
X_28848_ clknet_leaf_119_clock _01861_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_205_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_1200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_221_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15813_ _11263_ decode.regfile.registers_22\[13\] _11404_ _10978_ _11265_ VGND VGND
+ VPWR VPWR _11797_ sky130_fd_sc_hd__o2111a_1
X_18601_ memory.csr_read_data_out_reg\[19\] _09986_ _10078_ _10079_ VGND VGND VPWR
+ VPWR _03900_ sky130_fd_sc_hd__o22a_2
X_19581_ _04197_ _04198_ _03929_ _03933_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__o211ai_4
X_28779_ clknet_leaf_95_clock _01792_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16793_ decode.regfile.registers_23\[1\] _12714_ _12715_ _12756_ _12514_ VGND VGND
+ VPWR VPWR _12757_ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18532_ execute.csr_read_data_out_reg\[25\] _03659_ net117 _03666_ VGND VGND VPWR
+ VPWR _03831_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15744_ decode.regfile.registers_1\[11\] _11117_ _11057_ _11109_ VGND VGND VPWR VPWR
+ _11730_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18463_ _03730_ _03731_ _03740_ _03761_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__and4_1
XFILLER_0_158_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _11194_ decode.regfile.registers_12\[9\] decode.regfile.registers_13\[9\]
+ _11196_ VGND VGND VPWR VPWR _11663_ sky130_fd_sc_hd__o22a_1
XFILLER_0_213_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17414_ _12822_ decode.regfile.registers_21\[15\] _13164_ _13363_ VGND VGND VPWR
+ VPWR _13364_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_188_Left_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14626_ _10644_ _10653_ _10664_ _10668_ VGND VGND VPWR VPWR _10669_ sky130_fd_sc_hd__or4b_1
X_18394_ _03691_ _03692_ _03683_ _03671_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__nand4_2
XFILLER_0_157_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17345_ _13183_ _13293_ _13295_ _13296_ VGND VGND VPWR VPWR _13297_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14557_ decode.id_ex_ex_rd_reg\[4\] _10595_ _10596_ _10599_ VGND VGND VPWR VPWR _10600_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13508_ _09888_ csr.io_mem_pc\[2\] VGND VGND VPWR VPWR _09889_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17276_ decode.regfile.registers_2\[12\] _12835_ _12836_ _13228_ VGND VGND VPWR VPWR
+ _13229_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14488_ _10112_ _10530_ VGND VGND VPWR VPWR _10540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19015_ net314 _04307_ _04308_ _04313_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__o31a_1
XFILLER_0_70_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16227_ _11398_ _12199_ _12200_ _11246_ VGND VGND VPWR VPWR _12201_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_228_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16158_ _11243_ VGND VGND VPWR VPWR _12133_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_185_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15109_ _11105_ VGND VGND VPWR VPWR _11106_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_75_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_197_Left_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16089_ _11192_ _11318_ _11084_ decode.regfile.registers_5\[20\] _12065_ VGND VGND
+ VPWR VPWR _12066_ sky130_fd_sc_hd__o32a_1
XFILLER_0_121_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19917_ _03862_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1091 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19848_ _04303_ _05117_ _05118_ _04360_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__o31a_1
XFILLER_0_223_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19779_ _05045_ _05031_ _04525_ _05052_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_78_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_218_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21810_ net572 _06467_ _06475_ _10546_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22790_ net1739 _10817_ _07286_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21741_ net1168 _10878_ _06428_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24460_ _08409_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__clkbuf_1
X_21672_ _05691_ csr.minstret\[16\] _06366_ _06380_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__and4_1
XFILLER_0_114_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23411_ fetch.bht.bhtTable_target_pc\[8\]\[31\] fetch.bht.bhtTable_target_pc\[9\]\[31\]
+ fetch.bht.bhtTable_target_pc\[10\]\[31\] fetch.bht.bhtTable_target_pc\[11\]\[31\]
+ _07066_ _06661_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_43_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20623_ csr.mcycle\[25\] _05552_ _05618_ csr._csr_read_data_T_8\[25\] _05757_ VGND
+ VGND VPWR VPWR _05758_ sky130_fd_sc_hd__a221o_1
XFILLER_0_163_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24391_ net1509 execute.io_target_pc\[18\] _08367_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26130_ net1752 _09330_ _09369_ _09370_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23342_ execute.io_target_pc\[26\] _07090_ _10970_ _06037_ VGND VGND VPWR VPWR _07769_
+ sky130_fd_sc_hd__a211o_1
X_20554_ csr.mscratch\[16\] _05592_ _05611_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26061_ _08982_ _09330_ VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__nand2_1
X_23273_ _09956_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__buf_2
X_20485_ csr.minstret\[7\] _05571_ _05561_ csr.mcycle\[7\] _05637_ VGND VGND VPWR
+ VPWR _05638_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25012_ net2415 _08635_ _08721_ _06419_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22224_ _06672_ _06816_ _06818_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__a21oi_1
X_22155_ fetch.bht.bhtTable_tag\[14\]\[23\] fetch.bht.bhtTable_tag\[15\]\[23\] _06618_
+ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__mux2_1
X_29820_ clknet_leaf_307_clock _02833_ VGND VGND VPWR VPWR decode.regfile.registers_18\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21106_ net2425 _06044_ _06035_ _05856_ _05858_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__o311a_1
XFILLER_0_199_1260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22086_ fetch.bht.bhtTable_tag\[4\]\[7\] fetch.bht.bhtTable_tag\[5\]\[7\] _06680_
+ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__mux2_1
X_26963_ net201 _09862_ VGND VGND VPWR VPWR _09864_ sky130_fd_sc_hd__nand2_1
X_29751_ clknet_leaf_285_clock _02764_ VGND VGND VPWR VPWR decode.regfile.registers_15\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28702_ clknet_leaf_173_clock _01715_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_25914_ _08912_ _09243_ VGND VGND VPWR VPWR _09247_ sky130_fd_sc_hd__nand2_1
X_21037_ execute.csr_read_data_out_reg\[8\] _06002_ _05998_ VGND VGND VPWR VPWR _06004_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_121_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29682_ clknet_leaf_283_clock _02695_ VGND VGND VPWR VPWR decode.regfile.registers_13\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26894_ _09701_ VGND VGND VPWR VPWR _09825_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28633_ clknet_leaf_123_clock _01646_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_25845_ _08918_ _09200_ VGND VGND VPWR VPWR _09207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28564_ clknet_leaf_209_clock _01577_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_13790_ memory.csr_read_data_out_reg\[28\] _09988_ _10126_ VGND VGND VPWR VPWR _10127_
+ sky130_fd_sc_hd__o21ai_4
X_25776_ net654 _09156_ _09167_ _09153_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__o211a_1
X_22988_ _07125_ _07434_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__and2b_1
XFILLER_0_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27515_ clknet_leaf_28_clock _00544_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dfxtp_1
X_24727_ _08089_ net1489 _08542_ VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28495_ clknet_leaf_190_clock _01508_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21939_ _06565_ _06493_ _06566_ _06567_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27446_ clknet_leaf_147_clock _00475_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15460_ _11406_ VGND VGND VPWR VPWR _11453_ sky130_fd_sc_hd__buf_2
X_24658_ net1101 VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14411_ _10107_ _10487_ VGND VGND VPWR VPWR _10496_ sky130_fd_sc_hd__nand2_1
X_23609_ _07950_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15391_ _11363_ _11384_ _11385_ _11199_ VGND VGND VPWR VPWR _11386_ sky130_fd_sc_hd__o211a_1
X_27377_ clknet_leaf_21_clock _00406_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_24589_ net1516 execute.io_target_pc\[16\] _08473_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_189_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29116_ clknet_leaf_70_clock _02129_ VGND VGND VPWR VPWR csr.mcycle\[0\] sky130_fd_sc_hd__dfxtp_2
X_17130_ _12494_ VGND VGND VPWR VPWR _13087_ sky130_fd_sc_hd__buf_2
XFILLER_0_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26328_ _09417_ VGND VGND VPWR VPWR _09499_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14342_ _10122_ _10444_ VGND VGND VPWR VPWR _10456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29047_ clknet_leaf_124_clock _02060_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_17061_ decode.regfile.registers_6\[7\] _10602_ _12626_ _12645_ VGND VGND VPWR VPWR
+ _13019_ sky130_fd_sc_hd__o31a_1
XFILLER_0_122_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26259_ _09446_ VGND VGND VPWR VPWR _09459_ sky130_fd_sc_hd__clkbuf_4
X_14273_ net666 _10377_ _10415_ _10411_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16012_ decode.regfile.registers_1\[18\] _11539_ VGND VGND VPWR VPWR _11991_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_223_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_223_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ decode.regfile.registers_19\[29\] _10599_ _10588_ _12518_ VGND VGND VPWR
+ VPWR _03361_ sky130_fd_sc_hd__or4_1
XFILLER_0_97_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19702_ _04189_ _03894_ _04977_ _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__o31a_1
X_16914_ decode.regfile.registers_14\[4\] _10924_ _12589_ _10612_ VGND VGND VPWR VPWR
+ _12875_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17894_ _10938_ decode.regfile.registers_25\[27\] _13482_ _12811_ VGND VGND VPWR
+ VPWR _03294_ sky130_fd_sc_hd__or4_1
XFILLER_0_205_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19633_ _03938_ _04912_ _03924_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_217_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16845_ decode.regfile.registers_22\[2\] _12528_ _12805_ _12807_ _12687_ VGND VGND
+ VPWR VPWR _12808_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_192_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16776_ decode.regfile.registers_8\[1\] _10593_ _12549_ _12592_ _12605_ VGND VGND
+ VPWR VPWR _12740_ sky130_fd_sc_hd__a41o_1
X_19564_ _03929_ _04180_ _04253_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__mux2_1
X_13988_ _09993_ _10244_ VGND VGND VPWR VPWR _10252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15727_ _10956_ _11217_ _11085_ decode.regfile.registers_21\[10\] _11648_ VGND VGND
+ VPWR VPWR _11714_ sky130_fd_sc_hd__o32a_1
X_18515_ _03811_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__nand2_2
X_19495_ _04085_ _04225_ _04504_ _04186_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__a211o_1
XFILLER_0_220_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15658_ _10961_ VGND VGND VPWR VPWR _11646_ sky130_fd_sc_hd__clkbuf_4
X_18446_ net208 net206 _03744_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_201_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14609_ _10651_ VGND VGND VPWR VPWR _10652_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18377_ _09934_ decode.id_ex_ex_rs1_reg\[3\] VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__nand2_1
X_15589_ _11153_ decode.regfile.registers_0\[7\] VGND VGND VPWR VPWR _11579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17328_ decode.regfile.registers_13\[13\] _12775_ _13278_ _13279_ _12663_ VGND VGND
+ VPWR VPWR _13280_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17259_ _13183_ _13210_ _13211_ _13212_ VGND VGND VPWR VPWR _13213_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_77_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20270_ _05214_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_133_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2503 decode.id_ex_rs1_data_reg\[19\] VGND VGND VPWR VPWR net2730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 _10702_ VGND VGND VPWR VPWR net2741 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2525 execute.io_reg_pc\[0\] VGND VGND VPWR VPWR net2752 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2536 csr.minstret\[9\] VGND VGND VPWR VPWR net2763 sky130_fd_sc_hd__dlygate4sd3_1
X_23960_ _08150_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__clkbuf_1
Xhold1802 fetch.bht.bhtTable_target_pc\[2\]\[1\] VGND VGND VPWR VPWR net2029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2547 csr._mcycle_T_2\[22\] VGND VGND VPWR VPWR net2774 sky130_fd_sc_hd__buf_1
XFILLER_0_227_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1813 fetch.bht.bhtTable_tag\[5\]\[22\] VGND VGND VPWR VPWR net2040 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2558 decode.regfile.registers_30\[7\] VGND VGND VPWR VPWR net2785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2569 csr._mcycle_T_2\[10\] VGND VGND VPWR VPWR net2796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1824 decode.regfile.registers_15\[22\] VGND VGND VPWR VPWR net2051 sky130_fd_sc_hd__dlygate4sd3_1
X_22911_ _06834_ _07360_ _06849_ _07361_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__or4b_1
XFILLER_0_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1835 decode.regfile.registers_8\[19\] VGND VGND VPWR VPWR net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1846 fetch.bht.bhtTable_tag\[0\]\[14\] VGND VGND VPWR VPWR net2073 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23891_ net976 _08049_ _06179_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__mux2_1
Xhold1857 decode.regfile.registers_20\[11\] VGND VGND VPWR VPWR net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1868 decode.regfile.registers_18\[28\] VGND VGND VPWR VPWR net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25630_ net682 _09082_ _09083_ _09074_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__o211a_1
Xhold1879 decode.regfile.registers_23\[23\] VGND VGND VPWR VPWR net2106 sky130_fd_sc_hd__dlygate4sd3_1
X_22842_ net2090 _10881_ _09898_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25561_ net1966 _09039_ _09043_ _09033_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22773_ _06147_ net1839 _07276_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27300_ clknet_leaf_13_clock _00329_ VGND VGND VPWR VPWR decode.regfile.registers_31\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24512_ _08072_ net1860 _08428_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28280_ clknet_leaf_59_clock _01302_ VGND VGND VPWR VPWR csr._csr_read_data_T_8\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_21724_ net933 _06420_ _06421_ _06419_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25492_ _08943_ _08992_ VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27231_ clknet_leaf_2_clock _00260_ VGND VGND VPWR VPWR decode.regfile.registers_29\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_24443_ _08070_ net2137 _08400_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__mux2_1
X_21655_ csr._mcycle_T_2\[16\] _06321_ _06366_ _05691_ csr.minstret\[16\] VGND VGND
+ VPWR VPWR _06368_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_93_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20606_ csr.minstret\[23\] _05572_ _05582_ csr.mcycle\[23\] _05742_ VGND VGND VPWR
+ VPWR _05743_ sky130_fd_sc_hd__a221o_1
X_27162_ clknet_leaf_360_clock _00191_ VGND VGND VPWR VPWR decode.regfile.registers_27\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24374_ net1224 execute.io_target_pc\[10\] _08356_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21586_ csr.io_csr_write_address\[3\] csr.io_csr_write_address\[2\] csr.io_csr_write_enable
+ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__or3b_4
XFILLER_0_7_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26113_ net2378 _09356_ _09361_ _09359_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__o211a_1
X_23325_ fetch.bht.bhtTable_target_pc\[4\]\[25\] fetch.bht.bhtTable_target_pc\[5\]\[25\]
+ _07067_ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__mux2_1
X_20537_ csr.mscratch\[13\] _05593_ _05625_ _05672_ _05683_ VGND VGND VPWR VPWR _05684_
+ sky130_fd_sc_hd__o311a_2
XFILLER_0_127_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27093_ clknet_leaf_329_clock _00122_ VGND VGND VPWR VPWR decode.regfile.registers_25\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26044_ net2419 _09313_ _09321_ _09318_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__o211a_1
X_23256_ csr._csr_read_data_T_8\[21\] _06480_ csr.io_mret_vector\[21\] _07621_ VGND
+ VGND VPWR VPWR _07688_ sky130_fd_sc_hd__o22a_1
X_20468_ csr.mcycle\[5\] _05552_ _05575_ csr.minstret\[5\] VGND VGND VPWR VPWR _05623_
+ sky130_fd_sc_hd__a22o_1
X_22207_ fetch.bht.bhtTable_tag\[12\]\[24\] fetch.bht.bhtTable_tag\[13\]\[24\] fetch.bht.bhtTable_tag\[14\]\[24\]
+ fetch.bht.bhtTable_tag\[15\]\[24\] _06645_ _06651_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__mux4_1
X_23187_ fetch.bht.bhtTable_target_pc\[8\]\[17\] fetch.bht.bhtTable_target_pc\[9\]\[17\]
+ fetch.bht.bhtTable_target_pc\[10\]\[17\] fetch.bht.bhtTable_target_pc\[11\]\[17\]
+ _07106_ _07386_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__mux4_1
X_20399_ _05534_ _05538_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__nor2_4
X_29803_ clknet_leaf_296_clock _02816_ VGND VGND VPWR VPWR decode.regfile.registers_17\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_22138_ _06649_ _06732_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__or2b_1
X_27995_ clknet_leaf_221_clock _01017_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14960_ decode.immGen._imm_T_10\[3\] _10667_ _10975_ _10662_ VGND VGND VPWR VPWR
+ _10986_ sky130_fd_sc_hd__a22o_1
X_29734_ clknet_leaf_286_clock _02747_ VGND VGND VPWR VPWR decode.regfile.registers_15\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26946_ _10035_ _09849_ VGND VGND VPWR VPWR _09855_ sky130_fd_sc_hd__nand2_1
X_22069_ fetch.bht.bhtTable_tag\[8\]\[18\] fetch.bht.bhtTable_tag\[9\]\[18\] fetch.bht.bhtTable_tag\[10\]\[18\]
+ fetch.bht.bhtTable_tag\[11\]\[18\] _06646_ _06624_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__mux4_1
XFILLER_0_215_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13911_ _09993_ _10200_ VGND VGND VPWR VPWR _10207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_215_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26877_ _09404_ _09806_ VGND VGND VPWR VPWR _09815_ sky130_fd_sc_hd__nand2_1
X_29665_ clknet_leaf_287_clock _02678_ VGND VGND VPWR VPWR decode.regfile.registers_13\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_14891_ _10927_ VGND VGND VPWR VPWR _10928_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16630_ _12594_ VGND VGND VPWR VPWR _12595_ sky130_fd_sc_hd__clkbuf_4
X_28616_ clknet_leaf_100_clock _01629_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13842_ _10025_ _10164_ VGND VGND VPWR VPWR _10166_ sky130_fd_sc_hd__nand2_1
X_25828_ net1099 _09157_ _09196_ _09194_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29596_ clknet_leaf_289_clock _02609_ VGND VGND VPWR VPWR decode.regfile.registers_11\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16561_ _10925_ _12523_ _12525_ _11009_ VGND VGND VPWR VPWR _12526_ sky130_fd_sc_hd__and4b_1
X_28547_ clknet_leaf_167_clock _01560_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13773_ _10112_ _10075_ VGND VGND VPWR VPWR _10113_ sky130_fd_sc_hd__nand2_1
X_25759_ net693 _09156_ _09158_ _09153_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18300_ decode.id_ex_rs2_data_reg\[16\] _03605_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__and2_1
X_15512_ _11043_ decode.regfile.registers_4\[5\] _11503_ _10629_ _11083_ VGND VGND
+ VPWR VPWR _11504_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_97_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19280_ _04572_ _04573_ _04244_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__o21ai_1
X_28478_ clknet_leaf_222_clock _01491_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16492_ _10646_ _11298_ _12456_ _12457_ VGND VGND VPWR VPWR _12458_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_85_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18231_ csr.mcycle\[26\] csr.mcycle\[25\] csr.mcycle\[30\] _03565_ VGND VGND VPWR
+ VPWR _03566_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_216_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27429_ clknet_leaf_39_clock _00458_ VGND VGND VPWR VPWR decode.id_ex_regwrite_reg
+ sky130_fd_sc_hd__dfxtp_1
X_15443_ _11436_ decode.regfile.registers_26\[3\] _11349_ _10980_ _11347_ VGND VGND
+ VPWR VPWR _11437_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18162_ _10912_ _03464_ _10921_ decode.control.io_funct7\[0\] VGND VGND VPWR VPWR
+ _03509_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15374_ _11295_ VGND VGND VPWR VPWR _11369_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_212_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17113_ decode.regfile.registers_13\[8\] _12512_ _12723_ _12984_ VGND VGND VPWR VPWR
+ _13070_ sky130_fd_sc_hd__o31a_1
XFILLER_0_110_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14325_ net750 _10434_ _10446_ _10440_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__o211a_1
X_18093_ _03472_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17044_ _12494_ decode.regfile.registers_26\[6\] _13002_ _11010_ _11026_ VGND VGND
+ VPWR VPWR _13003_ sky130_fd_sc_hd__o2111a_1
Xhold409 csr._mcycle_T_3\[58\] VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ net2273 _10403_ _10406_ _10398_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_225_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_146_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14187_ _10117_ _10355_ VGND VGND VPWR VPWR _10366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_221_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18995_ net309 VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17946_ decode.regfile.registers_2\[29\] _12634_ _12628_ _03343_ VGND VGND VPWR VPWR
+ _03344_ sky130_fd_sc_hd__o211ai_2
Xhold1109 fetch.bht.bhtTable_target_pc\[15\]\[29\] VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_163_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17877_ _12601_ _03276_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__nand2_1
X_19616_ _04847_ _04896_ _04277_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__mux2_1
X_16828_ _11017_ _10588_ _12637_ _10605_ VGND VGND VPWR VPWR _12791_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_176_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19547_ _04083_ _04084_ net254 _04091_ _04081_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16759_ _12722_ VGND VGND VPWR VPWR _12723_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_66_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19478_ _04762_ _04763_ _04496_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__nand3_1
XFILLER_0_186_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_340 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_351 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_362 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18429_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__buf_4
XINSDIODE1_373 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_384 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21440_ _06235_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_135_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21371_ _06119_ net1287 _06188_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23110_ _07130_ _07549_ _07550_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__nand3_1
XFILLER_0_142_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20322_ decode.id_ex_pc_reg\[24\] _05490_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24090_ _08217_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold910 decode.regfile.registers_10\[8\] VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold921 decode.regfile.registers_5\[19\] VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 _01183_ VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold943 fetch.bht.bhtTable_target_pc\[11\]\[6\] VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__dlygate4sd3_1
X_23041_ execute.io_target_pc\[8\] _05864_ _07091_ _07485_ _07347_ VGND VGND VPWR
+ VPWR _07486_ sky130_fd_sc_hd__a311o_1
X_20253_ _10730_ decode.id_ex_pc_reg\[8\] _05433_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__and3_1
Xhold954 fetch.bht.bhtTable_target_pc\[11\]\[18\] VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 fetch.bht.bhtTable_tag\[10\]\[8\] VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 _08507_ VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold987 _10680_ VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold998 fetch.bht.bhtTable_target_pc\[13\]\[13\] VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__dlygate4sd3_1
X_20184_ _00574_ _05226_ _05384_ _05239_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_34_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2300 decode.regfile.registers_19\[20\] VGND VGND VPWR VPWR net2527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26800_ _09701_ VGND VGND VPWR VPWR _09771_ sky130_fd_sc_hd__buf_2
Xhold2311 decode.regfile.registers_24\[22\] VGND VGND VPWR VPWR net2538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2322 decode.regfile.registers_24\[26\] VGND VGND VPWR VPWR net2549 sky130_fd_sc_hd__dlygate4sd3_1
X_27780_ clknet_leaf_33_clock _00809_ VGND VGND VPWR VPWR memory.io_wb_readdata\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2333 csr._minstret_T_3\[32\] VGND VGND VPWR VPWR net2560 sky130_fd_sc_hd__dlygate4sd3_1
X_24992_ net2581 _08704_ _08707_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_216_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2344 decode.regfile.registers_11\[18\] VGND VGND VPWR VPWR net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1610 decode.regfile.registers_16\[19\] VGND VGND VPWR VPWR net1837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2355 decode.regfile.registers_6\[25\] VGND VGND VPWR VPWR net2582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 fetch.bht.bhtTable_target_pc\[14\]\[2\] VGND VGND VPWR VPWR net1848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26731_ _09408_ _09720_ VGND VGND VPWR VPWR _09731_ sky130_fd_sc_hd__nand2_1
Xhold2366 decode.regfile.registers_26\[29\] VGND VGND VPWR VPWR net2593 sky130_fd_sc_hd__dlygate4sd3_1
X_23943_ net1124 _08101_ _06156_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1632 decode.regfile.registers_13\[30\] VGND VGND VPWR VPWR net1859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2377 csr._csr_read_data_T_8\[19\] VGND VGND VPWR VPWR net2604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2388 decode.regfile.registers_12\[16\] VGND VGND VPWR VPWR net2615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1643 decode.regfile.registers_6\[2\] VGND VGND VPWR VPWR net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1654 fetch.bht.bhtTable_tag\[8\]\[24\] VGND VGND VPWR VPWR net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2399 csr.mtie VGND VGND VPWR VPWR net2626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1665 fetch.bht.bhtTable_target_pc\[15\]\[19\] VGND VGND VPWR VPWR net1892 sky130_fd_sc_hd__dlygate4sd3_1
X_29450_ clknet_leaf_262_clock _02463_ VGND VGND VPWR VPWR decode.regfile.registers_6\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1676 fetch.bht.bhtTable_target_pc\[13\]\[10\] VGND VGND VPWR VPWR net1903 sky130_fd_sc_hd__dlygate4sd3_1
X_26662_ _09415_ _09689_ VGND VGND VPWR VPWR _09691_ sky130_fd_sc_hd__nand2_1
X_23874_ _08103_ net1428 _07940_ VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__mux2_1
Xhold1687 _01222_ VGND VGND VPWR VPWR net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1698 decode.regfile.registers_10\[15\] VGND VGND VPWR VPWR net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28401_ clknet_leaf_142_clock _01414_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfxtp_4
X_25613_ _08990_ VGND VGND VPWR VPWR _09074_ sky130_fd_sc_hd__clkbuf_4
X_22825_ _07284_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__clkbuf_8
X_29381_ clknet_leaf_258_clock _02394_ VGND VGND VPWR VPWR decode.regfile.registers_4\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26593_ net1877 _09649_ _09651_ _09648_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__o211a_1
X_28332_ clknet_leaf_216_clock _01345_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25544_ _08918_ _09026_ VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__nand2_1
X_22756_ _06130_ net1659 _07265_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21707_ _05691_ csr.minstret\[16\] csr.minstret\[17\] csr.minstret\[18\] VGND VGND
+ VPWR VPWR _06408_ sky130_fd_sc_hd__and4_1
X_28263_ clknet_leaf_77_clock _01285_ VGND VGND VPWR VPWR csr._minstret_T_3\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25475_ _08925_ _08992_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22687_ csr._mcycle_T_2\[19\] _07223_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27214_ clknet_leaf_3_clock _00243_ VGND VGND VPWR VPWR decode.regfile.registers_28\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_229_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24426_ _08053_ net1496 _08389_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28194_ clknet_leaf_112_clock _01216_ VGND VGND VPWR VPWR csr.io_mret_vector\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_21638_ csr.minstret\[11\] _06349_ _06354_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_229_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27145_ clknet_leaf_358_clock _00174_ VGND VGND VPWR VPWR decode.regfile.registers_26\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24357_ net1179 execute.io_target_pc\[2\] _06141_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21569_ _06140_ net2315 _06295_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14110_ _10112_ _10312_ VGND VGND VPWR VPWR _10322_ sky130_fd_sc_hd__nand2_1
X_23308_ fetch.bht.bhtTable_target_pc\[8\]\[24\] fetch.bht.bhtTable_target_pc\[9\]\[24\]
+ fetch.bht.bhtTable_target_pc\[10\]\[24\] fetch.bht.bhtTable_target_pc\[11\]\[24\]
+ _07708_ _07710_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27076_ clknet_leaf_346_clock _00105_ VGND VGND VPWR VPWR decode.regfile.registers_24\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_15090_ _11086_ VGND VGND VPWR VPWR _11087_ sky130_fd_sc_hd__clkbuf_4
X_24288_ _08319_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14041_ net2520 _10271_ _10281_ _10275_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__o211a_1
X_26027_ _08948_ _09310_ VGND VGND VPWR VPWR _09312_ sky130_fd_sc_hd__nand2_1
X_23239_ _07653_ _07654_ _07672_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17800_ decode.regfile.registers_11\[25\] _12595_ _12772_ _12541_ VGND VGND VPWR
+ VPWR _03202_ sky130_fd_sc_hd__o2bb2a_1
X_15992_ _11948_ _11971_ _11454_ VGND VGND VPWR VPWR _11972_ sky130_fd_sc_hd__o21ai_1
X_18780_ net105 _03665_ _04078_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_219_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27978_ clknet_leaf_197_clock _01000_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14943_ _10971_ _10757_ _10672_ _10908_ VGND VGND VPWR VPWR _10972_ sky130_fd_sc_hd__or4_4
X_17731_ decode.regfile.registers_21\[23\] _12716_ _03111_ _03134_ _13164_ VGND VGND
+ VPWR VPWR _03135_ sky130_fd_sc_hd__o221a_1
X_29717_ clknet_leaf_284_clock _02730_ VGND VGND VPWR VPWR decode.regfile.registers_14\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26929_ net552 _09840_ VGND VGND VPWR VPWR _09845_ sky130_fd_sc_hd__nand2_1
X_14874_ _10915_ VGND VGND VPWR VPWR _10916_ sky130_fd_sc_hd__buf_2
X_29648_ clknet_leaf_280_clock _02661_ VGND VGND VPWR VPWR decode.regfile.registers_12\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_17662_ _12667_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19401_ _04166_ _04137_ _04234_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_218_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16613_ _12577_ VGND VGND VPWR VPWR _12578_ sky130_fd_sc_hd__buf_2
X_13825_ net1306 _10153_ _10156_ _10132_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17593_ decode.regfile.registers_13\[20\] _12927_ _12583_ _12663_ VGND VGND VPWR
+ VPWR _03000_ sky130_fd_sc_hd__a31o_1
X_29579_ clknet_leaf_266_clock _02592_ VGND VGND VPWR VPWR decode.regfile.registers_10\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16544_ _10601_ _12508_ VGND VGND VPWR VPWR _12509_ sky130_fd_sc_hd__nand2_4
X_19332_ _04234_ _04062_ _04487_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__o21ai_1
X_13756_ net2503 _10083_ _10098_ _10077_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19263_ _03638_ _04045_ _04504_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__a21oi_1
X_16475_ decode.regfile.registers_23\[30\] _11087_ _12417_ _12441_ VGND VGND VPWR
+ VPWR _12442_ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13687_ _09977_ _09978_ memory.io_wb_reg_pc\[12\] VGND VGND VPWR VPWR _10040_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18214_ _10910_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15426_ decode.regfile.registers_11\[3\] _11181_ _11184_ decode.regfile.registers_10\[3\]
+ VGND VGND VPWR VPWR _11420_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_143_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19194_ _04330_ _04480_ _04485_ _04409_ _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18145_ _03495_ _03493_ _03500_ net2122 VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__and4bb_1
Xclkbuf_leaf_340_clock clknet_5_5__leaf_clock VGND VGND VPWR VPWR clknet_leaf_340_clock
+ sky130_fd_sc_hd__clkbuf_8
X_15357_ _10990_ _11072_ _11065_ _10957_ VGND VGND VPWR VPWR _11352_ sky130_fd_sc_hd__and4_1
XFILLER_0_182_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire170 net171 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14308_ _10042_ _10431_ VGND VGND VPWR VPWR _10437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18076_ _03461_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__buf_1
XFILLER_0_123_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire181 _00656_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
Xhold206 decode.control.io_funct7\[4\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ _11283_ VGND VGND VPWR VPWR _11284_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_169_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire192 _10111_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_4
XFILLER_0_79_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold217 io_fetch_data[9] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 decode.io_wfi_out VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17027_ decode.regfile.registers_15\[6\] _12585_ _12983_ _12985_ VGND VGND VPWR VPWR
+ _12986_ sky130_fd_sc_hd__a22oi_1
X_14239_ net1939 _10390_ _10396_ _10385_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__o211a_1
Xhold239 decode.id_ex_memtoreg_reg\[0\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_355_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_355_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_91_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18978_ _04264_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__buf_4
XFILLER_0_225_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ decode.regfile.registers_23\[28\] _12714_ _03303_ _03327_ _12515_ VGND VGND
+ VPWR VPWR _03328_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_68_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20940_ _05951_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_124_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_1122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20871_ _05913_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22610_ csr._minstret_T_3\[51\] csr._minstret_T_3\[50\] csr._minstret_T_3\[49\] _07178_
+ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__and4_1
XFILLER_0_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23590_ _07929_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_220_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22541_ net78 _07065_ _07132_ _07134_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_27_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_170 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_181 execute.io_reg_pc\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_192 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25260_ _08099_ net1643 _09906_ VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22472_ _07066_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24211_ _08105_ net1281 _06251_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21423_ _06226_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25191_ net425 _08824_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_783 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24142_ _08244_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21354_ _06189_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20305_ _05340_ _10867_ _05473_ decode.id_ex_rdsel_reg VGND VGND VPWR VPWR _05480_
+ sky130_fd_sc_hd__a31o_1
X_28950_ clknet_leaf_124_clock _01963_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_24073_ net1283 execute.io_target_pc\[24\] _07991_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold740 fetch.bht.bhtTable_target_pc\[4\]\[18\] VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__dlygate4sd3_1
X_21285_ net994 _06149_ _06141_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__mux2_1
Xhold751 fetch.bht.bhtTable_target_pc\[2\]\[13\] VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold762 fetch.bht.bhtTable_target_pc\[2\]\[25\] VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23024_ _06248_ _07467_ _07469_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__o21ai_1
X_27901_ clknet_leaf_82_clock _00930_ VGND VGND VPWR VPWR csr._mcycle_T_2\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold773 decode.regfile.registers_29\[21\] VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20236_ _10834_ _10747_ decode.id_ex_pc_reg\[4\] VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__and3_1
X_28881_ clknet_leaf_103_clock _01894_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold784 fetch.bht.bhtTable_target_pc\[4\]\[11\] VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold795 fetch.bht.bhtTable_target_pc\[2\]\[17\] VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20167_ _05368_ _05369_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__and2b_1
X_27832_ clknet_leaf_321_clock _00861_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2130 decode.regfile.registers_10\[16\] VGND VGND VPWR VPWR net2357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2141 decode.regfile.registers_25\[31\] VGND VGND VPWR VPWR net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2152 decode.regfile.registers_3\[24\] VGND VGND VPWR VPWR net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2163 csr.mscratch\[21\] VGND VGND VPWR VPWR net2390 sky130_fd_sc_hd__dlygate4sd3_1
X_20098_ decode.id_ex_imm_reg\[13\] decode.id_ex_pc_reg\[13\] VGND VGND VPWR VPWR
+ _05311_ sky130_fd_sc_hd__nand2_1
X_24975_ _07199_ _08695_ _08696_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__nor3_1
X_27763_ clknet_leaf_315_clock _00792_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2174 decode.regfile.registers_25\[1\] VGND VGND VPWR VPWR net2401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1440 fetch.bht.bhtTable_target_pc\[10\]\[15\] VGND VGND VPWR VPWR net1667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2185 decode.regfile.registers_15\[17\] VGND VGND VPWR VPWR net2412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 decode.regfile.registers_16\[11\] VGND VGND VPWR VPWR net1678 sky130_fd_sc_hd__dlygate4sd3_1
X_29502_ clknet_leaf_251_clock _02515_ VGND VGND VPWR VPWR decode.regfile.registers_8\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_23926_ _08133_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__clkbuf_1
Xhold2196 csr._csr_read_data_T_8\[15\] VGND VGND VPWR VPWR net2423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26714_ net1041 _09709_ _09721_ _09717_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1462 fetch.bht.bhtTable_tag\[2\]\[11\] VGND VGND VPWR VPWR net1689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27694_ clknet_leaf_24_clock _00723_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1473 fetch.bht.bhtTable_tag\[15\]\[23\] VGND VGND VPWR VPWR net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 fetch.bht.bhtTable_target_pc\[3\]\[6\] VGND VGND VPWR VPWR net1711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_200_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 fetch.bht.bhtTable_tag\[13\]\[6\] VGND VGND VPWR VPWR net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1099 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26645_ net529 _09679_ _09681_ _09675_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__o211a_1
X_29433_ clknet_leaf_248_clock _02446_ VGND VGND VPWR VPWR decode.regfile.registers_5\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_23857_ _08092_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13610_ _09939_ _09940_ memory.io_wb_readdata\[3\] VGND VGND VPWR VPWR _09972_ sky130_fd_sc_hd__and3b_1
XFILLER_0_196_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22808_ _07299_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29364_ clknet_leaf_227_clock _02377_ VGND VGND VPWR VPWR decode.regfile.registers_3\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_26576_ net2133 _09636_ _09641_ _09635_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__o211a_1
X_14590_ _10632_ VGND VGND VPWR VPWR _10633_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23788_ _08046_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28315_ clknet_leaf_202_clock _01328_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13541_ _09915_ VGND VGND VPWR VPWR _09916_ sky130_fd_sc_hd__clkbuf_4
X_25527_ _09022_ VGND VGND VPWR VPWR _09023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22739_ _06113_ net1846 _09903_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__mux2_1
X_29295_ clknet_leaf_225_clock _02308_ VGND VGND VPWR VPWR decode.regfile.registers_1\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28246_ clknet_leaf_77_clock _01268_ VGND VGND VPWR VPWR csr._minstret_T_3\[46\]
+ sky130_fd_sc_hd__dfxtp_2
X_16260_ _11679_ decode.regfile.registers_27\[24\] _11869_ VGND VGND VPWR VPWR _12233_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25458_ _08910_ _08980_ VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15211_ _11207_ VGND VGND VPWR VPWR _11208_ sky130_fd_sc_hd__clkbuf_4
X_24409_ net973 execute.io_target_pc\[27\] _09911_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28177_ clknet_leaf_60_clock _01199_ VGND VGND VPWR VPWR csr.io_mret_vector\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16191_ _11250_ _11258_ decode.regfile.registers_27\[22\] _12135_ _12165_ VGND VGND
+ VPWR VPWR _12166_ sky130_fd_sc_hd__o32a_1
XFILLER_0_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25389_ _08935_ _08923_ VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27128_ clknet_leaf_354_clock _00157_ VGND VGND VPWR VPWR decode.regfile.registers_26\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_15142_ _11138_ VGND VGND VPWR VPWR _11139_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19950_ _05209_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__clkbuf_1
X_27059_ clknet_leaf_330_clock _00088_ VGND VGND VPWR VPWR decode.regfile.registers_24\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_15073_ net321 VGND VGND VPWR VPWR _11070_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14024_ net1549 _10271_ _10272_ _10262_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__o211a_1
X_18901_ _03919_ _03920_ _03921_ _03922_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_207_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19881_ _05149_ _04401_ _05150_ _04504_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__o31a_1
XFILLER_0_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18832_ _04126_ _04129_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__and2_2
XFILLER_0_208_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18763_ _03656_ _04059_ _03670_ _04061_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__o211a_4
XFILLER_0_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ _11153_ decode.regfile.registers_0\[17\] VGND VGND VPWR VPWR _11955_ sky130_fd_sc_hd__nand2_1
X_17714_ decode.regfile.registers_3\[23\] _10616_ _12729_ _12838_ VGND VGND VPWR VPWR
+ _03118_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14926_ _10642_ VGND VGND VPWR VPWR _10955_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18694_ execute.io_mem_memtoreg\[1\] execute.io_mem_memtoreg\[0\] net111 VGND VGND
+ VPWR VPWR _03993_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_72_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17645_ decode.regfile.registers_13\[21\] _12927_ _12587_ _12662_ VGND VGND VPWR
+ VPWR _03051_ sky130_fd_sc_hd__a31o_1
XFILLER_0_199_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14857_ decode.id_ex_pc_reg\[16\] _10875_ _10877_ decode.id_ex_pc_reg\[14\] _10899_
+ VGND VGND VPWR VPWR _10900_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_63_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13808_ _10142_ _09937_ VGND VGND VPWR VPWR _10143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14788_ decode.id_ex_pc_reg\[0\] csr.io_mem_pc\[0\] VGND VGND VPWR VPWR _10831_ sky130_fd_sc_hd__nor2_1
X_17576_ _13339_ _02981_ _02982_ _02983_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19315_ _04280_ _04019_ _04484_ _04606_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__o31a_1
XFILLER_0_58_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16527_ _10939_ _12491_ _11011_ _10928_ VGND VGND VPWR VPWR _12492_ sky130_fd_sc_hd__or4b_4
X_13739_ _09943_ memory.io_wb_aluresult\[20\] _09981_ memory.io_wb_readdata\[20\]
+ _09977_ VGND VGND VPWR VPWR _10084_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_220_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19246_ _04272_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16458_ decode.regfile.registers_2\[30\] _11190_ _11148_ _11151_ _12424_ VGND VGND
+ VPWR VPWR _12425_ sky130_fd_sc_hd__o311a_1
XFILLER_0_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15409_ _11238_ VGND VGND VPWR VPWR _11403_ sky130_fd_sc_hd__clkbuf_4
X_16389_ decode.regfile.registers_6\[28\] _10637_ _11136_ _12350_ _12357_ VGND VGND
+ VPWR VPWR _12358_ sky130_fd_sc_hd__o32a_1
X_19177_ _04350_ _04354_ _04264_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18128_ _03482_ _03480_ _03487_ decode.io_id_pc\[20\] VGND VGND VPWR VPWR _03492_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_81_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_294_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_294_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18059_ decode.control.io_opcode\[3\] _10583_ _10584_ _10998_ VGND VGND VPWR VPWR
+ _03451_ sky130_fd_sc_hd__and4b_1
XFILLER_0_44_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21070_ _06021_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__buf_1
XFILLER_0_223_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20021_ _05242_ _05244_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__xor2_1
XFILLER_0_158_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24760_ _08053_ net1848 _08563_ VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__mux2_1
X_21972_ net1590 _06588_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__or2_1
Xrebuffer10 _03744_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_1
XFILLER_0_197_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer21 _03686_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_1
X_23711_ _08006_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer32 _03763_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_232_clock clknet_5_29__leaf_clock VGND VGND VPWR VPWR clknet_leaf_232_clock
+ sky130_fd_sc_hd__clkbuf_8
X_20923_ _05937_ _05933_ net47 VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__and3_1
X_24691_ _08053_ net2124 _06306_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__mux2_1
Xrebuffer43 net269 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
Xrebuffer54 _07087_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__buf_1
Xclkbuf_5_18__f_clock clknet_2_2_0_clock VGND VGND VPWR VPWR clknet_5_18__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer65 _03739_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_178_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer76 csr.io_csr_address\[3\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd1_1
X_26430_ _09410_ _09545_ VGND VGND VPWR VPWR _09557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23642_ net1694 _10871_ _07961_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20854_ _05904_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer87 _04120_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_49_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer98 _03752_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26361_ net1771 _09505_ _09517_ _09512_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__o211a_1
X_23573_ _07931_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20785_ _05856_ net417 _05858_ _05863_ _01176_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28100_ clknet_leaf_75_clock _01122_ VGND VGND VPWR VPWR csr.minstret\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_147_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25312_ _08886_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29080_ clknet_leaf_186_clock _02093_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_22524_ _07109_ _07112_ _07076_ _07117_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_247_clock clknet_5_19__leaf_clock VGND VGND VPWR VPWR clknet_leaf_247_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26292_ _09424_ _09472_ VGND VGND VPWR VPWR _09478_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28031_ clknet_leaf_202_clock _01053_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer100 _09921_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_106_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25243_ _08851_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__clkbuf_1
X_22455_ _06618_ fetch.btb.btbTable\[13\]\[1\] fetch.bht.bhtTable_valid\[13\] _06687_
+ _07049_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__a311o_1
XFILLER_0_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer111 net336 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21406_ _06216_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25174_ _08813_ _09880_ _09884_ VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__or3b_2
XFILLER_0_44_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22386_ _06623_ _06978_ _06687_ _06980_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__a211oi_1
X_24125_ net1436 execute.io_target_pc\[17\] _08232_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21337_ _06155_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24056_ _08200_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__clkbuf_1
X_28933_ clknet_leaf_141_clock _01946_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_21268_ _10772_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__buf_2
Xhold570 decode.regfile.registers_29\[10\] VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 fetch.bht.bhtTable_tag\[1\]\[20\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold592 decode.regfile.registers_13\[12\] VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__dlygate4sd3_1
X_23007_ net227 _07343_ _07344_ _07453_ _06566_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__o311a_1
X_20219_ _04459_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__buf_4
XFILLER_0_198_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28864_ clknet_leaf_161_clock _01877_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_21199_ _06086_ _05868_ net2271 VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27815_ clknet_leaf_324_clock _00844_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_202_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28795_ clknet_leaf_173_clock _01808_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15760_ decode.regfile.registers_17\[11\] _11357_ _11745_ _11268_ VGND VGND VPWR
+ VPWR _11746_ sky130_fd_sc_hd__a211o_1
XFILLER_0_188_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24958_ _07199_ _08684_ _08685_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__nor3_1
X_27746_ clknet_leaf_35_clock _00775_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1270 fetch.bht.bhtTable_target_pc\[0\]\[13\] VGND VGND VPWR VPWR net1497 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _10733_ execute.io_target_pc\[31\] _10741_ _10742_ _10753_ VGND VGND VPWR
+ VPWR _10754_ sky130_fd_sc_hd__o2111ai_2
Xhold1281 decode.regfile.registers_28\[23\] VGND VGND VPWR VPWR net1508 sky130_fd_sc_hd__dlygate4sd3_1
X_23909_ _08124_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__clkbuf_1
Xhold1292 fetch.bht.bhtTable_target_pc\[4\]\[4\] VGND VGND VPWR VPWR net1519 sky130_fd_sc_hd__dlygate4sd3_1
X_15691_ _11050_ VGND VGND VPWR VPWR _11679_ sky130_fd_sc_hd__buf_2
X_24889_ csr._mcycle_T_3\[32\] _08636_ net620 VGND VGND VPWR VPWR _08638_ sky130_fd_sc_hd__a21oi_1
X_27677_ clknet_leaf_27_clock _00706_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14642_ _10684_ execute.io_target_pc\[30\] _10680_ execute.io_target_pc\[8\] VGND
+ VGND VPWR VPWR _10685_ sky130_fd_sc_hd__o2bb2a_1
X_17430_ _11021_ _12559_ _12534_ _12673_ decode.regfile.registers_16\[16\] VGND VGND
+ VPWR VPWR _13379_ sky130_fd_sc_hd__a32o_1
X_29416_ clknet_leaf_262_clock _02429_ VGND VGND VPWR VPWR decode.regfile.registers_5\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26628_ net1960 _09665_ _09671_ _09660_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29347_ clknet_leaf_230_clock _02360_ VGND VGND VPWR VPWR decode.regfile.registers_3\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_17361_ decode.regfile.registers_2\[14\] _10608_ _12635_ net209 VGND VGND VPWR VPWR
+ _13312_ sky130_fd_sc_hd__a31o_1
X_14573_ _10615_ VGND VGND VPWR VPWR _10616_ sky130_fd_sc_hd__buf_4
XFILLER_0_200_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26559_ net2165 _09622_ _09631_ _09619_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19100_ _04396_ _04310_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13524_ _09901_ VGND VGND VPWR VPWR _09902_ sky130_fd_sc_hd__clkbuf_8
X_16312_ _12281_ _12282_ VGND VGND VPWR VPWR _12283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17292_ _13242_ _13243_ _13244_ VGND VGND VPWR VPWR _13245_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_153_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29278_ clknet_leaf_243_clock _02291_ VGND VGND VPWR VPWR decode.regfile.registers_1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19031_ _03972_ _03974_ _04007_ _04268_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__o211a_2
XFILLER_0_36_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16243_ decode.regfile.registers_8\[24\] _11284_ _11287_ decode.regfile.registers_9\[24\]
+ _11381_ VGND VGND VPWR VPWR _12216_ sky130_fd_sc_hd__o221a_1
X_28229_ clknet_leaf_62_clock _01251_ VGND VGND VPWR VPWR csr.mscratch\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16174_ _12146_ _12147_ _12148_ VGND VGND VPWR VPWR _12149_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_209_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15125_ _11058_ _10631_ _10638_ _11121_ VGND VGND VPWR VPWR _11122_ sky130_fd_sc_hd__or4_4
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput108 net108 VGND VGND VPWR VPWR io_memory_address[17] sky130_fd_sc_hd__clkbuf_4
Xoutput119 net119 VGND VGND VPWR VPWR io_memory_address[27] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_112_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15056_ _11052_ VGND VGND VPWR VPWR _11053_ sky130_fd_sc_hd__clkbuf_4
X_19933_ _05200_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__inv_2
XFILLER_0_220_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14007_ _10048_ _10255_ VGND VGND VPWR VPWR _10263_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_183_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19864_ _04295_ _04775_ _04779_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_183_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput90 net90 VGND VGND VPWR VPWR io_fetch_address[30] sky130_fd_sc_hd__clkbuf_4
X_18815_ _03751_ _03752_ net251 net237 _04108_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__a311o_1
XFILLER_0_218_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19795_ _05068_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18746_ _04044_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_121_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15958_ _11250_ _11259_ decode.regfile.registers_27\[16\] _11911_ _11938_ VGND VGND
+ VPWR VPWR _11939_ sky130_fd_sc_hd__o32a_1
XFILLER_0_204_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14909_ decode.control.io_funct3\[0\] VGND VGND VPWR VPWR _10941_ sky130_fd_sc_hd__buf_2
X_18677_ _03971_ _03975_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__nor2_2
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15889_ _11756_ decode.regfile.registers_28\[14\] _11871_ _11681_ _11440_ VGND VGND
+ VPWR VPWR _11872_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_76_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17628_ decode.regfile.registers_9\[21\] _10594_ _12690_ _12533_ _12599_ VGND VGND
+ VPWR VPWR _03034_ sky130_fd_sc_hd__a41o_1
XFILLER_0_37_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17559_ decode.regfile.registers_8\[19\] _12892_ _12602_ _02966_ VGND VGND VPWR VPWR
+ _02967_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20570_ csr._minstret_T_3\[50\] _05577_ _05578_ _05711_ VGND VGND VPWR VPWR _05712_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19229_ _04520_ _04452_ _04521_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__o31a_1
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22240_ fetch.bht.bhtTable_tag\[2\]\[19\] fetch.bht.bhtTable_tag\[3\]\[19\] _06707_
+ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22171_ _06762_ _06764_ _06765_ _06673_ _06699_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21122_ _06053_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21053_ _06012_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__clkbuf_1
X_25930_ _09241_ VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__buf_2
XFILLER_0_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20004_ _05224_ _05229_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__xnor2_1
X_25861_ net1714 _09213_ _09216_ _09209_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__o211a_1
X_24812_ _08105_ net1486 _08585_ VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__mux2_1
X_27600_ clknet_leaf_152_clock _00629_ VGND VGND VPWR VPWR execute.io_target_pc\[9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_119_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28580_ clknet_leaf_127_clock _01593_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_171_clock clknet_5_24__leaf_clock VGND VGND VPWR VPWR clknet_leaf_171_clock
+ sky130_fd_sc_hd__clkbuf_8
X_25792_ net1221 _09170_ _09176_ _09169_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24743_ _08105_ net1136 _06283_ VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__mux2_1
X_27531_ clknet_leaf_155_clock _00560_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_69_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21955_ csr._mcycle_T_2\[2\] _06572_ _06577_ _06579_ VGND VGND VPWR VPWR _01222_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27462_ clknet_leaf_138_clock _00491_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[28\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20906_ _05932_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__clkbuf_1
X_24674_ _08520_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21886_ _06529_ _06519_ _06520_ _06530_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29201_ clknet_leaf_240_clock _02214_ VGND VGND VPWR VPWR fetch.btb.btbTable\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_104_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23625_ _09885_ _09887_ _09917_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__and3_4
X_26413_ net533 _09534_ _09547_ _09540_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_186_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_186_clock
+ sky130_fd_sc_hd__clkbuf_8
X_27393_ clknet_leaf_31_clock _00422_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20837_ net105 _05891_ _05887_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_13_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29132_ clknet_leaf_82_clock _02145_ VGND VGND VPWR VPWR csr.mcycle\[16\] sky130_fd_sc_hd__dfxtp_1
X_26344_ _09400_ _09502_ VGND VGND VPWR VPWR _09508_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23556_ net220 _07917_ _07922_ _05805_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20768_ _03452_ _05425_ csr.io_csr_address\[11\] VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__and3b_1
XFILLER_0_147_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22507_ _07100_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__buf_4
X_29063_ clknet_leaf_238_clock _02076_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26275_ _09406_ _09459_ VGND VGND VPWR VPWR _09468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23487_ net21 _07875_ _07882_ _07879_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20699_ _05809_ decode.id_ex_rs1_data_reg\[10\] _05798_ VGND VGND VPWR VPWR _05817_
+ sky130_fd_sc_hd__a21oi_1
X_25226_ _08842_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__clkbuf_1
X_28014_ clknet_leaf_193_clock _01036_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22438_ _06687_ _07026_ _07028_ _06641_ _07032_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__o311a_1
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25157_ net421 _08806_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22369_ net97 _06963_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24108_ net1173 execute.io_target_pc\[9\] _08221_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_124_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_202_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25088_ _06105_ net1900 _08596_ VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28916_ clknet_leaf_118_clock _01929_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_24039_ _08191_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__clkbuf_1
X_16930_ _12612_ _12887_ _12890_ VGND VGND VPWR VPWR _12891_ sky130_fd_sc_hd__o21ai_1
X_29896_ clknet_leaf_301_clock _02909_ VGND VGND VPWR VPWR decode.regfile.registers_20\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28847_ clknet_leaf_107_clock _01860_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_196_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16861_ _12523_ VGND VGND VPWR VPWR _12823_ sky130_fd_sc_hd__buf_2
XFILLER_0_205_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18600_ _03707_ decode.id_ex_imm_reg\[19\] VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_221_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_139_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_139_clock
+ sky130_fd_sc_hd__clkbuf_8
X_15812_ _11571_ net430 _11722_ _11723_ _11724_ VGND VGND VPWR VPWR _11796_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_137_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19580_ _04861_ _04860_ _04840_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__or3b_4
X_28778_ clknet_leaf_97_clock _01791_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16792_ decode.regfile.registers_21\[1\] _12716_ _12717_ _12754_ _12755_ VGND VGND
+ VPWR VPWR _12756_ sky130_fd_sc_hd__o221a_1
XFILLER_0_204_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18531_ _03814_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__nor2_1
X_15743_ decode.regfile.registers_2\[11\] _11296_ _11141_ _11109_ VGND VGND VPWR VPWR
+ _11729_ sky130_fd_sc_hd__a2bb2o_1
X_27729_ clknet_leaf_67_clock _00758_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18462_ _03719_ decode.io_wb_rd\[3\] VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15674_ _11650_ _11661_ VGND VGND VPWR VPWR _11662_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_155_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17413_ decode.regfile.registers_20\[15\] _12770_ _13361_ _13362_ _12537_ VGND VGND
+ VPWR VPWR _13363_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14625_ decode.control.io_opcode\[5\] decode.control.io_opcode\[4\] _10665_ _10667_
+ VGND VGND VPWR VPWR _10668_ sky130_fd_sc_hd__a31o_2
XFILLER_0_28_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18393_ decode.id_ex_ex_rs1_reg\[1\] decode.io_wb_rd\[1\] VGND VGND VPWR VPWR _03692_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_200_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17344_ _13087_ decode.regfile.registers_26\[13\] _13254_ _13047_ _13088_ VGND VGND
+ VPWR VPWR _13296_ sky130_fd_sc_hd__o2111a_1
X_14556_ _10598_ VGND VGND VPWR VPWR _10599_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13507_ csr.io_mem_pc\[3\] VGND VGND VPWR VPWR _09888_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17275_ decode.regfile.registers_1\[12\] _12631_ _12633_ _13227_ VGND VGND VPWR VPWR
+ _13228_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14487_ net478 _10533_ _10539_ _10535_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19014_ net314 _04307_ _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_114_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16226_ _11489_ decode.regfile.registers_28\[23\] decode.regfile.registers_29\[23\]
+ _11255_ VGND VGND VPWR VPWR _12200_ sky130_fd_sc_hd__o22a_1
XFILLER_0_141_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer1 _03655_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__buf_4
XFILLER_0_12_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16157_ _11761_ net600 _12098_ _12131_ _12132_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_185_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_185_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15108_ _10660_ _10655_ _10640_ _11104_ VGND VGND VPWR VPWR _11105_ sky130_fd_sc_hd__or4_2
XFILLER_0_139_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16088_ _11503_ _10629_ _11043_ _11083_ VGND VGND VPWR VPWR _12065_ sky130_fd_sc_hd__or4_1
XFILLER_0_139_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_181_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15039_ _11035_ VGND VGND VPWR VPWR _11036_ sky130_fd_sc_hd__buf_4
X_19916_ _03854_ _05169_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19847_ _04436_ _05036_ _04409_ _04947_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19778_ _05016_ _05018_ _05051_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_108_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18729_ _03972_ _03974_ _04007_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_78_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21740_ _06432_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21671_ csr.minstret\[17\] csr.minstret\[18\] csr.minstret\[19\] csr.minstret\[20\]
+ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__and4_1
XFILLER_0_114_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23410_ fetch.bht.bhtTable_target_pc\[12\]\[31\] fetch.bht.bhtTable_target_pc\[13\]\[31\]
+ fetch.bht.bhtTable_target_pc\[14\]\[31\] fetch.bht.bhtTable_target_pc\[15\]\[31\]
+ _07066_ _07070_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__mux4_1
X_20622_ csr.minstret\[25\] _05594_ _05595_ csr._minstret_T_3\[57\] VGND VGND VPWR
+ VPWR _05757_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24390_ net1478 VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_43_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23341_ _07764_ _07767_ _07084_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_138_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20553_ _05697_ _03587_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26060_ net2433 _09329_ _09331_ _09318_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23272_ _06248_ _10915_ _07688_ _07703_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_131_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20484_ csr.mtie _05517_ _05527_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25011_ net1733 _08710_ _08635_ csr.mcycle\[8\] VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__a211oi_1
X_22223_ _06817_ _06686_ _00003_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_41_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_41_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22154_ _06652_ _06748_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21105_ net132 _06043_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__nor2_1
X_29750_ clknet_leaf_294_clock _02763_ VGND VGND VPWR VPWR decode.regfile.registers_15\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_22085_ net299 VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__clkbuf_8
X_26962_ net1260 _09853_ _09863_ _09852_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_56_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28701_ clknet_leaf_177_clock _01714_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21036_ _06003_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__clkbuf_1
X_25913_ net2206 _09242_ _09246_ _09235_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__o211a_1
X_29681_ clknet_leaf_283_clock _02694_ VGND VGND VPWR VPWR decode.regfile.registers_13\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26893_ _09422_ _09819_ VGND VGND VPWR VPWR _09824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28632_ clknet_leaf_122_clock _01645_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25844_ net2362 _09199_ _09206_ _09194_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28563_ clknet_leaf_203_clock _01576_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_22987_ fetch.bht.bhtTable_target_pc\[4\]\[6\] fetch.bht.bhtTable_target_pc\[5\]\[6\]
+ _07123_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__mux2_1
X_25775_ _08922_ _09166_ VGND VGND VPWR VPWR _09167_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27514_ clknet_leaf_29_clock _00543_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24726_ _08547_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__clkbuf_1
X_21938_ csr._mcycle_T_2\[30\] _06496_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__or2_1
X_28494_ clknet_leaf_168_clock _01507_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24657_ net1100 execute.io_target_pc\[17\] _08508_ VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__mux2_1
X_27445_ clknet_leaf_147_clock _00474_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21869_ csr.io_mret_vector\[10\] _10878_ _06515_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14410_ net741 _10490_ _10495_ _10494_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__o211a_1
X_23608_ _06138_ net2013 _07941_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15390_ _11194_ decode.regfile.registers_12\[2\] decode.regfile.registers_13\[2\]
+ _11196_ VGND VGND VPWR VPWR _11385_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24588_ _08476_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__clkbuf_1
X_27376_ clknet_leaf_15_clock _00405_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29115_ clknet_leaf_18_clock _02128_ VGND VGND VPWR VPWR csr._mcycle_T_3\[63\] sky130_fd_sc_hd__dfxtp_1
X_14341_ net893 _10447_ _10455_ _10453_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23539_ net2778 _07903_ _07912_ _07907_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26327_ _09383_ _09492_ VGND VGND VPWR VPWR _09498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17060_ _13016_ _12732_ _13017_ VGND VGND VPWR VPWR _13018_ sky130_fd_sc_hd__a21o_1
X_29046_ clknet_leaf_125_clock _02059_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26258_ net480 _09447_ _09457_ _09458_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__o211a_1
X_14272_ _10142_ _10375_ VGND VGND VPWR VPWR _10415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16011_ _11371_ decode.regfile.registers_0\[18\] VGND VGND VPWR VPWR _11990_ sky130_fd_sc_hd__nand2_1
X_25209_ _08833_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26189_ net2418 _09395_ _09411_ _09394_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_223_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ decode.regfile.registers_18\[29\] _12565_ _03339_ _03359_ VGND VGND VPWR
+ VPWR _03360_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_223_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19701_ _04977_ _04974_ _04452_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_29_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16913_ _12852_ VGND VGND VPWR VPWR _12874_ sky130_fd_sc_hd__clkbuf_4
X_17893_ _12515_ _03290_ _03291_ _03292_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__a31o_1
X_29879_ clknet_leaf_300_clock _02892_ VGND VGND VPWR VPWR decode.regfile.registers_19\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19632_ _03912_ _04862_ _04863_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__and3_1
X_16844_ decode.regfile.registers_21\[2\] _12682_ _12806_ VGND VGND VPWR VPWR _12807_
+ sky130_fd_sc_hd__o21a_1
X_19563_ net309 _04371_ _04301_ _04649_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__or4b_1
X_16775_ _12736_ _12738_ VGND VGND VPWR VPWR _12739_ sky130_fd_sc_hd__nand2_1
X_13987_ net2685 _10243_ _10251_ _10249_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18514_ net349 _03809_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_17_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ decode.regfile.registers_20\[10\] _11452_ _11223_ _11712_ VGND VGND VPWR
+ VPWR _11713_ sky130_fd_sc_hd__a211o_1
XFILLER_0_198_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19494_ _04362_ _04767_ _04773_ _04778_ _04779_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_34_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18445_ _03734_ net292 _03743_ _03673_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nand4b_4
X_15657_ _11571_ decode.regfile.registers_30\[9\] _11039_ _11032_ _11033_ VGND VGND
+ VPWR VPWR _11645_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_200_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14608_ _10650_ VGND VGND VPWR VPWR _10651_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_38_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18376_ _09935_ decode.id_ex_ex_rs1_reg\[3\] _03671_ _03673_ _03674_ VGND VGND VPWR
+ VPWR _03675_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_172_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15588_ decode.regfile.registers_1\[7\] _11115_ _11056_ _11108_ VGND VGND VPWR VPWR
+ _11578_ sky130_fd_sc_hd__nand4_1
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17327_ _12499_ _12490_ _12511_ decode.regfile.registers_12\[13\] _12745_ VGND VGND
+ VPWR VPWR _13279_ sky130_fd_sc_hd__o32a_1
XFILLER_0_172_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14539_ decode.control.io_funct3\[1\] decode.control.io_funct3\[0\] _10581_ VGND
+ VGND VPWR VPWR _10582_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_56_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17258_ _13087_ decode.regfile.registers_26\[11\] _12814_ _13047_ _13088_ VGND VGND
+ VPWR VPWR _13212_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_77_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16209_ _12181_ _11533_ _12182_ VGND VGND VPWR VPWR _12183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17189_ decode.regfile.registers_1\[10\] _12778_ _12830_ _13143_ VGND VGND VPWR VPWR
+ _13144_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_11_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2504 decode.regfile.registers_16\[25\] VGND VGND VPWR VPWR net2731 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2515 decode.regfile.registers_9\[6\] VGND VGND VPWR VPWR net2742 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2526 decode.regfile.registers_0\[11\] VGND VGND VPWR VPWR net2753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2537 decode.csr_read_reg VGND VGND VPWR VPWR net2764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1803 fetch.bht.bhtTable_tag\[15\]\[7\] VGND VGND VPWR VPWR net2030 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2548 csr._mcycle_T_2\[7\] VGND VGND VPWR VPWR net2775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1814 fetch.bht.bhtTable_target_pc\[15\]\[4\] VGND VGND VPWR VPWR net2041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2559 net68 VGND VGND VPWR VPWR net2786 sky130_fd_sc_hd__dlygate4sd3_1
X_22910_ net80 _06833_ _06767_ net224 _06893_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__a221oi_1
Xhold1825 decode.regfile.registers_9\[19\] VGND VGND VPWR VPWR net2052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1836 decode.regfile.registers_22\[7\] VGND VGND VPWR VPWR net2063 sky130_fd_sc_hd__dlygate4sd3_1
X_23890_ _08114_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1847 fetch.bht.bhtTable_tag\[11\]\[11\] VGND VGND VPWR VPWR net2074 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1858 decode.regfile.registers_17\[2\] VGND VGND VPWR VPWR net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1869 csr._csr_read_data_T_8\[12\] VGND VGND VPWR VPWR net2096 sky130_fd_sc_hd__dlygate4sd3_1
X_22841_ _07316_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25560_ _08935_ _09036_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22772_ _07279_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24511_ _08436_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21723_ net2797 _06321_ _06420_ csr.minstret\[31\] VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_56_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25491_ decode.regfile.registers_2\[16\] _08995_ _09002_ _08991_ VGND VGND VPWR VPWR
+ _02335_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24442_ _08388_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_176_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27230_ clknet_leaf_2_clock _00259_ VGND VGND VPWR VPWR decode.regfile.registers_29\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_21654_ _05691_ _06366_ _06367_ _06352_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_163_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20605_ _05540_ csr.io_mret_vector\[23\] _05565_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__o21a_1
X_27161_ clknet_leaf_360_clock _00190_ VGND VGND VPWR VPWR decode.regfile.registers_27\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24373_ _08363_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21585_ csr.io_csr_write_address\[10\] csr.io_csr_write_address\[8\] csr.io_csr_write_address\[9\]
+ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__and3b_2
XFILLER_0_201_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26112_ _08958_ _09353_ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__nand2_1
X_23324_ fetch.bht.bhtTable_target_pc\[0\]\[25\] fetch.bht.bhtTable_target_pc\[1\]\[25\]
+ fetch.bht.bhtTable_target_pc\[2\]\[25\] fetch.bht.bhtTable_target_pc\[3\]\[25\]
+ _07098_ _07113_ VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20536_ csr.minstret\[13\] _05574_ _05586_ csr.mcycle\[13\] _05682_ VGND VGND VPWR
+ VPWR _05683_ sky130_fd_sc_hd__a221o_1
X_27092_ clknet_leaf_329_clock _00121_ VGND VGND VPWR VPWR decode.regfile.registers_25\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26043_ _08964_ _09310_ VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__nand2_1
X_23255_ net79 _07536_ _07537_ _07687_ _07535_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__o311a_1
XFILLER_0_104_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20467_ _05618_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__buf_4
XFILLER_0_162_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22206_ _06629_ _06796_ _06800_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_65_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23186_ fetch.bht.bhtTable_target_pc\[12\]\[17\] fetch.bht.bhtTable_target_pc\[13\]\[17\]
+ fetch.bht.bhtTable_target_pc\[14\]\[17\] fetch.bht.bhtTable_target_pc\[15\]\[17\]
+ _07384_ _07113_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__mux4_1
XFILLER_0_219_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20398_ _05540_ _05554_ csr.io_mret_vector\[0\] _05556_ _05557_ VGND VGND VPWR VPWR
+ _05558_ sky130_fd_sc_hd__o311a_1
XFILLER_0_219_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29802_ clknet_leaf_297_clock _02815_ VGND VGND VPWR VPWR decode.regfile.registers_17\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22137_ fetch.bht.bhtTable_tag\[4\]\[4\] fetch.bht.bhtTable_tag\[5\]\[4\] net302
+ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__mux2_1
X_27994_ clknet_leaf_236_clock _01016_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29733_ clknet_leaf_285_clock _02746_ VGND VGND VPWR VPWR decode.regfile.registers_15\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_22068_ _06659_ _06660_ _06661_ _06662_ _06633_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__o221a_1
XFILLER_0_206_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26945_ net659 _09853_ _09854_ _09852_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13910_ net2324 _10199_ _10205_ _10206_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__o211a_1
X_21019_ execute.csr_read_data_out_reg\[0\] _05989_ _05985_ VGND VGND VPWR VPWR _05994_
+ sky130_fd_sc_hd__and3_1
X_29664_ clknet_leaf_287_clock _02677_ VGND VGND VPWR VPWR decode.regfile.registers_13\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14890_ _10926_ VGND VGND VPWR VPWR _10927_ sky130_fd_sc_hd__buf_2
X_26876_ net1548 _09809_ _09814_ _09812_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28615_ clknet_leaf_115_clock _01628_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13841_ net511 _10153_ _10165_ _10162_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__o211a_1
X_25827_ _08975_ _09155_ VGND VGND VPWR VPWR _09196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29595_ clknet_leaf_270_clock _02608_ VGND VGND VPWR VPWR decode.regfile.registers_11\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_28546_ clknet_leaf_166_clock _01559_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16560_ _12524_ VGND VGND VPWR VPWR _12525_ sky130_fd_sc_hd__clkbuf_4
X_13772_ _10111_ VGND VGND VPWR VPWR _10112_ sky130_fd_sc_hd__clkbuf_8
X_25758_ _09025_ _09157_ VGND VGND VPWR VPWR _09158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15511_ _11129_ VGND VGND VPWR VPWR _11503_ sky130_fd_sc_hd__buf_4
XFILLER_0_35_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24709_ _08538_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28477_ clknet_leaf_236_clock _01490_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16491_ _11300_ decode.regfile.registers_0\[31\] VGND VGND VPWR VPWR _12457_ sky130_fd_sc_hd__nand2_1
X_25689_ net1710 _09111_ _09117_ _09115_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18230_ csr.mcycle\[28\] csr.mcycle\[27\] _03564_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_216_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15442_ _11435_ VGND VGND VPWR VPWR _11436_ sky130_fd_sc_hd__clkbuf_4
X_27428_ clknet_leaf_40_clock _00457_ VGND VGND VPWR VPWR decode.id_ex_memtoreg_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18161_ _11062_ _10577_ _10673_ _10911_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__nor4_1
X_15373_ decode.regfile.registers_3\[2\] _11292_ _11367_ _11178_ VGND VGND VPWR VPWR
+ _11368_ sky130_fd_sc_hd__o2bb2a_1
X_27359_ clknet_leaf_33_clock _00388_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17112_ decode.regfile.registers_12\[8\] _12794_ _13067_ _13068_ _12775_ VGND VGND
+ VPWR VPWR _13069_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_894 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14324_ _10081_ _10444_ VGND VGND VPWR VPWR _10446_ sky130_fd_sc_hd__nand2_1
X_18092_ _03469_ _03467_ _03465_ net2213 VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_123_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29029_ clknet_leaf_139_clock _02042_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17043_ _12759_ VGND VGND VPWR VPWR _13002_ sky130_fd_sc_hd__clkbuf_4
X_14255_ _10097_ _10400_ VGND VGND VPWR VPWR _10406_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14186_ net1066 _10359_ _10365_ _10357_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18994_ _04245_ _04271_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_104_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17945_ _12387_ _12932_ _10615_ _12933_ _03342_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_218_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17876_ decode.regfile.registers_8\[27\] _12725_ _03268_ _03275_ VGND VGND VPWR VPWR
+ _03276_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_105_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19615_ _03918_ _03934_ _04253_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__mux2_1
X_16827_ _12652_ VGND VGND VPWR VPWR _12790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19546_ _04745_ _04828_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__nand2_2
X_16758_ _12721_ VGND VGND VPWR VPWR _12722_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15709_ _11129_ _11298_ _11300_ decode.regfile.registers_0\[10\] VGND VGND VPWR VPWR
+ _11696_ sky130_fd_sc_hd__a2bb2o_1
X_19477_ _04119_ _04742_ _04107_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_61_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16689_ _12653_ VGND VGND VPWR VPWR _12654_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_330 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_341 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_352 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18428_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__buf_4
XINSDIODE1_363 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_374 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_385 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18359_ _03657_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_135_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21370_ _06197_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20321_ _05417_ _05367_ _05492_ _05454_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__o211a_1
Xhold900 fetch.bht.bhtTable_tag\[12\]\[5\] VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold911 decode.regfile.registers_11\[15\] VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold922 decode.regfile.registers_5\[14\] VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__dlygate4sd3_1
X_23040_ csr._csr_read_data_T_8\[8\] _06038_ csr.io_mret_vector\[8\] _06462_ VGND
+ VGND VPWR VPWR _07485_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20252_ _10910_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__clkbuf_4
Xhold933 decode.regfile.registers_17\[7\] VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold944 fetch.bht.bhtTable_tag\[11\]\[6\] VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 _08479_ VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 fetch.bht.bhtTable_target_pc\[11\]\[31\] VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold977 fetch.bht.bhtTable_tag\[1\]\[3\] VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold988 fetch.bht.bhtTable_tag\[0\]\[1\] VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__dlygate4sd3_1
X_20183_ _05382_ _05383_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_34_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold999 fetch.bht.bhtTable_target_pc\[11\]\[4\] VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2301 decode.regfile.registers_2\[30\] VGND VGND VPWR VPWR net2528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2312 decode.regfile.registers_19\[14\] VGND VGND VPWR VPWR net2539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2323 decode.regfile.registers_4\[18\] VGND VGND VPWR VPWR net2550 sky130_fd_sc_hd__dlygate4sd3_1
X_24991_ _08701_ csr.mcycle\[1\] csr.mcycle\[0\] csr.mcycle\[2\] VGND VGND VPWR VPWR
+ _08707_ sky130_fd_sc_hd__a31o_1
Xhold2334 csr._mcycle_T_3\[59\] VGND VGND VPWR VPWR net2561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1600 fetch.bht.bhtTable_target_pc\[7\]\[12\] VGND VGND VPWR VPWR net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2345 decode.regfile.registers_5\[6\] VGND VGND VPWR VPWR net2572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1611 fetch.bht.bhtTable_target_pc\[10\]\[9\] VGND VGND VPWR VPWR net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2356 execute.io_reg_pc\[14\] VGND VGND VPWR VPWR net2583 sky130_fd_sc_hd__dlygate4sd3_1
X_26730_ net749 _09723_ _09729_ _09730_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23942_ _08141_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__clkbuf_1
Xhold1622 fetch.bht.bhtTable_tag\[0\]\[23\] VGND VGND VPWR VPWR net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2367 decode.regfile.registers_4\[25\] VGND VGND VPWR VPWR net2594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 fetch.bht.bhtTable_target_pc\[10\]\[11\] VGND VGND VPWR VPWR net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2378 decode.regfile.registers_3\[28\] VGND VGND VPWR VPWR net2605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1644 net91 VGND VGND VPWR VPWR net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2389 csr._mcycle_T_3\[46\] VGND VGND VPWR VPWR net2616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1655 fetch.bht.bhtTable_tag\[6\]\[13\] VGND VGND VPWR VPWR net1882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23873_ execute.io_target_pc\[26\] VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__clkbuf_2
Xhold1666 fetch.bht.bhtTable_tag\[0\]\[18\] VGND VGND VPWR VPWR net1893 sky130_fd_sc_hd__dlygate4sd3_1
X_26661_ net2710 _09679_ _09690_ _09688_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__o211a_1
Xhold1677 fetch.bht.bhtTable_tag\[13\]\[21\] VGND VGND VPWR VPWR net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1688 decode.regfile.registers_17\[23\] VGND VGND VPWR VPWR net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1699 fetch.bht.bhtTable_target_pc\[10\]\[22\] VGND VGND VPWR VPWR net1926 sky130_fd_sc_hd__dlygate4sd3_1
X_28400_ clknet_leaf_142_clock _01413_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_2
X_22824_ _07307_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__clkbuf_1
X_25612_ _08912_ _09069_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29380_ clknet_leaf_257_clock _02393_ VGND VGND VPWR VPWR decode.regfile.registers_4\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_26592_ _09422_ _09645_ VGND VGND VPWR VPWR _09651_ sky130_fd_sc_hd__nand2_1
X_28331_ clknet_leaf_166_clock _01344_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_22755_ _07270_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25543_ net656 _09024_ _09032_ _09033_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21706_ csr.minstret\[14\] _06333_ _06355_ _06360_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__and4_1
XFILLER_0_164_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28262_ clknet_leaf_77_clock _01284_ VGND VGND VPWR VPWR csr._minstret_T_3\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_25474_ net2745 _08979_ _08993_ _08991_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22686_ net2256 _07222_ _07230_ _07221_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24425_ _08391_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27213_ clknet_leaf_3_clock _00242_ VGND VGND VPWR VPWR decode.regfile.registers_28\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21637_ _05613_ csr.minstret\[5\] csr.minstret\[10\] VGND VGND VPWR VPWR _06354_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_229_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28193_ clknet_leaf_112_clock _01215_ VGND VGND VPWR VPWR csr.io_mret_vector\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_229_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24356_ _08354_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27144_ clknet_leaf_358_clock _00173_ VGND VGND VPWR VPWR decode.regfile.registers_26\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21568_ _06304_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23307_ fetch.bht.bhtTable_target_pc\[12\]\[24\] fetch.bht.bhtTable_target_pc\[13\]\[24\]
+ fetch.bht.bhtTable_target_pc\[14\]\[24\] fetch.bht.bhtTable_target_pc\[15\]\[24\]
+ _07555_ _07710_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_185_Right_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20519_ csr.minstret\[11\] _05594_ _05595_ csr._minstret_T_3\[43\] VGND VGND VPWR
+ VPWR _05668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27075_ clknet_leaf_346_clock _00104_ VGND VGND VPWR VPWR decode.regfile.registers_24\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_24287_ _08049_ net1532 _06210_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21499_ _06128_ net1726 _06263_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14040_ _10128_ _10242_ VGND VGND VPWR VPWR _10281_ sky130_fd_sc_hd__nand2_1
X_23238_ _07659_ _07664_ _07671_ _07088_ VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26026_ decode.regfile.registers_9\[18\] _09300_ _09311_ _09305_ VGND VGND VPWR VPWR
+ _02561_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23169_ fetch.bht.bhtTable_target_pc\[10\]\[16\] fetch.bht.bhtTable_target_pc\[11\]\[16\]
+ _07108_ VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_207_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27977_ clknet_leaf_193_clock _00999_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15991_ _11106_ _11969_ _11970_ VGND VGND VPWR VPWR _11971_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17730_ decode.regfile.registers_19\[23\] _12678_ _03112_ _03133_ _12906_ VGND VGND
+ VPWR VPWR _03134_ sky130_fd_sc_hd__o221a_1
X_29716_ clknet_leaf_283_clock _02729_ VGND VGND VPWR VPWR decode.regfile.registers_14\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14942_ csr.io_trapped _10970_ VGND VGND VPWR VPWR _10971_ sky130_fd_sc_hd__or2_2
X_26928_ net1348 _09839_ _09844_ _09836_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_82_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17661_ _13183_ _03064_ _03065_ _03066_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__a31o_1
X_29647_ clknet_leaf_279_clock _02660_ VGND VGND VPWR VPWR decode.regfile.registers_12\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14873_ _10914_ VGND VGND VPWR VPWR _10915_ sky130_fd_sc_hd__clkbuf_4
X_26859_ net1681 _09795_ _09804_ _09799_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19400_ _04168_ _04682_ _04688_ _04505_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16612_ _10594_ _10598_ _10588_ _12511_ VGND VGND VPWR VPWR _12577_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_218_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ _09964_ _10154_ VGND VGND VPWR VPWR _10156_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_218_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17592_ decode.regfile.registers_15\[20\] _12555_ _10923_ _12876_ _13031_ VGND VGND
+ VPWR VPWR _02999_ sky130_fd_sc_hd__a41o_1
X_29578_ clknet_leaf_267_clock _02591_ VGND VGND VPWR VPWR decode.regfile.registers_10\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19331_ _04045_ _04234_ _04247_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28529_ clknet_leaf_234_clock _01542_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16543_ _10614_ VGND VGND VPWR VPWR _12508_ sky130_fd_sc_hd__buf_4
X_13755_ _10097_ _10075_ VGND VGND VPWR VPWR _10098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19262_ _04541_ _04393_ _04555_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16474_ decode.regfile.registers_21\[30\] _11267_ _11099_ _11228_ _12440_ VGND VGND
+ VPWR VPWR _12441_ sky130_fd_sc_hd__o311a_1
XFILLER_0_39_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13686_ _09943_ memory.io_wb_readdata\[12\] _10038_ VGND VGND VPWR VPWR _10039_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18213_ net2783 _11100_ _03548_ _03549_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__or4_1
XFILLER_0_156_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15425_ _11408_ _11417_ _11418_ VGND VGND VPWR VPWR _11419_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_183_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19193_ _04332_ _04486_ _04461_ _04317_ _04488_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__o311a_1
XFILLER_0_66_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18144_ _03501_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_91_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15356_ _11347_ _11348_ decode.regfile.registers_26\[2\] _11349_ _11350_ VGND VGND
+ VPWR VPWR _11351_ sky130_fd_sc_hd__a41o_1
XFILLER_0_198_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14307_ net554 _10434_ _10436_ _10427_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__o211a_1
Xwire171 _00677_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18075_ _10579_ _10667_ _10973_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15287_ _10645_ _10627_ _10635_ _11069_ VGND VGND VPWR VPWR _11283_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_169_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold207 decode.regfile.registers_31\[7\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 decode.regfile.registers_31\[29\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__buf_1
Xhold229 decode.regfile.registers_27\[31\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ _11020_ _12491_ _12666_ decode.regfile.registers_14\[6\] _12984_ VGND VGND
+ VPWR VPWR _12985_ sky130_fd_sc_hd__o32a_1
X_14238_ _10058_ _10387_ VGND VGND VPWR VPWR _10396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14169_ _10074_ _10355_ VGND VGND VPWR VPWR _10356_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _03835_ _03844_ _04230_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ decode.regfile.registers_21\[28\] _12682_ _03304_ _03326_ _12806_ VGND VGND
+ VPWR VPWR _03327_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17859_ _10929_ decode.regfile.registers_28\[26\] _02992_ VGND VGND VPWR VPWR _03260_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_124_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20870_ net121 _05903_ _05911_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19529_ _04251_ _04252_ _04768_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22540_ _06041_ _07133_ _06481_ _07065_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_27_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_160 _13356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_171 decode.id_ex_rs1_data_reg\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_182 execute.io_reg_pc\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_193 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22471_ _06619_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_1084 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24210_ _08279_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21422_ _06113_ net1314 _06219_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25190_ _09883_ _08813_ _09881_ VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24141_ net966 execute.io_target_pc\[25\] _06427_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__mux2_1
X_21353_ _06101_ net1077 _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20304_ _05340_ _05473_ _10867_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__a21oi_1
X_24072_ _08208_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21284_ csr.io_mem_pc\[29\] VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__buf_2
XFILLER_0_124_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold730 memory.csr_read_data_out_reg\[5\] VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__buf_1
Xhold741 _08237_ VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold752 _08163_ VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23023_ execute.io_target_pc\[7\] _05857_ _07091_ _07468_ _07347_ VGND VGND VPWR
+ VPWR _07469_ sky130_fd_sc_hd__a311oi_1
X_27900_ clknet_leaf_18_clock _00929_ VGND VGND VPWR VPWR csr._mcycle_T_2\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold763 fetch.bht.bhtTable_target_pc\[4\]\[31\] VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20235_ _05426_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__clkbuf_1
Xhold774 fetch.bht.bhtTable_target_pc\[4\]\[24\] VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__dlygate4sd3_1
X_28880_ clknet_leaf_120_clock _01893_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold785 fetch.bht.bhtTable_tag\[2\]\[8\] VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 _08168_ VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27831_ clknet_leaf_320_clock _00860_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20166_ decode.id_ex_imm_reg\[24\] decode.id_ex_pc_reg\[24\] VGND VGND VPWR VPWR
+ _05369_ sky130_fd_sc_hd__nand2_1
Xhold2120 csr._mcycle_T_3\[48\] VGND VGND VPWR VPWR net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2131 execute.csr_write_data_out_reg\[12\] VGND VGND VPWR VPWR net2358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2142 decode.regfile.registers_3\[27\] VGND VGND VPWR VPWR net2369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27762_ clknet_leaf_316_clock _00791_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2153 decode.regfile.registers_8\[16\] VGND VGND VPWR VPWR net2380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2164 _01241_ VGND VGND VPWR VPWR net2391 sky130_fd_sc_hd__dlygate4sd3_1
X_20097_ _05308_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__and2b_1
X_24974_ csr._mcycle_T_3\[60\] csr._mcycle_T_3\[59\] _08693_ VGND VGND VPWR VPWR _08696_
+ sky130_fd_sc_hd__and3_1
Xhold2175 csr._csr_read_data_T_8\[25\] VGND VGND VPWR VPWR net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29501_ clknet_leaf_251_clock _02514_ VGND VGND VPWR VPWR decode.regfile.registers_8\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1430 decode.regfile.registers_5\[16\] VGND VGND VPWR VPWR net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 fetch.bht.bhtTable_target_pc\[9\]\[26\] VGND VGND VPWR VPWR net1668 sky130_fd_sc_hd__dlygate4sd3_1
X_26713_ _09389_ _09720_ VGND VGND VPWR VPWR _09721_ sky130_fd_sc_hd__nand2_1
Xhold2186 decode.regfile.registers_8\[3\] VGND VGND VPWR VPWR net2413 sky130_fd_sc_hd__dlygate4sd3_1
X_23925_ net1272 _08083_ _08130_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__mux2_1
Xhold1452 fetch.bht.bhtTable_target_pc\[5\]\[17\] VGND VGND VPWR VPWR net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2197 decode.regfile.registers_15\[27\] VGND VGND VPWR VPWR net2424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1463 decode.regfile.registers_8\[7\] VGND VGND VPWR VPWR net1690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27693_ clknet_leaf_26_clock _00722_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1474 fetch.bht.bhtTable_target_pc\[14\]\[5\] VGND VGND VPWR VPWR net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1485 fetch.bht.bhtTable_target_pc\[3\]\[4\] VGND VGND VPWR VPWR net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29432_ clknet_leaf_247_clock _02445_ VGND VGND VPWR VPWR decode.regfile.registers_5\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_200_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 decode.regfile.registers_19\[17\] VGND VGND VPWR VPWR net1723 sky130_fd_sc_hd__dlygate4sd3_1
X_26644_ _09398_ _09676_ VGND VGND VPWR VPWR _09681_ sky130_fd_sc_hd__nand2_1
X_23856_ _08091_ net1073 _08079_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22807_ net959 _10803_ _07297_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__mux2_1
X_29363_ clknet_leaf_227_clock _02376_ VGND VGND VPWR VPWR decode.regfile.registers_3\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26575_ _09404_ _09632_ VGND VGND VPWR VPWR _09641_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23787_ _06149_ net1919 _08041_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20999_ execute.io_reg_pc\[24\] _05977_ _05973_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28314_ clknet_leaf_212_clock _01327_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13540_ csr.io_mem_pc\[5\] _09879_ VGND VGND VPWR VPWR _09915_ sky130_fd_sc_hd__and2b_1
X_25526_ _10150_ _03672_ _08903_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22738_ _07261_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__clkbuf_1
X_29294_ clknet_leaf_225_clock _02307_ VGND VGND VPWR VPWR decode.regfile.registers_1\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28245_ clknet_leaf_77_clock _01267_ VGND VGND VPWR VPWR csr._minstret_T_3\[45\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22669_ _06578_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__buf_2
XFILLER_0_137_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25457_ net1558 _08979_ _08983_ _08972_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15210_ _11206_ VGND VGND VPWR VPWR _11207_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24408_ _08381_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__clkbuf_1
X_28176_ clknet_leaf_57_clock _01198_ VGND VGND VPWR VPWR csr.io_mret_vector\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16190_ _11075_ _12163_ _12164_ _11236_ VGND VGND VPWR VPWR _12165_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25388_ _10047_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_11_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_998 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27127_ clknet_leaf_356_clock _00156_ VGND VGND VPWR VPWR decode.regfile.registers_26\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_15141_ _11091_ _10623_ _11137_ VGND VGND VPWR VPWR _11138_ sky130_fd_sc_hd__and3_2
X_24339_ _08101_ net2059 _06187_ VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15072_ _10654_ _10659_ VGND VGND VPWR VPWR _11069_ sky130_fd_sc_hd__nor2b_2
X_27058_ clknet_leaf_330_clock _00087_ VGND VGND VPWR VPWR decode.regfile.registers_24\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14023_ _10087_ _10268_ VGND VGND VPWR VPWR _10272_ sky130_fd_sc_hd__nand2_1
X_18900_ decode.id_ex_rs1_data_reg\[18\] _03908_ _03913_ _03700_ _03917_ VGND VGND
+ VPWR VPWR _04199_ sky130_fd_sc_hd__o221ai_4
X_26009_ _08931_ _09297_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19880_ _03802_ _05128_ _03791_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_207_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18831_ _04126_ _04129_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_160_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18762_ decode.id_ex_rs1_data_reg\[7\] _03908_ _04060_ _03914_ VGND VGND VPWR VPWR
+ _04061_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_199_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15974_ decode.regfile.registers_1\[17\] _11116_ _11056_ _11108_ VGND VGND VPWR VPWR
+ _11954_ sky130_fd_sc_hd__nand4_1
XFILLER_0_101_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17713_ decode.regfile.registers_4\[23\] decode.regfile.registers_5\[23\] _12882_
+ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__mux2_1
X_14925_ _10953_ VGND VGND VPWR VPWR _10954_ sky130_fd_sc_hd__clkbuf_2
X_18693_ execute.csr_read_data_out_reg\[1\] execute.io_mem_memtoreg\[0\] execute.io_mem_memtoreg\[1\]
+ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_215_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17644_ decode.regfile.registers_12\[21\] _12489_ _11019_ _12541_ VGND VGND VPWR
+ VPWR _03050_ sky130_fd_sc_hd__or4_1
X_14856_ decode.id_ex_pc_reg\[14\] _10877_ _10880_ _10694_ _10898_ VGND VGND VPWR
+ VPWR _10899_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_72_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13807_ _10141_ VGND VGND VPWR VPWR _10142_ sky130_fd_sc_hd__buf_4
X_17575_ _13250_ decode.regfile.registers_24\[19\] _13170_ _13083_ _13367_ VGND VGND
+ VPWR VPWR _02983_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_221_Right_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14787_ decode.id_ex_pc_reg\[0\] csr.io_mem_pc\[0\] VGND VGND VPWR VPWR _10830_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19314_ _04279_ _04019_ _04473_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_202_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16526_ _12490_ VGND VGND VPWR VPWR _12491_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13738_ _09937_ VGND VGND VPWR VPWR _10083_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19245_ _04492_ _04536_ _04538_ _04539_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__a22o_1
X_16457_ _11300_ decode.regfile.registers_0\[30\] _11155_ _12423_ VGND VGND VPWR VPWR
+ _12424_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13669_ _10024_ VGND VGND VPWR VPWR _10025_ sky130_fd_sc_hd__buf_4
XFILLER_0_183_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_213_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15408_ _10962_ net2126 _11039_ _11032_ _11033_ VGND VGND VPWR VPWR _11402_ sky130_fd_sc_hd__o2111a_1
X_19176_ _04364_ _04351_ _04277_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16388_ _12351_ _12355_ _12356_ VGND VGND VPWR VPWR _12357_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18127_ _03491_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15339_ _11334_ VGND VGND VPWR VPWR _11335_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_182_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18058_ _03450_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17009_ _12694_ VGND VGND VPWR VPWR _12968_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20020_ _04018_ _10711_ _05243_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21971_ _06573_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer11 net237 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23710_ net1365 csr.io_mem_pc\[18\] _08003_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__mux2_1
X_20922_ _05941_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer22 _03686_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24690_ _08528_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer33 _03739_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_1
XFILLER_0_96_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer44 net205 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__buf_6
Xrebuffer55 _10765_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer66 _03710_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_222_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23641_ _07968_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20853_ net465 _05903_ _05899_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__and3_1
Xrebuffer77 _03752_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_1
Xrebuffer88 _03745_ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__buf_6
XFILLER_0_178_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer99 _03752_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__buf_1
XFILLER_0_193_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23572_ _06103_ net1563 _07930_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__mux2_1
X_26360_ _09415_ _09515_ VGND VGND VPWR VPWR _09517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20784_ _05865_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22523_ _07115_ _07116_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__and2b_1
XFILLER_0_181_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25311_ _08880_ decode.regfile.registers_0\[17\] VGND VGND VPWR VPWR _08886_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_46_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26291_ net2376 _09475_ _09477_ _09471_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28030_ clknet_leaf_198_clock _01052_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[6\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25242_ _08081_ net1612 _08848_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__mux2_1
X_22454_ _06617_ fetch.btb.btbTable\[12\]\[1\] fetch.bht.bhtTable_valid\[12\] VGND
+ VGND VPWR VPWR _07049_ sky130_fd_sc_hd__and3b_1
Xrebuffer101 net327 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer112 _05041_ VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_91_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21405_ _06153_ net2118 _06210_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25173_ _08815_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22385_ _06622_ _06979_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_59_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24124_ _08235_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__clkbuf_1
X_21336_ _06178_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__clkbuf_1
X_24055_ net900 execute.io_target_pc\[15\] _08198_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__mux2_1
X_28932_ clknet_leaf_130_clock _01945_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_21267_ _06137_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__clkbuf_1
Xhold560 fetch.bht.bhtTable_tag\[3\]\[16\] VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold571 fetch.bht.bhtTable_tag\[2\]\[19\] VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23006_ _06248_ _07450_ _07452_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold582 decode.regfile.registers_23\[0\] VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__dlygate4sd3_1
X_20218_ _05223_ _05224_ _05412_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__o21ai_1
Xhold593 decode.regfile.registers_5\[12\] VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__dlygate4sd3_1
X_28863_ clknet_leaf_181_clock _01876_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21198_ _06094_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27814_ clknet_leaf_325_clock _00843_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_202_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20149_ _05352_ _05354_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__xnor2_1
X_28794_ clknet_leaf_129_clock _01807_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_202_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_216_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27745_ clknet_leaf_326_clock _00774_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_24957_ csr._mcycle_T_3\[54\] csr._mcycle_T_3\[53\] _08682_ VGND VGND VPWR VPWR _08685_
+ sky130_fd_sc_hd__and3_1
Xhold1260 fetch.bht.bhtTable_tag\[13\]\[17\] VGND VGND VPWR VPWR net1487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14710_ _10743_ execute.io_target_pc\[28\] _10745_ _10752_ VGND VGND VPWR VPWR _10753_
+ sky130_fd_sc_hd__o211a_1
Xhold1271 fetch.bht.bhtTable_tag\[8\]\[2\] VGND VGND VPWR VPWR net1498 sky130_fd_sc_hd__dlygate4sd3_1
X_23908_ net1024 _08066_ _08119_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__mux2_1
Xhold1282 fetch.bht.bhtTable_target_pc\[8\]\[18\] VGND VGND VPWR VPWR net1509 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_194_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _11236_ _11674_ _11675_ _11677_ VGND VGND VPWR VPWR _11678_ sky130_fd_sc_hd__a31o_1
Xhold1293 decode.regfile.registers_23\[4\] VGND VGND VPWR VPWR net1520 sky130_fd_sc_hd__dlygate4sd3_1
X_27676_ clknet_leaf_30_clock _00705_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_24888_ net1800 _08636_ _08637_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__o21a_1
X_29415_ clknet_leaf_257_clock _02428_ VGND VGND VPWR VPWR decode.regfile.registers_5\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14641_ decode.id_ex_pc_reg\[30\] VGND VGND VPWR VPWR _10684_ sky130_fd_sc_hd__inv_2
X_26627_ _09381_ _09666_ VGND VGND VPWR VPWR _09671_ sky130_fd_sc_hd__nand2_1
X_23839_ _08080_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29346_ clknet_leaf_256_clock _02359_ VGND VGND VPWR VPWR decode.regfile.registers_3\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_17360_ decode.regfile.registers_4\[14\] _12617_ _12619_ decode.regfile.registers_5\[14\]
+ _12622_ VGND VGND VPWR VPWR _13311_ sky130_fd_sc_hd__a221oi_1
X_26558_ _09387_ _09623_ VGND VGND VPWR VPWR _09631_ sky130_fd_sc_hd__nand2_1
X_14572_ _10614_ VGND VGND VPWR VPWR _10615_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_354_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_354_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16311_ decode.regfile.registers_3\[26\] _11614_ _11367_ _11178_ VGND VGND VPWR VPWR
+ _12282_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_32_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13523_ _09900_ _09880_ _09883_ _09887_ VGND VGND VPWR VPWR _09901_ sky130_fd_sc_hd__or4bb_4
X_25509_ _08960_ _09005_ VGND VGND VPWR VPWR _09013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29277_ clknet_leaf_241_clock _02290_ VGND VGND VPWR VPWR decode.regfile.registers_1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_17291_ decode.regfile.registers_18\[12\] _10924_ _12568_ _12524_ _11008_ VGND VGND
+ VPWR VPWR _13244_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26489_ net623 _09578_ _09591_ _09582_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_153_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19030_ _04325_ _04326_ _04328_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__a21oi_2
X_28228_ clknet_leaf_83_clock _01250_ VGND VGND VPWR VPWR csr.mscratch\[30\] sky130_fd_sc_hd__dfxtp_1
X_16242_ _12207_ _12214_ _11175_ VGND VGND VPWR VPWR _12215_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28159_ clknet_leaf_66_clock _01181_ VGND VGND VPWR VPWR csr.meie sky130_fd_sc_hd__dfxtp_1
X_16173_ decode.regfile.registers_9\[22\] _11280_ _11134_ _11509_ VGND VGND VPWR VPWR
+ _12148_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_209_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15124_ _11120_ VGND VGND VPWR VPWR _11121_ sky130_fd_sc_hd__clkbuf_8
Xoutput109 net109 VGND VGND VPWR VPWR io_memory_address[18] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_112_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19932_ _05199_ _04855_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__nand2_4
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15055_ _11051_ VGND VGND VPWR VPWR _11052_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_112_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14006_ net1220 _10258_ _10261_ _10262_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__o211a_1
X_19863_ _04883_ _05113_ _05114_ _05133_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_183_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput80 net80 VGND VGND VPWR VPWR io_fetch_address[21] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput91 net91 VGND VGND VPWR VPWR io_fetch_address[31] sky130_fd_sc_hd__clkbuf_4
X_18814_ _03759_ _04110_ decode.id_ex_rs2_data_reg\[12\] net315 _03726_ VGND VGND
+ VPWR VPWR _04113_ sky130_fd_sc_hd__o221a_1
X_19794_ net339 _05043_ _05067_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18745_ _03656_ _04041_ _03669_ _04043_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__o211a_1
X_15957_ _11075_ _11936_ _11937_ _11236_ VGND VGND VPWR VPWR _11938_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_307_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_307_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_121_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14908_ _10940_ _10577_ _10673_ _10911_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__nor4_1
XFILLER_0_204_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18676_ _03706_ decode.id_ex_imm_reg\[3\] _03972_ _03974_ VGND VGND VPWR VPWR _03975_
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_204_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15888_ _11066_ VGND VGND VPWR VPWR _11871_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_86_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17627_ decode.regfile.registers_15\[21\] _10612_ _10619_ _12589_ _13031_ VGND VGND
+ VPWR VPWR _03033_ sky130_fd_sc_hd__a41o_1
X_14839_ _10881_ _10817_ _10816_ _10878_ VGND VGND VPWR VPWR _10882_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17558_ _02963_ _02964_ _02965_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__a21o_1
XFILLER_0_175_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16509_ decode.regfile.registers_19\[31\] _11406_ _11325_ _12474_ VGND VGND VPWR
+ VPWR _12475_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_119_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17489_ _12719_ _13436_ VGND VGND VPWR VPWR _13437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19228_ _03638_ _04504_ _04039_ _04522_ _04308_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__o311a_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19159_ _04024_ _04455_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_41_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22170_ fetch.bht.bhtTable_tag\[8\]\[13\] fetch.bht.bhtTable_tag\[9\]\[13\] fetch.bht.bhtTable_tag\[10\]\[13\]
+ fetch.bht.bhtTable_tag\[11\]\[13\] _06754_ _06622_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21121_ _06050_ _06046_ net825 VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21052_ execute.csr_read_data_out_reg\[15\] _06002_ _06010_ VGND VGND VPWR VPWR _06012_
+ sky130_fd_sc_hd__and3_1
X_20003_ _04261_ decode.id_ex_pc_reg\[1\] VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__xnor2_1
X_25860_ _08933_ _09210_ VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__nand2_1
X_24811_ _08592_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25791_ _08939_ _09166_ VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27530_ clknet_leaf_155_clock _00559_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_2_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24742_ _08555_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21954_ _06578_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27461_ clknet_leaf_137_clock _00490_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20905_ _05925_ _05921_ net38 VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__and3_1
X_24673_ net1465 execute.io_target_pc\[25\] _07285_ VGND VGND VPWR VPWR _08520_ sky130_fd_sc_hd__mux2_1
X_21885_ net806 _06521_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29200_ clknet_leaf_240_clock _02213_ VGND VGND VPWR VPWR fetch.btb.btbTable\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26412_ _09392_ _09545_ VGND VGND VPWR VPWR _09547_ sky130_fd_sc_hd__nand2_1
X_23624_ _07958_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__clkbuf_1
X_20836_ _05894_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27392_ clknet_leaf_31_clock _00421_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29131_ clknet_leaf_82_clock _02144_ VGND VGND VPWR VPWR csr.mcycle\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_194_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26343_ net612 _09505_ _09507_ _09499_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_13_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23555_ net2298 _07918_ _07915_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__or3b_1
XFILLER_0_181_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20767_ _05852_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22506_ _07070_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__buf_4
X_29062_ clknet_leaf_218_clock _02075_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23486_ decode.control.io_funct7\[3\] _07876_ _07873_ VGND VGND VPWR VPWR _07882_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26274_ net2524 _09462_ _09467_ _09458_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20698_ _00514_ _05656_ _05816_ net182 net2707 VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28013_ clknet_leaf_188_clock _01035_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_25225_ _08064_ net1406 _08837_ VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__mux2_1
X_22437_ _07029_ _06690_ _06672_ _07031_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__a211o_1
XFILLER_0_162_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22368_ _06959_ _06962_ _06640_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__mux2_4
X_25156_ _10556_ _10557_ _06281_ _10568_ VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__or4b_2
XFILLER_0_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24107_ _08226_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__clkbuf_1
X_21319_ net1409 _10803_ _06168_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25087_ _08771_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22299_ _06642_ _06742_ _06746_ _06752_ net88 VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__o311a_1
XFILLER_0_131_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28915_ clknet_leaf_140_clock _01928_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_24038_ net1518 execute.io_target_pc\[7\] _08187_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold390 decode.regfile.registers_29\[2\] VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__dlygate4sd3_1
X_29895_ clknet_leaf_301_clock _02908_ VGND VGND VPWR VPWR decode.regfile.registers_20\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_28846_ clknet_leaf_86_clock _01859_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_16860_ _12681_ VGND VGND VPWR VPWR _12822_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_196_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15811_ _11761_ net427 _11762_ _11795_ _11760_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_221_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28777_ clknet_leaf_96_clock _01790_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16791_ _10599_ _10924_ _12500_ _10935_ VGND VGND VPWR VPWR _12755_ sky130_fd_sc_hd__or4_2
X_25989_ net2261 _09286_ _09290_ _09277_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__o211a_1
X_18530_ _03828_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__buf_2
X_27728_ clknet_leaf_65_clock _00757_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_15742_ decode.regfile.registers_11\[11\] _11071_ _11470_ _11278_ VGND VGND VPWR
+ VPWR _11728_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1090 fetch.bht.bhtTable_tag\[11\]\[25\] VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18461_ _03673_ _03732_ _03733_ _03742_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__and4_1
XFILLER_0_217_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15673_ _11651_ _11659_ _11660_ VGND VGND VPWR VPWR _11661_ sky130_fd_sc_hd__o21a_1
X_27659_ clknet_leaf_26_clock _00688_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_293_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_293_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17412_ decode.regfile.registers_19\[15\] _10599_ _10589_ _12518_ _12543_ VGND VGND
+ VPWR VPWR _13362_ sky130_fd_sc_hd__o41a_1
XFILLER_0_68_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _10666_ VGND VGND VPWR VPWR _10667_ sky130_fd_sc_hd__clkbuf_4
X_18392_ decode.io_wb_rd\[4\] decode.id_ex_ex_rs1_reg\[4\] VGND VGND VPWR VPWR _03691_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_213_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29329_ clknet_leaf_226_clock _02342_ VGND VGND VPWR VPWR decode.regfile.registers_2\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17343_ _12915_ decode.regfile.registers_25\[13\] _13045_ _13294_ VGND VGND VPWR
+ VPWR _13295_ sky130_fd_sc_hd__or4_1
XFILLER_0_138_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14555_ _10597_ VGND VGND VPWR VPWR _10598_ sky130_fd_sc_hd__buf_4
XFILLER_0_172_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13506_ _09881_ _09884_ _09885_ _09887_ net393 VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__a41o_1
X_17274_ _12530_ _12616_ _12557_ decode.regfile.registers_0\[12\] VGND VGND VPWR VPWR
+ _13227_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14486_ _10107_ _10530_ VGND VGND VPWR VPWR _10539_ sky130_fd_sc_hd__nand2_1
X_19013_ _03635_ _03634_ net257 _04311_ _04299_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__o32a_1
XFILLER_0_181_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16225_ _11250_ _11258_ decode.regfile.registers_27\[23\] _12170_ _12198_ VGND VGND
+ VPWR VPWR _12199_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_114_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer2 net228 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_1
XFILLER_0_141_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16156_ _11248_ VGND VGND VPWR VPWR _12132_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_185_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_231_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_231_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_110_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15107_ _10650_ _10632_ VGND VGND VPWR VPWR _11104_ sky130_fd_sc_hd__nand2_2
XFILLER_0_107_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16087_ _11045_ _11410_ _12063_ VGND VGND VPWR VPWR _12064_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_224_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19915_ _04443_ _04242_ _04817_ _04879_ _05182_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15038_ _10659_ _10654_ VGND VGND VPWR VPWR _11035_ sky130_fd_sc_hd__and2_2
XFILLER_0_220_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19846_ _04325_ _05070_ _04317_ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_88_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_246_clock clknet_5_19__leaf_clock VGND VGND VPWR VPWR clknet_leaf_246_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_208_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16989_ decode.regfile.registers_16\[5\] _12575_ _12926_ _12948_ VGND VGND VPWR VPWR
+ _12949_ sky130_fd_sc_hd__o22a_1
X_19777_ _03852_ _03839_ _03851_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_218_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18728_ _09974_ _03771_ _03969_ _03970_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_140_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18659_ _03903_ _03939_ _03948_ _03957_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_78_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21670_ csr._mcycle_T_2\[20\] _06329_ _06378_ csr.minstret\[20\] VGND VGND VPWR VPWR
+ _06379_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_4_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20621_ csr.minstret\[25\] _05574_ _05586_ csr.mcycle\[25\] _05755_ VGND VGND VPWR
+ VPWR _05756_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23340_ _07765_ _07766_ _07081_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20552_ csr.mcycle\[15\] _05588_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_138_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23271_ _07064_ _07689_ _07690_ _07702_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20483_ _05534_ csr.minstret\[7\] _05538_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22222_ fetch.bht.bhtTable_tag\[0\]\[20\] fetch.bht.bhtTable_tag\[1\]\[20\] fetch.bht.bhtTable_tag\[2\]\[20\]
+ fetch.bht.bhtTable_tag\[3\]\[20\] net303 _06620_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__mux4_1
XFILLER_0_162_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25010_ _06331_ _08635_ _08720_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__nor3_1
XFILLER_0_6_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22153_ fetch.bht.bhtTable_tag\[12\]\[23\] fetch.bht.bhtTable_tag\[13\]\[23\] _06618_
+ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21104_ net100 net111 execute.io_mem_memwrite VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22084_ _06615_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__buf_6
X_26961_ _10073_ _09862_ VGND VGND VPWR VPWR _09863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28700_ clknet_leaf_175_clock _01713_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25912_ _08910_ _09243_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__nand2_1
X_21035_ execute.csr_read_data_out_reg\[7\] _06002_ _05998_ VGND VGND VPWR VPWR _06003_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_227_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29680_ clknet_leaf_283_clock _02693_ VGND VGND VPWR VPWR decode.regfile.registers_13\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_26892_ net1755 _09822_ _09823_ _09812_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28631_ clknet_leaf_117_clock _01644_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_25843_ _08916_ _09200_ VGND VGND VPWR VPWR _09206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28562_ clknet_leaf_202_clock _01575_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25774_ _09155_ VGND VGND VPWR VPWR _09166_ sky130_fd_sc_hd__clkbuf_4
X_22986_ fetch.bht.bhtTable_target_pc\[0\]\[6\] fetch.bht.bhtTable_target_pc\[1\]\[6\]
+ fetch.bht.bhtTable_target_pc\[2\]\[6\] fetch.bht.bhtTable_target_pc\[3\]\[6\] _07407_
+ _07115_ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__mux4_1
X_27513_ clknet_leaf_15_clock _00542_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dfxtp_1
X_24725_ _08087_ net1720 _08542_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28493_ clknet_leaf_197_clock _01506_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21937_ _03449_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__buf_4
XFILLER_0_167_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27444_ clknet_leaf_151_clock _00473_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_24656_ _08511_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__clkbuf_1
X_21868_ _06516_ _06494_ _06495_ _06517_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23607_ _07949_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27375_ clknet_leaf_9_clock _00404_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_20819_ net128 _05879_ _05875_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__and3_1
X_24587_ net828 execute.io_target_pc\[15\] _08473_ VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21799_ csr._mcycle_T_2\[7\] _06467_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__or2b_1
XFILLER_0_166_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_189_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29114_ clknet_leaf_70_clock _02127_ VGND VGND VPWR VPWR csr._mcycle_T_3\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26326_ net758 _09491_ _09497_ _09484_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__o211a_1
X_14340_ _10117_ _10444_ VGND VGND VPWR VPWR _10455_ sky130_fd_sc_hd__nand2_1
X_23538_ net2152 _07904_ _07901_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__or3b_1
XFILLER_0_167_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_189_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29045_ clknet_leaf_115_clock _02058_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26257_ _09417_ VGND VGND VPWR VPWR _09458_ sky130_fd_sc_hd__clkbuf_4
X_14271_ net1151 _10403_ _10414_ _10411_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23469_ net14 _07861_ _07871_ _07865_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__o211a_2
XFILLER_0_107_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16010_ decode.regfile.registers_5\[18\] _11192_ _11139_ VGND VGND VPWR VPWR _11989_
+ sky130_fd_sc_hd__and3_1
X_25208_ _10572_ net2750 _08832_ VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26188_ _09410_ _09390_ VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_227_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25139_ _03528_ _07250_ _08798_ _10998_ _03458_ VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_148_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17961_ decode.regfile.registers_16\[29\] _13011_ _12579_ _03358_ VGND VGND VPWR
+ VPWR _03359_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_223_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19700_ _04937_ _04193_ _03963_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__a21oi_1
X_16912_ _10931_ decode.regfile.registers_30\[4\] _12487_ VGND VGND VPWR VPWR _12873_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_218_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17892_ _12712_ decode.regfile.registers_24\[27\] _12997_ _12998_ _11025_ VGND VGND
+ VPWR VPWR _03292_ sky130_fd_sc_hd__o2111a_1
X_29878_ clknet_leaf_300_clock _02891_ VGND VGND VPWR VPWR decode.regfile.registers_19\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16843_ _12755_ VGND VGND VPWR VPWR _12806_ sky130_fd_sc_hd__clkbuf_4
X_19631_ _04204_ _04206_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__and2_1
X_28829_ clknet_leaf_179_clock _01842_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19562_ _04408_ _04209_ _04620_ _03933_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__or4_1
X_16774_ decode.regfile.registers_7\[1\] _12610_ _12737_ decode.regfile.registers_6\[1\]
+ VGND VGND VPWR VPWR _12738_ sky130_fd_sc_hd__a22oi_1
X_13986_ _09984_ _10244_ VGND VGND VPWR VPWR _10251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18513_ net196 _03772_ _03775_ _03806_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__a211oi_4
XTAP_TAPCELL_ROW_17_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15725_ decode.regfile.registers_19\[10\] _11453_ _11688_ _11711_ _11454_ VGND VGND
+ VPWR VPWR _11712_ sky130_fd_sc_hd__o221a_1
X_19493_ net66 _10908_ _10758_ _03636_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__or4b_4
XFILLER_0_125_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18444_ _09934_ csr.io_csr_address\[3\] _03740_ _03742_ VGND VGND VPWR VPWR _03743_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15656_ _11344_ net435 _11610_ _11644_ _11249_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__o221a_1
XFILLER_0_185_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_199_Right_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14607_ _10649_ VGND VGND VPWR VPWR _10650_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18375_ decode.io_wb_rd\[4\] _03652_ decode.id_ex_ex_rs1_reg\[1\] _09931_ VGND VGND
+ VPWR VPWR _03674_ sky130_fd_sc_hd__o22a_1
X_15587_ decode.regfile.registers_3\[7\] _11157_ _11140_ _11145_ VGND VGND VPWR VPWR
+ _11577_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17326_ _13266_ _13277_ _12591_ VGND VGND VPWR VPWR _13278_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14538_ decode.control.io_opcode\[6\] decode.control.io_opcode\[5\] decode.control.io_opcode\[4\]
+ _10580_ VGND VGND VPWR VPWR _10581_ sky130_fd_sc_hd__and4_1
XFILLER_0_83_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_1160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17257_ _12915_ decode.regfile.registers_25\[11\] _13045_ _12812_ VGND VGND VPWR
+ VPWR _13211_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14469_ _10069_ _10517_ VGND VGND VPWR VPWR _10529_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_77_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_170_clock clknet_5_24__leaf_clock VGND VGND VPWR VPWR clknet_leaf_170_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16208_ decode.regfile.registers_7\[23\] _11092_ _11167_ _11134_ VGND VGND VPWR VPWR
+ _12182_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_133_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17188_ _12934_ _10592_ _12558_ decode.regfile.registers_0\[10\] VGND VGND VPWR VPWR
+ _13143_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16139_ _11046_ decode.regfile.registers_12\[21\] _10650_ _11052_ _10632_ VGND VGND
+ VPWR VPWR _12115_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_122_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_185_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_185_clock
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_102_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2505 csr._minstret_T_3\[50\] VGND VGND VPWR VPWR net2732 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2516 execute.io_wfi_out VGND VGND VPWR VPWR net2743 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2527 csr._mcycle_T_2\[20\] VGND VGND VPWR VPWR net2754 sky130_fd_sc_hd__buf_1
Xhold2538 csr._csr_read_data_T_8\[11\] VGND VGND VPWR VPWR net2765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1804 fetch.bht.bhtTable_target_pc\[7\]\[26\] VGND VGND VPWR VPWR net2031 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2549 decode.regfile.registers_30\[15\] VGND VGND VPWR VPWR net2776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1815 csr.mscratch\[3\] VGND VGND VPWR VPWR net2042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1826 fetch.bht.bhtTable_tag\[7\]\[24\] VGND VGND VPWR VPWR net2053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19829_ _05076_ _05052_ _05100_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__o21bai_2
Xhold1837 fetch.bht.bhtTable_target_pc\[14\]\[18\] VGND VGND VPWR VPWR net2064 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1848 fetch.bht.bhtTable_target_pc\[9\]\[10\] VGND VGND VPWR VPWR net2075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 fetch.bht.bhtTable_tag\[5\]\[19\] VGND VGND VPWR VPWR net2086 sky130_fd_sc_hd__dlygate4sd3_1
X_22840_ net1435 _10821_ _09898_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22771_ _06145_ net1176 _07276_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24510_ _08070_ net1613 _08428_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21722_ csr.minstret\[29\] csr.minstret\[30\] _06415_ VGND VGND VPWR VPWR _06420_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_56_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25490_ _08941_ _08992_ VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_123_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_123_clock
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_111_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24441_ _08399_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__clkbuf_1
X_21653_ csr._mcycle_T_2\[15\] _06329_ _06366_ _05691_ VGND VGND VPWR VPWR _06367_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20604_ csr.mscratch\[23\] _03718_ _05554_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__or3_1
X_27160_ clknet_leaf_356_clock _00189_ VGND VGND VPWR VPWR decode.regfile.registers_27\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24372_ net1187 execute.io_target_pc\[9\] _08356_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__mux2_1
X_21584_ csr.io_csr_write_address\[5\] csr.io_csr_write_address\[4\] csr.io_csr_write_address\[7\]
+ csr.io_csr_write_address\[6\] VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__nor4_2
XFILLER_0_47_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26111_ net2703 _09356_ _09360_ _09359_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__o211a_1
X_23323_ _07749_ _07750_ _07081_ VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__mux2_1
X_20535_ _05541_ csr.io_mret_vector\[13\] _05602_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27091_ clknet_leaf_328_clock _00120_ VGND VGND VPWR VPWR decode.regfile.registers_25\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_138_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_138_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26042_ decode.regfile.registers_9\[25\] _09313_ _09320_ _09318_ VGND VGND VPWR VPWR
+ _02568_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23254_ _07619_ _07573_ _07620_ _07686_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__a31o_1
X_20466_ _05621_ _05219_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22205_ _06652_ _06797_ _06632_ _06799_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23185_ _07417_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__buf_2
X_20397_ csr.mscratch\[0\] _03718_ _05554_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__or3_1
XFILLER_0_127_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22136_ _06729_ _06730_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__nand2_1
X_29801_ clknet_leaf_297_clock _02814_ VGND VGND VPWR VPWR decode.regfile.registers_17\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_27993_ clknet_leaf_235_clock _01015_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22067_ fetch.bht.bhtTable_tag\[4\]\[18\] fetch.bht.bhtTable_tag\[5\]\[18\] _06646_
+ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__mux2_1
X_29732_ clknet_leaf_286_clock _02745_ VGND VGND VPWR VPWR decode.regfile.registers_15\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_26944_ _10030_ _09849_ VGND VGND VPWR VPWR _09854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21018_ _05993_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__clkbuf_1
X_29663_ clknet_leaf_271_clock _02676_ VGND VGND VPWR VPWR decode.regfile.registers_13\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_26875_ _09402_ _09806_ VGND VGND VPWR VPWR _09814_ sky130_fd_sc_hd__nand2_1
X_28614_ clknet_leaf_96_clock _01627_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13840_ _10015_ _10164_ VGND VGND VPWR VPWR _10165_ sky130_fd_sc_hd__nand2_1
X_25826_ net2239 _09157_ _09195_ _09194_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29594_ clknet_leaf_289_clock _02607_ VGND VGND VPWR VPWR decode.regfile.registers_11\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28545_ clknet_leaf_195_clock _01558_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13771_ memory.csr_read_data_out_reg\[25\] _09989_ _10110_ VGND VGND VPWR VPWR _10111_
+ sky130_fd_sc_hd__o21ai_2
X_25757_ _09155_ VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__buf_2
X_22969_ _06461_ _06041_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__nand2_2
XFILLER_0_58_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15510_ _11500_ _11501_ VGND VGND VPWR VPWR _11502_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24708_ _08070_ net1903 _08531_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28476_ clknet_leaf_222_clock _01489_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16490_ decode.regfile.registers_1\[31\] _11539_ VGND VGND VPWR VPWR _12456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25688_ _08912_ _09112_ VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15441_ _10957_ VGND VGND VPWR VPWR _11435_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27427_ clknet_leaf_40_clock _00456_ VGND VGND VPWR VPWR decode.id_ex_memtoreg_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_24639_ _08502_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_216_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_216_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18160_ _03508_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15372_ _11293_ VGND VGND VPWR VPWR _11367_ sky130_fd_sc_hd__buf_4
X_27358_ clknet_leaf_41_clock _00387_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[31\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17111_ _12499_ _12541_ _12490_ decode.regfile.registers_11\[8\] _12878_ VGND VGND
+ VPWR VPWR _13068_ sky130_fd_sc_hd__o32a_1
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14323_ net1059 _10434_ _10445_ _10440_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__o211a_1
X_26309_ _09441_ _09446_ VGND VGND VPWR VPWR _09487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18091_ _03471_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27289_ clknet_leaf_8_clock _00318_ VGND VGND VPWR VPWR decode.regfile.registers_31\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29028_ clknet_leaf_128_clock _02041_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_17042_ _10938_ decode.regfile.registers_25\[6\] _12505_ _12811_ VGND VGND VPWR VPWR
+ _13001_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14254_ net2493 _10403_ _10405_ _10398_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14185_ _10112_ _10355_ VGND VGND VPWR VPWR _10365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18993_ _04273_ _04278_ _04288_ _04291_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__a211o_1
XFILLER_0_209_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17944_ _12631_ decode.regfile.registers_0\[29\] VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__nand2_1
X_17875_ _03269_ _03273_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_105_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19614_ _04894_ _04414_ _04508_ _04242_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__and4b_1
X_16826_ _12654_ _12788_ VGND VGND VPWR VPWR _12789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_1332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16757_ _11017_ _10606_ _10935_ VGND VGND VPWR VPWR _12721_ sky130_fd_sc_hd__or3_1
X_19545_ _04827_ _04106_ _04104_ _04756_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__and4b_1
XFILLER_0_159_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13969_ _10147_ _10198_ VGND VGND VPWR VPWR _10239_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_40_clock clknet_5_6__leaf_clock VGND VGND VPWR VPWR clknet_leaf_40_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15708_ decode.regfile.registers_1\[10\] _11117_ _11057_ _11157_ VGND VGND VPWR VPWR
+ _11695_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_66_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16688_ _12652_ VGND VGND VPWR VPWR _12653_ sky130_fd_sc_hd__clkbuf_4
X_19476_ _04119_ net271 _04742_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__or3_1
XINSDIODE1_320 execute.io_target_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_0_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_0_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_331 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_342 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15639_ _11048_ decode.regfile.registers_12\[8\] _10651_ _11054_ _10633_ VGND VGND
+ VPWR VPWR _11628_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18427_ decode.id_ex_immsrc_reg VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_29_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_353 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_364 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_375 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_386 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_55_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_55_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_135_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18358_ execute.io_mem_memtoreg\[1\] execute.io_mem_memtoreg\[0\] VGND VGND VPWR
+ VPWR _03657_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_135_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17309_ _13055_ net430 _13097_ VGND VGND VPWR VPWR _13261_ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18289_ _03609_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20320_ _05490_ _05491_ _05420_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold901 fetch.bht.bhtTable_tag\[8\]\[15\] VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold912 fetch.bht.bhtTable_target_pc\[1\]\[6\] VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 fetch.bht.bhtTable_tag\[6\]\[15\] VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__dlygate4sd3_1
X_20251_ _05417_ _05274_ _05438_ _05414_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_9_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold934 fetch.bht.bhtTable_target_pc\[11\]\[5\] VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold945 decode.regfile.registers_21\[7\] VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold956 fetch.bht.bhtTable_tag\[4\]\[25\] VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 decode.regfile.registers_18\[7\] VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 fetch.bht.bhtTable_tag\[15\]\[14\] VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__dlygate4sd3_1
X_20182_ decode.id_ex_imm_reg\[25\] _10790_ _05381_ _05380_ VGND VGND VPWR VPWR _05383_
+ sky130_fd_sc_hd__o211ai_1
Xhold989 fetch.bht.bhtTable_tag\[1\]\[14\] VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2302 decode.regfile.registers_4\[27\] VGND VGND VPWR VPWR net2529 sky130_fd_sc_hd__dlygate4sd3_1
X_24990_ net569 _08701_ net1617 _06318_ _08706_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__a311oi_1
Xhold2313 decode.regfile.registers_6\[18\] VGND VGND VPWR VPWR net2540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2324 csr._csr_read_data_T_8\[16\] VGND VGND VPWR VPWR net2551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2335 decode.regfile.registers_10\[1\] VGND VGND VPWR VPWR net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1601 fetch.bht.bhtTable_target_pc\[6\]\[17\] VGND VGND VPWR VPWR net1828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2346 decode.regfile.registers_13\[23\] VGND VGND VPWR VPWR net2573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1612 fetch.bht.bhtTable_tag\[10\]\[22\] VGND VGND VPWR VPWR net1839 sky130_fd_sc_hd__dlygate4sd3_1
X_23941_ net907 _08099_ _06156_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__mux2_1
Xhold2357 fetch.btb.btbTable\[14\]\[1\] VGND VGND VPWR VPWR net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1623 decode.regfile.registers_3\[12\] VGND VGND VPWR VPWR net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2368 decode.regfile.registers_4\[28\] VGND VGND VPWR VPWR net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1634 fetch.bht.bhtTable_tag\[4\]\[17\] VGND VGND VPWR VPWR net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2379 decode.regfile.registers_6\[7\] VGND VGND VPWR VPWR net2606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1645 fetch.bht.bhtTable_tag\[14\]\[24\] VGND VGND VPWR VPWR net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1656 fetch.bht.bhtTable_tag\[3\]\[8\] VGND VGND VPWR VPWR net1883 sky130_fd_sc_hd__dlygate4sd3_1
X_26660_ _09412_ _09689_ VGND VGND VPWR VPWR _09690_ sky130_fd_sc_hd__nand2_1
Xhold1667 fetch.bht.bhtTable_tag\[5\]\[10\] VGND VGND VPWR VPWR net1894 sky130_fd_sc_hd__dlygate4sd3_1
X_23872_ _08102_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__clkbuf_1
Xhold1678 fetch.bht.bhtTable_tag\[14\]\[15\] VGND VGND VPWR VPWR net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1689 fetch.bht.bhtTable_tag\[14\]\[19\] VGND VGND VPWR VPWR net1916 sky130_fd_sc_hd__dlygate4sd3_1
X_25611_ net1394 _09068_ _09072_ _09059_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__o211a_1
X_22823_ net1299 _10773_ _07297_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__mux2_1
X_26591_ net1669 _09649_ _09650_ _09648_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_212_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28330_ clknet_leaf_184_clock _01343_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25542_ _08990_ VGND VGND VPWR VPWR _09033_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22754_ _06128_ net1046 _07265_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_891 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21705_ net584 _06404_ _06406_ _06352_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__a211oi_1
X_28261_ clknet_leaf_78_clock _01283_ VGND VGND VPWR VPWR csr._minstret_T_3\[61\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25473_ _08922_ _08992_ VGND VGND VPWR VPWR _08993_ sky130_fd_sc_hd__nand2_1
X_22685_ csr._mcycle_T_2\[18\] _07223_ VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__or2_1
XFILLER_0_212_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27212_ clknet_leaf_364_clock _00241_ VGND VGND VPWR VPWR decode.regfile.registers_28\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_24424_ _08051_ net869 _08389_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28192_ clknet_leaf_113_clock _01214_ VGND VGND VPWR VPWR csr.io_mret_vector\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_21636_ net606 net1443 _06350_ _06353_ _06336_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27143_ clknet_leaf_358_clock _00172_ VGND VGND VPWR VPWR decode.regfile.registers_26\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_24355_ net1492 execute.io_target_pc\[1\] _06141_ VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__mux2_1
X_21567_ _06138_ net2476 _06295_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23306_ fetch.bht.bhtTable_target_pc\[0\]\[24\] fetch.bht.bhtTable_target_pc\[1\]\[24\]
+ fetch.bht.bhtTable_target_pc\[2\]\[24\] fetch.bht.bhtTable_target_pc\[3\]\[24\]
+ _07555_ _07710_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20518_ csr.io_mret_vector\[11\] _05580_ _05581_ csr.mscratch\[11\] _05666_ VGND
+ VGND VPWR VPWR _05667_ sky130_fd_sc_hd__a221o_1
X_27074_ clknet_leaf_346_clock _00103_ VGND VGND VPWR VPWR decode.regfile.registers_24\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_24286_ _08318_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__clkbuf_1
X_21498_ _06266_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26025_ _08945_ _09310_ VGND VGND VPWR VPWR _09311_ sky130_fd_sc_hd__nand2_1
X_23237_ _07666_ _07668_ _07670_ _07075_ _06740_ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__a221o_1
Xclkbuf_5_9__f_clock clknet_2_1_0_clock VGND VGND VPWR VPWR clknet_5_9__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_20449_ _05592_ csr.io_mret_vector\[3\] _05603_ _05605_ VGND VGND VPWR VPWR _05606_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23168_ fetch.bht.bhtTable_target_pc\[12\]\[16\] fetch.bht.bhtTable_target_pc\[13\]\[16\]
+ fetch.bht.bhtTable_target_pc\[14\]\[16\] fetch.bht.bhtTable_target_pc\[15\]\[16\]
+ _07439_ _07112_ VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22119_ fetch.bht.bhtTable_tag\[14\]\[3\] fetch.bht.bhtTable_tag\[15\]\[3\] _06674_
+ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__mux2_1
X_23099_ fetch.bht.bhtTable_target_pc\[0\]\[12\] fetch.bht.bhtTable_target_pc\[1\]\[12\]
+ fetch.bht.bhtTable_target_pc\[2\]\[12\] fetch.bht.bhtTable_target_pc\[3\]\[12\]
+ _07107_ _07071_ VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__mux4_1
X_27976_ clknet_leaf_208_clock _00998_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_15990_ decode.regfile.registers_18\[17\] _10955_ _11114_ _11094_ _10976_ VGND VGND
+ VPWR VPWR _11970_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_219_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14941_ csr.io_mret VGND VGND VPWR VPWR _10970_ sky130_fd_sc_hd__clkbuf_4
X_29715_ clknet_leaf_284_clock _02728_ VGND VGND VPWR VPWR decode.regfile.registers_14\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_26927_ net210 _09840_ VGND VGND VPWR VPWR _09844_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_202_Right_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17660_ _02986_ decode.regfile.registers_26\[21\] _13254_ _13484_ _02987_ VGND VGND
+ VPWR VPWR _03066_ sky130_fd_sc_hd__o2111a_1
X_14872_ _10670_ decode.id_ex_memread_reg VGND VGND VPWR VPWR _10914_ sky130_fd_sc_hd__or2b_1
X_29646_ clknet_leaf_279_clock _02659_ VGND VGND VPWR VPWR decode.regfile.registers_12\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_26858_ _09385_ _09796_ VGND VGND VPWR VPWR _09804_ sky130_fd_sc_hd__nand2_1
X_16611_ _12575_ VGND VGND VPWR VPWR _12576_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_215_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13823_ net809 _10153_ _10155_ _10132_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__o211a_1
X_25809_ net2344 _09183_ _09186_ _09182_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17591_ decode.regfile.registers_18\[20\] _10924_ _12568_ _12524_ _10612_ VGND VGND
+ VPWR VPWR _02998_ sky130_fd_sc_hd__o2111a_1
X_29577_ clknet_leaf_273_clock _02590_ VGND VGND VPWR VPWR decode.regfile.registers_10\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_207_Left_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26789_ net1002 _09752_ _09764_ _09758_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_218_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28528_ clknet_leaf_218_clock _01541_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16542_ _12506_ VGND VGND VPWR VPWR _12507_ sky130_fd_sc_hd__buf_2
X_19330_ _04408_ _04620_ _04621_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__or3_1
XFILLER_0_134_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13754_ _10096_ VGND VGND VPWR VPWR _10097_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19261_ _04280_ _04282_ _04554_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__or3_1
XFILLER_0_169_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28459_ clknet_leaf_149_clock _01472_ VGND VGND VPWR VPWR decode.io_id_pc\[17\] sky130_fd_sc_hd__dfxtp_1
X_16473_ decode.regfile.registers_20\[30\] _11103_ _11327_ _12439_ VGND VGND VPWR
+ VPWR _12440_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13685_ _09939_ memory.io_wb_aluresult\[12\] _09940_ VGND VGND VPWR VPWR _10038_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_195_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18212_ _11347_ _03529_ _11011_ _12636_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__or4b_1
X_15424_ decode.regfile.registers_8\[3\] _11285_ _11365_ decode.regfile.registers_9\[3\]
+ _11132_ VGND VGND VPWR VPWR _11418_ sky130_fd_sc_hd__o221a_1
XFILLER_0_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19192_ _04045_ _04320_ _04487_ _04332_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_122_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18143_ _03495_ _03493_ _03500_ net2103 VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_143_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15355_ _11079_ _10979_ _10958_ _11080_ VGND VGND VPWR VPWR _11350_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14306_ _10036_ _10431_ VGND VGND VPWR VPWR _10436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18074_ _03460_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15286_ decode.regfile.registers_9\[1\] _11280_ _11281_ _11183_ VGND VGND VPWR VPWR
+ _11282_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_216_Left_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire172 _01316_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold208 decode.regfile.registers_31\[8\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkdlybuf4s25_1
Xwire183 _05815_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_151_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17025_ _12669_ VGND VGND VPWR VPWR _12984_ sky130_fd_sc_hd__clkbuf_4
Xhold219 decode.regfile.registers_30\[8\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14237_ net1622 _10390_ _10395_ _10385_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14168_ _10331_ VGND VGND VPWR VPWR _10355_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18976_ net188 _03812_ _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__mux2_1
X_14099_ _10087_ _10312_ VGND VGND VPWR VPWR _10316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ decode.regfile.registers_19\[28\] _12679_ _12545_ _03325_ VGND VGND VPWR
+ VPWR _03326_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17858_ _02990_ _03068_ decode.regfile.registers_27\[26\] _13487_ VGND VGND VPWR
+ VPWR _03259_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_225_Left_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16809_ _12722_ VGND VGND VPWR VPWR _12772_ sky130_fd_sc_hd__clkbuf_4
X_17789_ decode.regfile.registers_1\[25\] _12636_ _13145_ _12835_ VGND VGND VPWR VPWR
+ _03191_ sky130_fd_sc_hd__a31o_1
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19528_ _04180_ _04181_ _03989_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19459_ net265 _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__xor2_1
XFILLER_0_147_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_150 _12597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_161 _13433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_172 decode.id_ex_rs1_data_reg\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_183 execute.io_target_pc\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22470_ _10758_ _10914_ _07064_ _03590_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_194 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1096 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21421_ _06225_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24140_ _08243_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__clkbuf_1
X_21352_ _06187_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20303_ _05478_ _05219_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24071_ net1190 execute.io_target_pc\[23\] _08198_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__mux2_1
X_21283_ _06148_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__clkbuf_1
Xhold720 fetch.bht.bhtTable_tag\[11\]\[9\] VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold731 fetch.bht.bhtTable_tag\[3\]\[18\] VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold742 decode.regfile.registers_12\[30\] VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold753 fetch.bht.bhtTable_tag\[1\]\[7\] VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__dlygate4sd3_1
X_23022_ csr._csr_read_data_T_8\[7\] _06038_ csr.io_mret_vector\[7\] _06462_ VGND
+ VGND VPWR VPWR _07468_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_57_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20234_ _03581_ _05424_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__and3b_1
Xhold764 fetch.bht.bhtTable_target_pc\[14\]\[9\] VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold775 decode.regfile.registers_19\[8\] VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold786 fetch.bht.bhtTable_target_pc\[12\]\[16\] VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 fetch.bht.bhtTable_target_pc\[1\]\[8\] VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__dlygate4sd3_1
X_27830_ clknet_leaf_321_clock _00859_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20165_ decode.id_ex_imm_reg\[24\] decode.id_ex_pc_reg\[24\] VGND VGND VPWR VPWR
+ _05368_ sky130_fd_sc_hd__nor2_1
Xhold2110 decode.regfile.registers_6\[27\] VGND VGND VPWR VPWR net2337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2121 execute.csr_write_data_out_reg\[10\] VGND VGND VPWR VPWR net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2132 decode.regfile.registers_5\[28\] VGND VGND VPWR VPWR net2359 sky130_fd_sc_hd__dlygate4sd3_1
X_27761_ clknet_leaf_318_clock _00790_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_20096_ decode.id_ex_imm_reg\[14\] decode.id_ex_pc_reg\[14\] VGND VGND VPWR VPWR
+ _05309_ sky130_fd_sc_hd__nand2_1
Xhold2143 decode.regfile.registers_1\[12\] VGND VGND VPWR VPWR net2370 sky130_fd_sc_hd__dlygate4sd3_1
X_24973_ net2365 _08693_ net699 VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__a21oi_1
Xhold2154 decode.regfile.registers_4\[21\] VGND VGND VPWR VPWR net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1420 fetch.bht.bhtTable_target_pc\[13\]\[4\] VGND VGND VPWR VPWR net1647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2165 decode.regfile.registers_24\[21\] VGND VGND VPWR VPWR net2392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1431 fetch.bht.bhtTable_target_pc\[7\]\[16\] VGND VGND VPWR VPWR net1658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2176 decode.regfile.registers_24\[29\] VGND VGND VPWR VPWR net2403 sky130_fd_sc_hd__dlygate4sd3_1
X_26712_ _09708_ VGND VGND VPWR VPWR _09720_ sky130_fd_sc_hd__clkbuf_4
X_29500_ clknet_leaf_251_clock _02513_ VGND VGND VPWR VPWR decode.regfile.registers_8\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23924_ _08132_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__clkbuf_1
Xhold1442 decode.regfile.registers_16\[20\] VGND VGND VPWR VPWR net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2187 decode.regfile.registers_23\[19\] VGND VGND VPWR VPWR net2414 sky130_fd_sc_hd__dlygate4sd3_1
X_27692_ clknet_leaf_26_clock _00721_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1453 fetch.bht.bhtTable_tag\[9\]\[4\] VGND VGND VPWR VPWR net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2198 execute.exception_out_reg VGND VGND VPWR VPWR net2425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 execute.csr_write_data_out_reg\[16\] VGND VGND VPWR VPWR net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 fetch.bht.bhtTable_target_pc\[11\]\[20\] VGND VGND VPWR VPWR net1702 sky130_fd_sc_hd__dlygate4sd3_1
X_29431_ clknet_leaf_261_clock _02444_ VGND VGND VPWR VPWR decode.regfile.registers_5\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1486 fetch.bht.bhtTable_target_pc\[5\]\[21\] VGND VGND VPWR VPWR net1713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26643_ net653 _09679_ _09680_ _09675_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23855_ execute.io_target_pc\[20\] VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__clkbuf_2
Xhold1497 decode.regfile.registers_17\[16\] VGND VGND VPWR VPWR net1724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22806_ _07298_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__clkbuf_1
X_29362_ clknet_leaf_227_clock _02375_ VGND VGND VPWR VPWR decode.regfile.registers_3\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_26574_ net1924 _09636_ _09640_ _09635_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23786_ _08045_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ _05982_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__clkbuf_1
X_28313_ clknet_leaf_208_clock _01326_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25525_ net2185 _08980_ _09021_ _09017_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22737_ _06111_ net2177 _09903_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__mux2_1
X_29293_ clknet_leaf_231_clock _02306_ VGND VGND VPWR VPWR decode.regfile.registers_1\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_213_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28244_ clknet_leaf_77_clock _01266_ VGND VGND VPWR VPWR csr._minstret_T_3\[44\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25456_ _08982_ _08980_ VGND VGND VPWR VPWR _08983_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22668_ csr._mcycle_T_2\[11\] _07210_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24407_ net988 execute.io_target_pc\[26\] _09911_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28175_ clknet_leaf_57_clock _01197_ VGND VGND VPWR VPWR csr.io_mret_vector\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_21619_ csr.minstret\[6\] _06340_ _06341_ _06331_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__a211oi_1
X_25387_ net2370 _08928_ _08934_ _08927_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22599_ csr._minstret_T_3\[47\] _07174_ net1978 VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15140_ _11055_ VGND VGND VPWR VPWR _11137_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_11_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27126_ clknet_leaf_351_clock _00155_ VGND VGND VPWR VPWR decode.regfile.registers_26\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24338_ _08345_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15071_ _10961_ decode.regfile.registers_28\[0\] _11067_ _11038_ _10994_ VGND VGND
+ VPWR VPWR _11068_ sky130_fd_sc_hd__o2111a_1
X_27057_ clknet_leaf_330_clock _00086_ VGND VGND VPWR VPWR decode.regfile.registers_24\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_24269_ _08097_ net1546 _08300_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__mux2_1
X_14022_ _10242_ VGND VGND VPWR VPWR _10271_ sky130_fd_sc_hd__clkbuf_4
X_26008_ net551 _09300_ _09301_ _09292_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_207_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18830_ _03890_ decode.id_ex_imm_reg\[8\] _04127_ _04128_ VGND VGND VPWR VPWR _04129_
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_101_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15973_ decode.regfile.registers_3\[17\] _11109_ _11140_ _11145_ VGND VGND VPWR VPWR
+ _11953_ sky130_fd_sc_hd__a31o_1
X_18761_ memory.csr_read_data_out_reg\[7\] _09986_ _10002_ _10006_ VGND VGND VPWR
+ VPWR _04060_ sky130_fd_sc_hd__o22a_1
X_27959_ clknet_leaf_189_clock _00981_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14924_ _10949_ _10950_ _10952_ VGND VGND VPWR VPWR _10953_ sky130_fd_sc_hd__or3_1
XFILLER_0_117_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17712_ decode.regfile.registers_10\[23\] _12790_ _12878_ VGND VGND VPWR VPWR _03116_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18692_ net207 net206 _09963_ net203 VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_188_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_215_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14855_ decode.id_ex_pc_reg\[12\] _10880_ _10883_ _10897_ VGND VGND VPWR VPWR _10898_
+ sky130_fd_sc_hd__o211ai_1
X_17643_ _03047_ _03048_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__nand2_1
X_29629_ clknet_leaf_288_clock _02642_ VGND VGND VPWR VPWR decode.regfile.registers_12\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13806_ memory.csr_read_data_out_reg\[30\] _09989_ _10140_ VGND VGND VPWR VPWR _10141_
+ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_63_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17574_ _13081_ _13168_ decode.regfile.registers_23\[19\] _13041_ VGND VGND VPWR
+ VPWR _02982_ sky130_fd_sc_hd__or4_1
X_14786_ _09928_ _10828_ VGND VGND VPWR VPWR _10829_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19313_ _04588_ _04596_ _04605_ _04459_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__o31a_2
X_16525_ _12489_ VGND VGND VPWR VPWR _12490_ sky130_fd_sc_hd__clkbuf_4
X_13737_ net1946 _10027_ _10082_ _10077_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_158_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16456_ decode.regfile.registers_1\[30\] _11115_ _11056_ _11108_ VGND VGND VPWR VPWR
+ _12423_ sky130_fd_sc_hd__and4_1
XFILLER_0_129_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19244_ _03635_ _03634_ _03637_ _03633_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__and4b_2
XFILLER_0_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13668_ memory.csr_read_data_out_reg\[9\] _09988_ _10022_ _10023_ VGND VGND VPWR
+ VPWR _10024_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_144_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15407_ _11344_ net801 _11345_ _11401_ _11249_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__o221a_1
XFILLER_0_183_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19175_ _04269_ _04468_ _04470_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16387_ _11042_ decode.regfile.registers_4\[28\] _11190_ _10628_ _11083_ VGND VGND
+ VPWR VPWR _12356_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_22_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13599_ memory.csr_read_data_out_reg\[1\] _09941_ _09959_ _09962_ VGND VGND VPWR
+ VPWR _09963_ sky130_fd_sc_hd__o22ai_4
X_18126_ _03482_ _03480_ _03487_ decode.io_id_pc\[19\] VGND VGND VPWR VPWR _03491_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_147_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15338_ _11059_ _10977_ _10955_ _11072_ VGND VGND VPWR VPWR _11334_ sky130_fd_sc_hd__or4b_1
XFILLER_0_147_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18057_ _10965_ _10972_ _10969_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__and4bb_1
X_15269_ _10989_ VGND VGND VPWR VPWR _11265_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_188_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17008_ _12495_ VGND VGND VPWR VPWR _12967_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18959_ _04251_ _04252_ _04257_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__a21o_1
XFILLER_0_226_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21970_ _06571_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer12 net238 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_1
X_20921_ _05937_ _05933_ net46 VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__and3_1
Xrebuffer23 _03757_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__buf_1
XFILLER_0_55_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer34 _04229_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer45 _03784_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer56 _04105_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd1_1
X_23640_ net1039 csr.io_mem_pc\[12\] _07961_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__mux2_1
Xrebuffer67 net293 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_1
X_20852_ _05866_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__clkbuf_2
Xrebuffer78 _03752_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer89 net360 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23571_ _09914_ net338 _07930_ net521 VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20783_ _05864_ _09954_ net2670 VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25310_ _08885_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22522_ fetch.bht.bhtTable_target_pc\[0\]\[1\] fetch.bht.bhtTable_target_pc\[1\]\[1\]
+ _07099_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26290_ _09422_ _09472_ VGND VGND VPWR VPWR _09477_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25241_ _08850_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22453_ _06699_ _07039_ _07041_ _07047_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__a31o_1
XFILLER_0_146_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer102 net328 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer113 _08633_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__buf_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21404_ _06215_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25172_ _10573_ net2751 _08814_ VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22384_ fetch.bht.bhtTable_tag\[4\]\[9\] fetch.bht.bhtTable_tag\[5\]\[9\] _06878_
+ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_27__f_clock clknet_2_3_0_clock VGND VGND VPWR VPWR clknet_5_27__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_161_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24123_ net919 execute.io_target_pc\[16\] _08232_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21335_ net1941 _10773_ _06168_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24054_ _08199_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__clkbuf_1
X_28931_ clknet_leaf_130_clock _01944_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21266_ net1517 _06136_ _06120_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold550 csr._mcycle_T_2\[6\] VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__clkbuf_2
Xhold561 decode.id_ex_imm_reg\[0\] VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 fetch.bht.bhtTable_target_pc\[2\]\[19\] VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold583 fetch.bht.bhtTable_target_pc\[4\]\[27\] VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__dlygate4sd3_1
X_23005_ execute.io_target_pc\[6\] _05857_ _07091_ _07451_ _07348_ VGND VGND VPWR
+ VPWR _07452_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_60_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20217_ _05411_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28862_ clknet_leaf_176_clock _01875_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold594 fetch.bht.bhtTable_tag\[3\]\[1\] VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd3_1
X_21197_ _06086_ _05868_ net1899 VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20148_ decode.id_ex_imm_reg\[20\] _10867_ _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__a21o_1
X_27813_ clknet_leaf_320_clock _00842_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_28793_ clknet_leaf_123_clock _01806_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_202_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20079_ _00559_ _05228_ _05294_ _05231_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__o22a_1
X_24956_ csr._mcycle_T_3\[53\] _08682_ net948 VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__a21oi_1
X_27744_ clknet_leaf_34_clock _00773_ VGND VGND VPWR VPWR memory.io_wb_memtoreg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1250 fetch.bht.bhtTable_target_pc\[8\]\[17\] VGND VGND VPWR VPWR net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 fetch.bht.bhtTable_target_pc\[14\]\[28\] VGND VGND VPWR VPWR net1488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23907_ _08123_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_194_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1272 decode.regfile.registers_3\[15\] VGND VGND VPWR VPWR net1499 sky130_fd_sc_hd__dlygate4sd3_1
X_27675_ clknet_leaf_30_clock _00704_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[17\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold1283 _08373_ VGND VGND VPWR VPWR net1510 sky130_fd_sc_hd__dlygate4sd3_1
X_24887_ csr._mcycle_T_3\[32\] _08636_ _07179_ VGND VGND VPWR VPWR _08637_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_194_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1294 decode.regfile.registers_30\[18\] VGND VGND VPWR VPWR net1521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14640_ _10680_ execute.io_target_pc\[8\] _10682_ execute.io_target_pc\[15\] VGND
+ VGND VPWR VPWR _10683_ sky130_fd_sc_hd__a22oi_1
X_26626_ net1360 _09665_ _09670_ _09660_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__o211a_1
X_29414_ clknet_leaf_262_clock _02427_ VGND VGND VPWR VPWR decode.regfile.registers_5\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_23838_ _08078_ net1928 _08079_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29345_ clknet_leaf_230_clock _02358_ VGND VGND VPWR VPWR decode.regfile.registers_3\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_14571_ decode.immGen._imm_T_24\[15\] VGND VGND VPWR VPWR _10614_ sky130_fd_sc_hd__clkbuf_8
X_26557_ net870 _09622_ _09630_ _09619_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23769_ _08036_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16310_ decode.regfile.registers_2\[26\] _11369_ _11297_ _11121_ _12280_ VGND VGND
+ VPWR VPWR _12281_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_68_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13522_ fetch.bht.bhtTable_tag_MPORT_en VGND VGND VPWR VPWR _09900_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25508_ net2587 _09008_ _09012_ _09004_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29276_ clknet_leaf_243_clock _02289_ VGND VGND VPWR VPWR decode.regfile.registers_1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_17290_ decode.regfile.registers_17\[12\] _12719_ _12565_ VGND VGND VPWR VPWR _13243_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26488_ _09392_ _09589_ VGND VGND VPWR VPWR _09591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28227_ clknet_leaf_84_clock net2625 VGND VGND VPWR VPWR csr.mscratch\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16241_ _11291_ _12212_ _12213_ VGND VGND VPWR VPWR _12214_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25439_ net194 VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_180_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28158_ clknet_leaf_66_clock _01180_ VGND VGND VPWR VPWR csr.msie sky130_fd_sc_hd__dfxtp_1
X_16172_ decode.regfile.registers_8\[22\] _11045_ _11175_ VGND VGND VPWR VPWR _12147_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_209_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15123_ _10659_ decode.immGen._imm_T_24\[2\] VGND VGND VPWR VPWR _11120_ sky130_fd_sc_hd__or2_1
X_27109_ clknet_leaf_358_clock _00138_ VGND VGND VPWR VPWR decode.regfile.registers_25\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_149_Left_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28089_ clknet_leaf_167_clock _01111_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19931_ _05183_ _05197_ _05198_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__o21bai_2
X_15054_ _10660_ _10655_ VGND VGND VPWR VPWR _11051_ sky130_fd_sc_hd__nand2_2
XFILLER_0_220_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14005_ _10131_ VGND VGND VPWR VPWR _10262_ sky130_fd_sc_hd__buf_2
XFILLER_0_142_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19862_ _04508_ _04301_ _04736_ _05119_ _05132_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__o311a_1
Xoutput70 net70 VGND VGND VPWR VPWR io_fetch_address[12] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput81 net81 VGND VGND VPWR VPWR io_fetch_address[22] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput92 net92 VGND VGND VPWR VPWR io_fetch_address[3] sky130_fd_sc_hd__clkbuf_4
X_18813_ _04108_ _03914_ _03687_ decode.id_ex_rs1_data_reg\[12\] _04111_ VGND VGND
+ VPWR VPWR _04112_ sky130_fd_sc_hd__o221a_4
X_19793_ _04439_ _04679_ _05059_ _05066_ _04949_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_218_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18744_ decode.id_ex_rs1_data_reg\[5\] net246 _04042_ net355 VGND VGND VPWR VPWR
+ _04043_ sky130_fd_sc_hd__o22a_1
X_15956_ decode.regfile.registers_25\[16\] _11483_ _11484_ decode.regfile.registers_24\[16\]
+ VGND VGND VPWR VPWR _11937_ sky130_fd_sc_hd__o22a_1
XFILLER_0_204_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_158_Left_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14907_ _10939_ VGND VGND VPWR VPWR _10940_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_188_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15887_ _11679_ decode.regfile.registers_27\[14\] _11869_ VGND VGND VPWR VPWR _11870_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_78_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18675_ decode.id_ex_rs2_data_reg\[3\] net315 _03973_ VGND VGND VPWR VPWR _03974_
+ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_86_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_1290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17626_ _13451_ net668 _13492_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__o21a_1
X_14838_ csr.io_mem_pc\[8\] VGND VGND VPWR VPWR _10881_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14769_ csr.io_mem_pc\[11\] VGND VGND VPWR VPWR _10812_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17557_ decode.regfile.registers_7\[19\] _10617_ _13020_ _12843_ VGND VGND VPWR VPWR
+ _02965_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16508_ decode.regfile.registers_18\[31\] _11269_ _11271_ _12473_ VGND VGND VPWR
+ VPWR _12474_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17488_ decode.regfile.registers_16\[17\] _13011_ _13419_ _13435_ VGND VGND VPWR
+ VPWR _13436_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_15_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19227_ _04054_ net310 _04394_ _03638_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__o211ai_1
X_16439_ decode.regfile.registers_19\[29\] _11049_ _11215_ _11217_ _11454_ VGND VGND
+ VPWR VPWR _12407_ sky130_fd_sc_hd__o41a_1
XFILLER_0_128_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_167_Left_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19158_ _04332_ _04373_ net318 net257 VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18109_ _03481_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__clkbuf_1
X_19089_ _04371_ _04270_ _04372_ _04385_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__a311o_1
XFILLER_0_48_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21120_ _06052_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21051_ _06011_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20002_ _05226_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24810_ _08103_ net1652 _08585_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__mux2_1
X_25790_ net473 _09170_ _09175_ _09169_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24741_ _08103_ net1343 _06283_ VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21953_ _10130_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_2_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27460_ clknet_leaf_138_clock _00489_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[26\]
+ sky130_fd_sc_hd__dfxtp_4
X_20904_ _05931_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24672_ _08519_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21884_ csr.io_mret_vector\[14\] _10872_ _06515_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26411_ net628 _09534_ _09546_ _09540_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__o211a_1
X_23623_ _06153_ net1841 _07952_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27391_ clknet_leaf_328_clock _00420_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_20835_ net104 _05891_ _05887_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29130_ clknet_leaf_82_clock _02143_ VGND VGND VPWR VPWR csr.mcycle\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26342_ _09398_ _09502_ VGND VGND VPWR VPWR _09507_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23554_ net221 _07917_ _07921_ _05805_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20766_ _03452_ _05425_ csr.io_csr_address\[10\] VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__and3b_1
XFILLER_0_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22505_ _07098_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__buf_4
X_29061_ clknet_leaf_215_clock _02074_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_26273_ _09404_ _09459_ VGND VGND VPWR VPWR _09467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23485_ net20 _07875_ _07881_ _07879_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20697_ _05813_ decode.id_ex_rs1_data_reg\[9\] VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28012_ clknet_leaf_190_clock _01034_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25224_ _08841_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__clkbuf_1
X_22436_ _06621_ _07030_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__and2b_1
XFILLER_0_165_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25155_ _08805_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22367_ _06960_ _06961_ _06626_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24106_ net1715 execute.io_target_pc\[8\] _08221_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__mux2_1
X_21318_ _06169_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25086_ _06103_ net1539 _08596_ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__mux2_1
X_22298_ net220 _06892_ _06739_ net68 VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__a2bb2o_1
X_28914_ clknet_leaf_106_clock _01927_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_24037_ _08190_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__clkbuf_1
X_21249_ _06125_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__clkbuf_1
Xhold380 _01127_ VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold391 decode.regfile.registers_3\[10\] VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__dlygate4sd3_1
X_29894_ clknet_leaf_340_clock _02907_ VGND VGND VPWR VPWR decode.regfile.registers_20\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28845_ clknet_leaf_102_clock _01858_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_196_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15810_ _11445_ _11793_ _11794_ VGND VGND VPWR VPWR _11795_ sky130_fd_sc_hd__o21a_1
X_16790_ decode.regfile.registers_19\[1\] _12678_ _12718_ _12753_ _12544_ VGND VGND
+ VPWR VPWR _12754_ sky130_fd_sc_hd__o221a_1
X_28776_ clknet_leaf_99_clock _01789_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_25988_ _08910_ _09287_ VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_221_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15741_ decode.regfile.registers_14\[11\] _11360_ _11274_ decode.regfile.registers_15\[11\]
+ _11202_ VGND VGND VPWR VPWR _11727_ sky130_fd_sc_hd__a221o_1
X_24939_ csr._mcycle_T_3\[48\] csr._mcycle_T_3\[47\] csr._mcycle_T_3\[46\] _08668_
+ _03579_ VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__a41o_1
X_27727_ clknet_leaf_67_clock _00756_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1080 fetch.bht.bhtTable_target_pc\[4\]\[22\] VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 fetch.bht.bhtTable_target_pc\[3\]\[19\] VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15672_ decode.regfile.registers_8\[9\] _11284_ _11287_ decode.regfile.registers_9\[9\]
+ _11131_ VGND VGND VPWR VPWR _11660_ sky130_fd_sc_hd__o221a_1
X_18460_ _03758_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__buf_6
X_27658_ clknet_leaf_25_clock _00687_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ decode.control.io_opcode\[4\] _10580_ decode.control.io_opcode\[5\] VGND
+ VGND VPWR VPWR _10666_ sky130_fd_sc_hd__and3b_1
X_17411_ decode.regfile.registers_18\[15\] _12571_ _13359_ _13360_ _12561_ VGND VGND
+ VPWR VPWR _13361_ sky130_fd_sc_hd__a221o_1
XFILLER_0_197_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26609_ _09566_ VGND VGND VPWR VPWR _09660_ sky130_fd_sc_hd__clkbuf_4
X_18391_ memory.csr_read_data_out_reg\[31\] _09988_ _10144_ _10145_ VGND VGND VPWR
+ VPWR _03690_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27589_ clknet_leaf_150_clock _00618_ VGND VGND VPWR VPWR csr.io_mem_pc\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17342_ _12512_ VGND VGND VPWR VPWR _13294_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_173_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29328_ clknet_leaf_226_clock _02341_ VGND VGND VPWR VPWR decode.regfile.registers_2\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14554_ decode.immGen._imm_T_24\[18\] VGND VGND VPWR VPWR _10597_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_166_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13505_ _09886_ VGND VGND VPWR VPWR _09887_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17273_ decode.regfile.registers_4\[12\] _12618_ _12620_ decode.regfile.registers_5\[12\]
+ _12737_ VGND VGND VPWR VPWR _13226_ sky130_fd_sc_hd__a221o_1
X_29259_ clknet_leaf_233_clock _02272_ VGND VGND VPWR VPWR decode.regfile.registers_0\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_14485_ net485 _10533_ _10538_ _10535_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19012_ decode.id_ex_aluop_reg\[3\] decode.id_ex_aluop_reg\[2\] decode.id_ex_aluop_reg\[1\]
+ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__or3b_1
X_16224_ _11074_ _12196_ _12197_ _11236_ VGND VGND VPWR VPWR _12198_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer3 net229 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16155_ _11445_ _12129_ _12130_ VGND VGND VPWR VPWR _12131_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15106_ _11102_ VGND VGND VPWR VPWR _11103_ sky130_fd_sc_hd__buf_2
XFILLER_0_80_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_185_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16086_ decode.regfile.registers_4\[20\] _11410_ _12058_ _12062_ VGND VGND VPWR VPWR
+ _12063_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_107_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19914_ _05093_ _04436_ _04428_ _05181_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__o211a_1
X_15037_ _10950_ _11034_ _10969_ net470 _11004_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__o311a_1
XFILLER_0_139_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19845_ _05056_ _04261_ _04263_ _05115_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19776_ _05047_ net212 _05048_ _05049_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__and4b_1
X_16988_ _12928_ _12946_ _12852_ _12947_ VGND VGND VPWR VPWR _12948_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18727_ _03983_ _03989_ _04003_ _04006_ _04025_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_84_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15939_ decode.regfile.registers_5\[16\] _11291_ _11918_ _11919_ VGND VGND VPWR VPWR
+ _11920_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_140_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18658_ _03953_ _03954_ _03956_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_91_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17609_ decode.regfile.registers_17\[20\] _12578_ _12564_ VGND VGND VPWR VPWR _03016_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18589_ _03887_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20620_ _05541_ csr.io_mret_vector\[25\] _05602_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_175_Left_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20551_ _05577_ _05538_ _05691_ _05537_ _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__o311a_1
XFILLER_0_11_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23270_ execute.io_target_pc\[21\] _07090_ _07089_ _07701_ _06032_ VGND VGND VPWR
+ VPWR _07702_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20482_ _05632_ _05635_ _05630_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__o21a_2
X_22221_ fetch.bht.bhtTable_tag\[4\]\[20\] fetch.bht.bhtTable_tag\[5\]\[20\] fetch.bht.bhtTable_tag\[6\]\[20\]
+ fetch.bht.bhtTable_tag\[7\]\[20\] _06809_ _06649_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22152_ fetch.bht.bhtTable_tag\[8\]\[23\] fetch.bht.bhtTable_tag\[9\]\[23\] fetch.bht.bhtTable_tag\[10\]\[23\]
+ fetch.bht.bhtTable_tag\[11\]\[23\] _06618_ _06623_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__mux4_2
XFILLER_0_125_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21103_ _05856_ _06035_ _05858_ _06042_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__a31o_1
X_22083_ _06677_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__buf_4
X_26960_ _09838_ VGND VGND VPWR VPWR _09862_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_184_Left_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_353_clock clknet_5_1__leaf_clock VGND VGND VPWR VPWR clknet_leaf_353_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_7_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25911_ net2498 _09242_ _09245_ _09235_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__o211a_1
X_21034_ _05864_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26891_ _09420_ _09819_ VGND VGND VPWR VPWR _09823_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28630_ clknet_leaf_123_clock _01643_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_25842_ net1650 _09199_ _09205_ _09194_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28561_ clknet_leaf_211_clock _01574_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_25773_ net2606 _09156_ _09165_ _09153_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22985_ net94 _07343_ _07344_ _07432_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__o31a_1
XFILLER_0_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24724_ _08546_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__clkbuf_1
X_27512_ clknet_leaf_15_clock _00541_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28492_ clknet_leaf_186_clock _01505_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_21936_ csr.io_mret_vector\[30\] _10777_ _06481_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27443_ clknet_leaf_152_clock _00472_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_24655_ net1013 execute.io_target_pc\[16\] _08508_ VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__mux2_1
X_21867_ csr._mcycle_T_2\[9\] _06497_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23606_ _06136_ net2144 _07941_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_193_Left_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20818_ _05884_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__clkbuf_1
X_27374_ clknet_leaf_9_clock _00403_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_24586_ _08475_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_1188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21798_ _06457_ net217 _06458_ _06466_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__and4b_2
XFILLER_0_49_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29113_ clknet_leaf_17_clock _02126_ VGND VGND VPWR VPWR csr._mcycle_T_3\[61\] sky130_fd_sc_hd__dfxtp_1
X_26325_ _09381_ _09492_ VGND VGND VPWR VPWR _09497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23537_ _06887_ _07903_ _07911_ _07907_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_189_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20749_ _05831_ _05813_ decode.id_ex_rs1_data_reg\[31\] _05845_ _00718_ VGND VGND
+ VPWR VPWR _00750_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29044_ clknet_leaf_119_clock _02057_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14270_ _10136_ _10375_ VGND VGND VPWR VPWR _10414_ sky130_fd_sc_hd__nand2_1
X_26256_ _09387_ _09448_ VGND VGND VPWR VPWR _09457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23468_ _10981_ _07862_ _07859_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__or3b_1
XFILLER_0_150_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_306_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_306_clock
+ sky130_fd_sc_hd__clkbuf_8
X_25207_ net412 _08832_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__xnor2_1
X_22419_ _07013_ _06677_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__or2b_1
X_26187_ _10068_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__buf_4
X_23399_ fetch.bht.bhtTable_target_pc\[8\]\[30\] fetch.bht.bhtTable_target_pc\[9\]\[30\]
+ fetch.bht.bhtTable_target_pc\[10\]\[30\] fetch.bht.bhtTable_target_pc\[11\]\[30\]
+ _07106_ _07070_ VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25138_ _08797_ _03535_ decode.control.io_funct7\[5\] VGND VGND VPWR VPWR _08798_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_227_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25069_ csr._mcycle_T_2\[27\] _08712_ _08759_ csr.mcycle\[27\] VGND VGND VPWR VPWR
+ _08760_ sky130_fd_sc_hd__a211oi_1
X_17960_ decode.regfile.registers_15\[29\] _12584_ _03356_ _03357_ _13031_ VGND VGND
+ VPWR VPWR _03358_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_223_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16911_ _12707_ VGND VGND VPWR VPWR _12872_ sky130_fd_sc_hd__clkbuf_4
X_17891_ _11014_ _10936_ decode.regfile.registers_23\[27\] _12995_ VGND VGND VPWR
+ VPWR _03291_ sky130_fd_sc_hd__or4_1
X_29877_ clknet_leaf_300_clock _02890_ VGND VGND VPWR VPWR decode.regfile.registers_19\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19630_ _04887_ _04899_ _04908_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__o31ai_1
X_28828_ clknet_leaf_181_clock _01841_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16842_ decode.regfile.registers_20\[2\] _12771_ _12803_ _12804_ _12538_ VGND VGND
+ VPWR VPWR _12805_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19561_ _04211_ _04446_ _04826_ _04843_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a31o_1
X_28759_ clknet_leaf_133_clock _01772_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13985_ net1876 _10243_ _10250_ _10249_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__o211a_1
X_16773_ _12621_ VGND VGND VPWR VPWR _12737_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18512_ net196 _03772_ _03775_ _03806_ _03810_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__a2111o_1
X_15724_ _11059_ _11149_ _11128_ decode.regfile.registers_17\[10\] _11710_ VGND VGND
+ VPWR VPWR _11711_ sky130_fd_sc_hd__o221a_1
X_19492_ _04386_ _04774_ _04777_ _04295_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_17_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18443_ _03741_ decode.io_wb_rd\[2\] VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15655_ _11445_ _11642_ _11643_ _11246_ VGND VGND VPWR VPWR _11644_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14606_ _10648_ VGND VGND VPWR VPWR _10649_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_174_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15586_ decode.regfile.registers_7\[7\] _11092_ _11142_ _11165_ VGND VGND VPWR VPWR
+ _11576_ sky130_fd_sc_hd__a31o_1
X_18374_ decode.io_wb_rd\[4\] _10196_ _03672_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_145_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14537_ decode.control.io_opcode\[3\] decode.control.io_opcode\[2\] decode.control.io_opcode\[1\]
+ decode.control.io_opcode\[0\] VGND VGND VPWR VPWR _10580_ sky130_fd_sc_hd__and4bb_2
X_17325_ decode.regfile.registers_10\[13\] _12600_ _13275_ _13276_ _12724_ VGND VGND
+ VPWR VPWR _13277_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_84_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17256_ _12516_ _13207_ _13208_ _13209_ VGND VGND VPWR VPWR _13210_ sky130_fd_sc_hd__a31o_1
X_14468_ net399 _10520_ _10528_ _10522_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16207_ decode.regfile.registers_6\[23\] _10638_ _11136_ _12174_ _12180_ VGND VGND
+ VPWR VPWR _12181_ sky130_fd_sc_hd__o32a_1
XFILLER_0_141_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17187_ decode.regfile.registers_2\[10\] _12835_ _12836_ decode.regfile.registers_3\[10\]
+ _12838_ VGND VGND VPWR VPWR _13142_ sky130_fd_sc_hd__a221oi_2
XTAP_TAPCELL_ROW_133_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14399_ _10081_ _10487_ VGND VGND VPWR VPWR _10489_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_133_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16138_ _11382_ decode.regfile.registers_10\[21\] _11364_ _12113_ VGND VGND VPWR
+ VPWR _12114_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_216_Right_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_224_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16069_ decode.regfile.registers_25\[19\] _11333_ _11336_ decode.regfile.registers_24\[19\]
+ VGND VGND VPWR VPWR _12047_ sky130_fd_sc_hd__o22a_1
XFILLER_0_227_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2506 csr.mcycle\[20\] VGND VGND VPWR VPWR net2733 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2517 decode.regfile.registers_1\[18\] VGND VGND VPWR VPWR net2744 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2528 decode.regfile.registers_0\[31\] VGND VGND VPWR VPWR net2755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2539 csr._mcycle_T_3\[45\] VGND VGND VPWR VPWR net2766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1805 fetch.bht.bhtTable_tag\[15\]\[24\] VGND VGND VPWR VPWR net2032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1816 decode.regfile.registers_17\[1\] VGND VGND VPWR VPWR net2043 sky130_fd_sc_hd__dlygate4sd3_1
X_19828_ _03814_ _03829_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1827 fetch.bht.bhtTable_tag\[14\]\[3\] VGND VGND VPWR VPWR net2054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1838 decode.regfile.registers_10\[2\] VGND VGND VPWR VPWR net2065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1849 fetch.bht.bhtTable_tag\[0\]\[24\] VGND VGND VPWR VPWR net2076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19759_ _03872_ _03844_ _04307_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22770_ _07278_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21721_ net1009 _06417_ _06418_ _06419_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_91_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24440_ _08068_ net1826 _08389_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21652_ _06320_ _06365_ csr.io_inst_retired VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_192_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20603_ _05740_ _03588_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24371_ _08362_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__clkbuf_1
X_21583_ _06312_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26110_ _08956_ _09353_ VGND VGND VPWR VPWR _09360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23322_ fetch.bht.bhtTable_target_pc\[8\]\[25\] fetch.bht.bhtTable_target_pc\[9\]\[25\]
+ fetch.bht.bhtTable_target_pc\[10\]\[25\] fetch.bht.bhtTable_target_pc\[11\]\[25\]
+ _07384_ _07386_ VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20534_ csr.minstret\[13\] _05575_ _05622_ csr._csr_read_data_T_8\[13\] _05680_ VGND
+ VGND VPWR VPWR _05681_ sky130_fd_sc_hd__a221o_2
XFILLER_0_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27090_ clknet_leaf_329_clock _00119_ VGND VGND VPWR VPWR decode.regfile.registers_25\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26041_ _08962_ _09310_ VGND VGND VPWR VPWR _09320_ sky130_fd_sc_hd__nand2_1
X_23253_ csr._csr_read_data_T_8\[20\] _06480_ csr.io_mret_vector\[20\] _07621_ _07685_
+ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__o221a_1
X_20465_ _05612_ _05615_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__a21oi_4
X_22204_ _06798_ _06623_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__or2b_1
X_23184_ _10672_ VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__buf_2
X_20396_ _05534_ _05555_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__nand2_2
XFILLER_0_207_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29800_ clknet_leaf_292_clock _02813_ VGND VGND VPWR VPWR decode.regfile.registers_17\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22135_ _06649_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_292_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_292_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27992_ clknet_leaf_221_clock _01014_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29731_ clknet_leaf_291_clock _02744_ VGND VGND VPWR VPWR decode.regfile.registers_15\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_22066_ _06652_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__buf_4
X_26943_ _09838_ VGND VGND VPWR VPWR _09853_ sky130_fd_sc_hd__clkbuf_4
X_21017_ _05949_ _05945_ net479 VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__and3_1
X_29662_ clknet_leaf_288_clock _02675_ VGND VGND VPWR VPWR decode.regfile.registers_13\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26874_ net817 _09809_ _09813_ _09812_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__o211a_1
X_28613_ clknet_leaf_136_clock _01626_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25825_ _08973_ _09155_ VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__nand2_1
X_29593_ clknet_leaf_252_clock _02606_ VGND VGND VPWR VPWR decode.regfile.registers_10\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28544_ clknet_leaf_187_clock _01557_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13770_ memory.io_wb_reg_pc\[25\] _10001_ _10005_ _10109_ VGND VGND VPWR VPWR _10110_
+ sky130_fd_sc_hd__a211o_1
X_25756_ _09155_ VGND VGND VPWR VPWR _09156_ sky130_fd_sc_hd__clkbuf_4
X_22968_ _06461_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24707_ _08537_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__clkbuf_1
X_21919_ csr._mcycle_T_2\[24\] _06545_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_230_clock clknet_5_19__leaf_clock VGND VGND VPWR VPWR clknet_leaf_230_clock
+ sky130_fd_sc_hd__clkbuf_8
X_28475_ clknet_leaf_217_clock _01488_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25687_ net1757 _09111_ _09116_ _09115_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__o211a_1
X_22899_ net98 _06717_ _06698_ net225 VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15440_ decode.regfile.registers_25\[3\] _11333_ _11336_ decode.regfile.registers_24\[3\]
+ VGND VGND VPWR VPWR _11434_ sky130_fd_sc_hd__o22a_1
X_24638_ net974 execute.io_target_pc\[8\] _08497_ VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__mux2_1
X_27426_ clknet_leaf_54_clock _00455_ VGND VGND VPWR VPWR decode.id_ex_pcsel_reg sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_216_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_216_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15371_ decode.regfile.registers_8\[2\] _11285_ _11365_ decode.regfile.registers_9\[2\]
+ VGND VGND VPWR VPWR _11366_ sky130_fd_sc_hd__o22ai_1
X_24569_ _08466_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__clkbuf_1
X_27357_ clknet_leaf_49_clock _00386_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[30\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_245_clock clknet_5_25__leaf_clock VGND VGND VPWR VPWR clknet_leaf_245_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14322_ _10074_ _10444_ VGND VGND VPWR VPWR _10445_ sky130_fd_sc_hd__nand2_1
X_17110_ _12654_ _13065_ _13066_ VGND VGND VPWR VPWR _13067_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_1123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18090_ _03469_ _03467_ _03465_ net1377 VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__and4bb_1
X_26308_ net1165 _09475_ _09486_ _09484_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27288_ clknet_leaf_7_clock _00317_ VGND VGND VPWR VPWR decode.regfile.registers_31\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17041_ _12515_ _12994_ _12996_ _12999_ VGND VGND VPWR VPWR _13000_ sky130_fd_sc_hd__a31o_1
X_29027_ clknet_leaf_126_clock _02040_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_14253_ _10092_ _10400_ VGND VGND VPWR VPWR _10405_ sky130_fd_sc_hd__nand2_1
X_26239_ _09446_ VGND VGND VPWR VPWR _09447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14184_ net696 _10359_ _10364_ _10357_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18992_ _04290_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_167_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17943_ decode.regfile.registers_4\[29\] decode.regfile.registers_5\[29\] _10615_
+ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__mux2_1
X_29929_ clknet_leaf_339_clock _02942_ VGND VGND VPWR VPWR decode.regfile.registers_21\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17874_ decode.regfile.registers_4\[27\] _12548_ _12531_ decode.regfile.registers_5\[27\]
+ _12625_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19613_ _03972_ _03974_ _04007_ _04420_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_105_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16825_ decode.regfile.registers_9\[2\] _12603_ _12777_ _12787_ VGND VGND VPWR VPWR
+ _12788_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_191_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_215_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap1 _03812_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_2
X_19544_ _04095_ _04186_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_176_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16756_ decode.regfile.registers_15\[1\] _10611_ _10618_ _12588_ _12672_ VGND VGND
+ VPWR VPWR _12720_ sky130_fd_sc_hd__a41o_1
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13968_ net2637 _10200_ _10238_ _10232_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15707_ decode.regfile.registers_3\[10\] _11110_ _11141_ _11146_ VGND VGND VPWR VPWR
+ _11694_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_66_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19475_ net271 _04757_ _04760_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__o21bai_1
X_13899_ _10198_ VGND VGND VPWR VPWR _10200_ sky130_fd_sc_hd__buf_2
X_16687_ _12651_ VGND VGND VPWR VPWR _12652_ sky130_fd_sc_hd__clkbuf_4
XINSDIODE1_310 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_321 execute.io_target_pc\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_332 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18426_ net356 VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15638_ decode.regfile.registers_11\[8\] _11072_ _11205_ _11407_ _11626_ VGND VGND
+ VPWR VPWR _11627_ sky130_fd_sc_hd__a311o_1
XINSDIODE1_343 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_354 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_365 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_376 _11062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_387 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18357_ net228 VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_173_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15569_ decode.regfile.registers_21\[6\] _11267_ _11098_ _11227_ _11559_ VGND VGND
+ VPWR VPWR _11560_ sky130_fd_sc_hd__o311a_1
XFILLER_0_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17308_ net427 _12709_ _13220_ _13260_ _13219_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__o221a_1
XFILLER_0_142_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18288_ decode.id_ex_rs2_data_reg\[10\] _03605_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17239_ decode.regfile.registers_2\[11\] _12835_ _12836_ decode.regfile.registers_3\[11\]
+ _12838_ VGND VGND VPWR VPWR _13193_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold902 fetch.bht.bhtTable_target_pc\[10\]\[20\] VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold913 decode.regfile.registers_14\[16\] VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__dlygate4sd3_1
X_20250_ _05436_ _05437_ _05418_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold924 decode.regfile.registers_28\[29\] VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 fetch.bht.bhtTable_tag\[1\]\[16\] VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold946 fetch.bht.bhtTable_target_pc\[4\]\[9\] VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 fetch.bht.bhtTable_target_pc\[7\]\[20\] VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 fetch.bht.bhtTable_tag\[4\]\[11\] VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__dlygate4sd3_1
X_20181_ _05374_ _05380_ _05381_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__a21oi_1
Xhold979 csr.mscratch\[19\] VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2303 csr._minstret_T_3\[55\] VGND VGND VPWR VPWR net2530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2314 csr.mcycle\[16\] VGND VGND VPWR VPWR net2541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2325 decode.regfile.registers_19\[29\] VGND VGND VPWR VPWR net2552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23940_ _08140_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__clkbuf_1
Xhold2336 decode.id_ex_rs1_data_reg\[24\] VGND VGND VPWR VPWR net2563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1602 fetch.bht.bhtTable_target_pc\[6\]\[30\] VGND VGND VPWR VPWR net1829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2347 decode.regfile.registers_15\[24\] VGND VGND VPWR VPWR net2574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1613 fetch.bht.bhtTable_target_pc\[0\]\[14\] VGND VGND VPWR VPWR net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2358 decode.regfile.registers_11\[8\] VGND VGND VPWR VPWR net2585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 fetch.bht.bhtTable_tag\[6\]\[23\] VGND VGND VPWR VPWR net1851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 decode.regfile.registers_13\[24\] VGND VGND VPWR VPWR net2596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1635 decode.regfile.registers_27\[26\] VGND VGND VPWR VPWR net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1646 fetch.bht.bhtTable_tag\[9\]\[18\] VGND VGND VPWR VPWR net1873 sky130_fd_sc_hd__dlygate4sd3_1
X_23871_ _08101_ net2026 _07940_ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1657 fetch.bht.bhtTable_target_pc\[13\]\[17\] VGND VGND VPWR VPWR net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1668 fetch.bht.bhtTable_target_pc\[5\]\[1\] VGND VGND VPWR VPWR net1895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1679 fetch.bht.bhtTable_target_pc\[15\]\[7\] VGND VGND VPWR VPWR net1906 sky130_fd_sc_hd__dlygate4sd3_1
X_25610_ _08910_ _09069_ VGND VGND VPWR VPWR _09072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_224_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22822_ _07306_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26590_ _09420_ _09645_ VGND VGND VPWR VPWR _09650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25541_ _08916_ _09026_ VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__nand2_1
X_22753_ _07269_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21704_ csr._mcycle_T_2\[27\] _06321_ _06405_ csr.minstret\[27\] VGND VGND VPWR VPWR
+ _06406_ sky130_fd_sc_hd__a211oi_1
X_28260_ clknet_leaf_92_clock _01282_ VGND VGND VPWR VPWR csr._minstret_T_3\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_25472_ _08978_ VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22684_ net2630 _07222_ _07229_ _07221_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__o211a_1
X_24423_ _08390_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__clkbuf_1
X_27211_ clknet_leaf_364_clock _00240_ VGND VGND VPWR VPWR decode.regfile.registers_28\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28191_ clknet_leaf_113_clock _01213_ VGND VGND VPWR VPWR csr.io_mret_vector\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_21635_ csr._mcycle_T_2\[11\] _06325_ _06350_ csr.minstret\[10\] csr.minstret\[11\]
+ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_87_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27142_ clknet_leaf_359_clock _00171_ VGND VGND VPWR VPWR decode.regfile.registers_26\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_24354_ _08353_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21566_ _06303_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23305_ fetch.bht.bhtTable_target_pc\[4\]\[24\] fetch.bht.bhtTable_target_pc\[5\]\[24\]
+ fetch.bht.bhtTable_target_pc\[6\]\[24\] fetch.bht.bhtTable_target_pc\[7\]\[24\]
+ _07708_ _07103_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20517_ csr.minstret\[11\] _05573_ _05585_ csr.mcycle\[11\] _05665_ VGND VGND VPWR
+ VPWR _05666_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27073_ clknet_leaf_346_clock _00102_ VGND VGND VPWR VPWR decode.regfile.registers_24\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24285_ _08113_ net1780 _06218_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21497_ _06126_ net2066 _06263_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26024_ _09285_ VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__buf_2
X_23236_ fetch.bht.bhtTable_target_pc\[4\]\[19\] fetch.bht.bhtTable_target_pc\[5\]\[19\]
+ fetch.bht.bhtTable_target_pc\[6\]\[19\] fetch.bht.bhtTable_target_pc\[7\]\[19\]
+ _07669_ _07100_ VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20448_ csr.mcycle\[3\] _05582_ _05581_ csr.mscratch\[3\] _05604_ VGND VGND VPWR
+ VPWR _05605_ sky130_fd_sc_hd__a221o_1
X_23167_ _07602_ _07603_ _07406_ VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__mux2_1
X_20379_ _05541_ _03737_ _05516_ net358 VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_219_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22118_ _06685_ _06712_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__and2b_1
X_23098_ fetch.bht.bhtTable_target_pc\[4\]\[12\] fetch.bht.bhtTable_target_pc\[5\]\[12\]
+ fetch.bht.bhtTable_target_pc\[6\]\[12\] fetch.bht.bhtTable_target_pc\[7\]\[12\]
+ _07107_ _07114_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__mux4_1
X_27975_ clknet_leaf_210_clock _00997_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29714_ clknet_leaf_283_clock _02727_ VGND VGND VPWR VPWR decode.regfile.registers_14\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_22049_ _06643_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__clkbuf_8
X_14940_ _10968_ VGND VGND VPWR VPWR _10969_ sky130_fd_sc_hd__clkbuf_4
X_26926_ net725 _09839_ _09843_ _09836_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_162_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29645_ clknet_leaf_277_clock _02658_ VGND VGND VPWR VPWR decode.regfile.registers_12\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_14871_ _10909_ VGND VGND VPWR VPWR _10913_ sky130_fd_sc_hd__clkbuf_2
X_26857_ net1047 _09795_ _09803_ _09799_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16610_ _12574_ VGND VGND VPWR VPWR _12575_ sky130_fd_sc_hd__clkbuf_4
X_13822_ _09950_ _10154_ VGND VGND VPWR VPWR _10155_ sky130_fd_sc_hd__nand2_1
X_25808_ _08956_ _09179_ VGND VGND VPWR VPWR _09186_ sky130_fd_sc_hd__nand2_1
X_17590_ _10930_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__buf_2
X_29576_ clknet_leaf_267_clock _02589_ VGND VGND VPWR VPWR decode.regfile.registers_10\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_218_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26788_ _09389_ _09763_ VGND VGND VPWR VPWR _09764_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_218_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28527_ clknet_leaf_217_clock _01540_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16541_ _12505_ VGND VGND VPWR VPWR _12506_ sky130_fd_sc_hd__clkbuf_4
X_13753_ memory.csr_read_data_out_reg\[22\] _09989_ _10095_ VGND VGND VPWR VPWR _10096_
+ sky130_fd_sc_hd__o21ai_4
X_25739_ _08962_ _09136_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19260_ _04045_ _04054_ _03971_ _04321_ _04254_ _04352_ VGND VGND VPWR VPWR _04554_
+ sky130_fd_sc_hd__mux4_1
X_28458_ clknet_leaf_149_clock _01471_ VGND VGND VPWR VPWR decode.io_id_pc\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13684_ net594 _10027_ _10037_ _10020_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16472_ decode.regfile.registers_19\[30\] _11406_ _11325_ _12438_ VGND VGND VPWR
+ VPWR _12439_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18211_ decode.immGen._imm_T_10\[3\] _03519_ _03530_ _03547_ VGND VGND VPWR VPWR
+ _03548_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_184_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_184_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_182_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27409_ clknet_leaf_10_clock _00438_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[18\]
+ sky130_fd_sc_hd__dfxtp_4
X_15423_ _10648_ _10624_ _11085_ _11409_ _11416_ VGND VGND VPWR VPWR _11417_ sky130_fd_sc_hd__o32a_2
XFILLER_0_109_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19191_ _03986_ _03985_ _03984_ _03987_ _04070_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__a311o_1
X_28389_ clknet_leaf_58_clock _01402_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_5_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18142_ _10915_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__clkbuf_4
X_15354_ _11080_ VGND VGND VPWR VPWR _11349_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_171_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14305_ net797 _10434_ _10435_ _10427_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18073_ _10965_ _10972_ _11000_ _10018_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_53_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15285_ _11133_ VGND VGND VPWR VPWR _11281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire173 net174 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_169_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_199_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_199_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_169_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14236_ _10053_ _10387_ VGND VGND VPWR VPWR _10395_ sky130_fd_sc_hd__nand2_1
X_17024_ _12659_ _12981_ _12982_ _12664_ VGND VGND VPWR VPWR _12983_ sky130_fd_sc_hd__a211o_1
Xhold209 decode.regfile.registers_31\[22\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_1
XFILLER_0_151_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14167_ net902 _10346_ _10354_ _10344_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_91_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_122_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_122_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14098_ _10286_ VGND VGND VPWR VPWR _10315_ sky130_fd_sc_hd__clkbuf_4
X_18975_ _04230_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17926_ _12566_ _03323_ _03324_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17857_ _12968_ _03255_ _03256_ _03257_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_137_clock clknet_5_13__leaf_clock VGND VGND VPWR VPWR clknet_leaf_137_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_178_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16808_ _12770_ VGND VGND VPWR VPWR _12771_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17788_ decode.regfile.registers_3\[25\] _12836_ _10610_ _12626_ VGND VGND VPWR VPWR
+ _03190_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19527_ _04091_ net254 VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16739_ _11027_ _11015_ _11012_ _12542_ _10973_ VGND VGND VPWR VPWR _12704_ sky130_fd_sc_hd__o41a_4
XFILLER_0_18_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19458_ _04334_ net279 _04744_ _04721_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_159_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_140 _12395_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_151 _12597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_162 clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18409_ _03707_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__clkbuf_8
XINSDIODE1_173 decode.id_ex_rs2_data_reg\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19389_ _04291_ _04369_ _04358_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_184 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_195 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21420_ _06111_ net1656 _06219_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21351_ _06186_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20302_ _05476_ _05477_ _05416_ _05344_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__o2bb2a_1
X_24070_ _08207_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21282_ net1917 _06147_ _06141_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold710 decode.regfile.registers_8\[12\] VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 csr._mcycle_T_3\[54\] VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold732 fetch.bht.bhtTable_tag\[12\]\[11\] VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23021_ _07391_ _07392_ _07463_ _07466_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__a31o_1
Xhold743 fetch.bht.bhtTable_tag\[10\]\[23\] VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__dlygate4sd3_1
X_20233_ _03582_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold754 fetch.bht.bhtTable_target_pc\[1\]\[12\] VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold765 fetch.bht.bhtTable_target_pc\[12\]\[7\] VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold776 fetch.bht.bhtTable_tag\[12\]\[20\] VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold787 decode.regfile.registers_20\[31\] VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20164_ _05222_ _05367_ _05228_ _00571_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__o22a_1
Xhold798 decode.regfile.registers_19\[7\] VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2100 decode.regfile.registers_5\[11\] VGND VGND VPWR VPWR net2327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2111 decode.regfile.registers_17\[20\] VGND VGND VPWR VPWR net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2122 decode.regfile.registers_3\[25\] VGND VGND VPWR VPWR net2349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2133 decode.regfile.registers_24\[1\] VGND VGND VPWR VPWR net2360 sky130_fd_sc_hd__dlygate4sd3_1
X_27760_ clknet_leaf_322_clock _00789_ VGND VGND VPWR VPWR memory.io_wb_aluresult\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_20095_ decode.id_ex_imm_reg\[14\] decode.id_ex_pc_reg\[14\] VGND VGND VPWR VPWR
+ _05308_ sky130_fd_sc_hd__nor2_1
Xhold2144 decode.regfile.registers_7\[15\] VGND VGND VPWR VPWR net2371 sky130_fd_sc_hd__dlygate4sd3_1
X_24972_ net2365 _08693_ _08694_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__o21a_1
Xhold1410 decode.regfile.registers_22\[15\] VGND VGND VPWR VPWR net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2155 decode.regfile.registers_1\[11\] VGND VGND VPWR VPWR net2382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1421 fetch.bht.bhtTable_tag\[10\]\[11\] VGND VGND VPWR VPWR net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2166 decode.regfile.registers_14\[18\] VGND VGND VPWR VPWR net2393 sky130_fd_sc_hd__dlygate4sd3_1
X_26711_ net1194 _09709_ _09719_ _09717_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__o211a_1
X_23923_ net1296 _08081_ _08130_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1432 fetch.bht.bhtTable_tag\[10\]\[14\] VGND VGND VPWR VPWR net1659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2177 decode.regfile.registers_8\[29\] VGND VGND VPWR VPWR net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1443 fetch.bht.bhtTable_target_pc\[15\]\[12\] VGND VGND VPWR VPWR net1670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2188 csr.mcycle\[8\] VGND VGND VPWR VPWR net2415 sky130_fd_sc_hd__dlygate4sd3_1
X_27691_ clknet_leaf_24_clock _00720_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2199 decode.regfile.registers_4\[13\] VGND VGND VPWR VPWR net2426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 decode.regfile.registers_20\[6\] VGND VGND VPWR VPWR net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 fetch.bht.bhtTable_tag\[14\]\[17\] VGND VGND VPWR VPWR net1692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29430_ clknet_leaf_260_clock _02443_ VGND VGND VPWR VPWR decode.regfile.registers_5\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1476 _08481_ VGND VGND VPWR VPWR net1703 sky130_fd_sc_hd__dlygate4sd3_1
X_23854_ _08090_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__clkbuf_1
X_26642_ _09396_ _09676_ VGND VGND VPWR VPWR _09680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1487 decode.regfile.registers_7\[12\] VGND VGND VPWR VPWR net1714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1498 fetch.bht.bhtTable_target_pc\[6\]\[9\] VGND VGND VPWR VPWR net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22805_ net952 _10868_ _07297_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29361_ clknet_leaf_227_clock _02374_ VGND VGND VPWR VPWR decode.regfile.registers_3\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_23785_ _06147_ net2121 _08041_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__mux2_1
X_26573_ _09402_ _09632_ VGND VGND VPWR VPWR _09640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20997_ execute.io_reg_pc\[23\] _05977_ _05973_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__and3_1
XFILLER_0_223_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28312_ clknet_leaf_220_clock _01325_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22736_ _07260_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__clkbuf_1
X_25524_ _08975_ _08978_ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_213_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29292_ clknet_leaf_231_clock _02305_ VGND VGND VPWR VPWR decode.regfile.registers_1\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28243_ clknet_leaf_77_clock _01265_ VGND VGND VPWR VPWR csr._minstret_T_3\[43\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_48_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25455_ net211 VGND VGND VPWR VPWR _08982_ sky130_fd_sc_hd__buf_4
XFILLER_0_165_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22667_ net2568 _07208_ _07219_ _07164_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24406_ _08380_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__clkbuf_1
X_21618_ net2676 _06329_ _06340_ csr.minstret\[6\] VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_192_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28174_ clknet_leaf_57_clock _01196_ VGND VGND VPWR VPWR csr.io_mret_vector\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_25386_ _08933_ _08923_ VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__nand2_1
X_22598_ csr._minstret_T_3\[47\] _07174_ _07175_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_124_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24337_ _08099_ net1819 _06187_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27125_ clknet_leaf_351_clock _00154_ VGND VGND VPWR VPWR decode.regfile.registers_26\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_21549_ _06294_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15070_ _11066_ VGND VGND VPWR VPWR _11067_ sky130_fd_sc_hd__buf_4
X_27056_ clknet_leaf_330_clock _00085_ VGND VGND VPWR VPWR decode.regfile.registers_24\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24268_ _08309_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14021_ net1866 _10258_ _10270_ _10262_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__o211a_1
X_26007_ _08929_ _09297_ VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23219_ _07651_ _07652_ _07063_ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__and3b_1
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24199_ _08093_ net1713 _08266_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_207_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18760_ execute.io_reg_pc\[7\] _03777_ _03665_ net129 _04058_ VGND VGND VPWR VPWR
+ _04059_ sky130_fd_sc_hd__o221a_1
X_27958_ clknet_leaf_186_clock _00980_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_160_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ _11042_ decode.regfile.registers_4\[17\] VGND VGND VPWR VPWR _11952_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_54_clock
+ sky130_fd_sc_hd__clkbuf_8
X_17711_ decode.regfile.registers_13\[23\] _12927_ _12588_ _12663_ VGND VGND VPWR
+ VPWR _03115_ sky130_fd_sc_hd__a31o_1
X_14923_ decode.control.io_opcode\[5\] _10951_ VGND VGND VPWR VPWR _10952_ sky130_fd_sc_hd__nor2_2
X_26909_ net2355 _09822_ _09832_ _09825_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18691_ net208 net206 net236 _03598_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_136_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27889_ clknet_leaf_24_clock _00918_ VGND VGND VPWR VPWR csr._mcycle_T_2\[10\] sky130_fd_sc_hd__dfxtp_2
X_17642_ decode.regfile.registers_11\[21\] _12724_ _12722_ _12540_ VGND VGND VPWR
+ VPWR _03048_ sky130_fd_sc_hd__o2bb2a_1
X_29628_ clknet_leaf_288_clock _02641_ VGND VGND VPWR VPWR decode.regfile.registers_12\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14854_ _10680_ _10884_ _10885_ _10886_ _10896_ VGND VGND VPWR VPWR _10897_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_216_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13805_ memory.io_wb_readdata\[30\] _10004_ _10139_ VGND VGND VPWR VPWR _10140_ sky130_fd_sc_hd__a21o_1
X_17573_ decode.regfile.registers_22\[19\] _12527_ _02979_ _02980_ _12686_ VGND VGND
+ VPWR VPWR _02981_ sky130_fd_sc_hd__a221o_1
X_29559_ clknet_leaf_274_clock _02572_ VGND VGND VPWR VPWR decode.regfile.registers_9\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14785_ csr.io_mem_pc\[2\] csr.io_mem_pc\[3\] csr.io_mem_pc\[4\] VGND VGND VPWR VPWR
+ _10828_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_69_clock clknet_5_2__leaf_clock VGND VGND VPWR VPWR clknet_leaf_69_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19312_ _04601_ _04604_ _04415_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_158_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16524_ _12488_ VGND VGND VPWR VPWR _12489_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_158_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13736_ _10081_ _10075_ VGND VGND VPWR VPWR _10082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19243_ _03704_ _04537_ _04270_ _04536_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__a31o_1
X_16455_ decode.regfile.registers_3\[30\] _11110_ _11141_ _11145_ VGND VGND VPWR VPWR
+ _12422_ sky130_fd_sc_hd__a31o_1
X_13667_ _10012_ memory.io_wb_aluresult\[9\] _09978_ memory.io_wb_reg_pc\[9\] _09995_
+ VGND VGND VPWR VPWR _10023_ sky130_fd_sc_hd__a221o_2
X_15406_ _11346_ _11253_ _11064_ decode.regfile.registers_29\[2\] _11400_ VGND VGND
+ VPWR VPWR _11401_ sky130_fd_sc_hd__o221a_1
X_19174_ _04279_ _04019_ _04469_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_22_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16386_ _12353_ _11369_ _11614_ _12354_ VGND VGND VPWR VPWR _12355_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_22_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13598_ _09960_ _09961_ memory.io_wb_reg_pc\[1\] VGND VGND VPWR VPWR _09962_ sky130_fd_sc_hd__o21a_1
XFILLER_0_183_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18125_ _03490_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15337_ _11332_ VGND VGND VPWR VPWR _11333_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18056_ _09954_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 _00701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15268_ _10977_ VGND VGND VPWR VPWR _11264_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17007_ _10930_ decode.regfile.registers_28\[6\] _12698_ VGND VGND VPWR VPWR _12966_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14219_ net688 _10376_ _10384_ _10385_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__o211a_1
X_15199_ _11195_ VGND VGND VPWR VPWR _11196_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18958_ _03918_ _04255_ _04256_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_52_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17909_ decode.regfile.registers_2\[28\] _12834_ net209 decode.regfile.registers_3\[28\]
+ _12837_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__a221oi_1
X_18889_ _04121_ _04179_ _04184_ _04187_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_206_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20920_ _05940_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer13 _03757_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__buf_1
Xrebuffer24 net252 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer35 net261 VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_1
Xrebuffer46 net204 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__buf_1
XFILLER_0_156_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20851_ _05902_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer57 net283 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer68 net293 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_1
Xrebuffer79 _03752_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23570_ _07929_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__clkbuf_8
X_20782_ _03590_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22521_ _07114_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__buf_4
XFILLER_0_187_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25240_ _08078_ net1542 _08848_ VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22452_ _07044_ _07046_ _06623_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer103 _09921_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21403_ _06151_ net2053 _06210_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__mux2_1
Xrebuffer114 _08633_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__buf_1
X_25171_ net413 _08814_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22383_ fetch.bht.bhtTable_tag\[6\]\[9\] fetch.bht.bhtTable_tag\[7\]\[9\] _06617_
+ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24122_ _08234_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__clkbuf_1
X_21334_ _06177_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24053_ net1069 execute.io_target_pc\[14\] _08198_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__mux2_1
X_28930_ clknet_leaf_135_clock _01943_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21265_ csr.io_mem_pc\[23\] VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__buf_2
Xhold540 fetch.bht.bhtTable_target_pc\[12\]\[21\] VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _01226_ VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold562 fetch.bht.bhtTable_tag\[3\]\[3\] VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__dlygate4sd3_1
X_23004_ csr._csr_read_data_T_8\[6\] _06038_ csr.io_mret_vector\[6\] _06462_ VGND
+ VGND VPWR VPWR _07451_ sky130_fd_sc_hd__a22o_1
X_20216_ decode.id_ex_rdsel_reg VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold573 decode.regfile.registers_6\[16\] VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28861_ clknet_leaf_178_clock _01874_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold584 decode.regfile.registers_4\[3\] VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd3_1
X_21196_ _06093_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__clkbuf_1
Xhold595 decode.regfile.registers_31\[20\] VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__buf_1
XFILLER_0_204_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27812_ clknet_leaf_35_clock _00841_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20147_ _05341_ _05347_ _05345_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__and3_1
X_28792_ clknet_leaf_121_clock _01805_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_202_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27743_ clknet_leaf_35_clock _00772_ VGND VGND VPWR VPWR memory.io_wb_memtoreg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_20078_ _05290_ _05293_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__and2_1
X_24955_ net2638 _08682_ _08683_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__o21a_1
Xhold1240 decode.regfile.registers_5\[4\] VGND VGND VPWR VPWR net1467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1251 _08372_ VGND VGND VPWR VPWR net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 fetch.bht.bhtTable_target_pc\[13\]\[19\] VGND VGND VPWR VPWR net1489 sky130_fd_sc_hd__dlygate4sd3_1
X_23906_ net752 _08064_ _08119_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__mux2_1
Xhold1273 fetch.bht.bhtTable_target_pc\[12\]\[22\] VGND VGND VPWR VPWR net1500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27674_ clknet_leaf_31_clock _00703_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[16\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold1284 fetch.bht.bhtTable_target_pc\[10\]\[13\] VGND VGND VPWR VPWR net1511 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24886_ csr.mcycle\[31\] _08628_ _08632_ _08635_ VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__and4_2
XFILLER_0_224_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 fetch.bht.bhtTable_target_pc\[9\]\[29\] VGND VGND VPWR VPWR net1522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29413_ clknet_leaf_257_clock _02426_ VGND VGND VPWR VPWR decode.regfile.registers_5\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_26625_ _09379_ _09666_ VGND VGND VPWR VPWR _09670_ sky130_fd_sc_hd__nand2_1
X_23837_ _07929_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_185_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29344_ clknet_leaf_230_clock _02357_ VGND VGND VPWR VPWR decode.regfile.registers_3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14570_ decode.id_ex_ex_rd_reg\[1\] VGND VGND VPWR VPWR _10613_ sky130_fd_sc_hd__inv_2
XFILLER_0_196_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23768_ _06130_ net1320 _08030_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__mux2_1
X_26556_ _09385_ _09623_ VGND VGND VPWR VPWR _09630_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13521_ _09899_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__clkbuf_1
X_25507_ _08958_ _09005_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29275_ clknet_leaf_241_clock _02288_ VGND VGND VPWR VPWR decode.regfile.registers_1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_22719_ decode.control.io_funct3\[0\] _10943_ decode.control.io_funct3\[2\] VGND
+ VGND VPWR VPWR _07250_ sky130_fd_sc_hd__and3b_1
X_23699_ net1186 _10871_ _07992_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__mux2_1
X_26487_ net624 _09578_ _09590_ _09582_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28226_ clknet_leaf_87_clock net2159 VGND VGND VPWR VPWR csr.mscratch\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16240_ decode.regfile.registers_5\[24\] _11313_ _11410_ _11462_ _11314_ VGND VGND
+ VPWR VPWR _12213_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_153_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25438_ net2408 _08951_ _08969_ _08950_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25369_ net2434 _08906_ _08921_ _07247_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__o211a_1
X_28157_ clknet_leaf_66_clock _01179_ VGND VGND VPWR VPWR csr.msip sky130_fd_sc_hd__dfxtp_1
X_16171_ _11136_ _12144_ _12145_ VGND VGND VPWR VPWR _12146_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27108_ clknet_leaf_348_clock _00137_ VGND VGND VPWR VPWR decode.regfile.registers_25\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_15122_ _11118_ VGND VGND VPWR VPWR _11119_ sky130_fd_sc_hd__clkbuf_4
X_28088_ clknet_leaf_195_clock _01110_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19930_ _04317_ _04439_ _04468_ _04949_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__a31o_1
X_15053_ _11049_ VGND VGND VPWR VPWR _11050_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27039_ clknet_leaf_345_clock _00068_ VGND VGND VPWR VPWR decode.regfile.registers_23\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14004_ _10042_ _10255_ VGND VGND VPWR VPWR _10261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19861_ _04620_ _05120_ _05121_ _05131_ _04301_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__o221ai_4
Xoutput71 net71 VGND VGND VPWR VPWR io_fetch_address[13] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput82 net82 VGND VGND VPWR VPWR io_fetch_address[23] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18812_ _03768_ _03769_ _03770_ _04110_ _03669_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__o41a_2
Xoutput93 net93 VGND VGND VPWR VPWR io_fetch_address[4] sky130_fd_sc_hd__clkbuf_4
X_19792_ _04675_ _04924_ _04360_ _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18743_ memory.csr_read_data_out_reg\[5\] _10010_ _09991_ VGND VGND VPWR VPWR _04042_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_218_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15955_ decode.regfile.registers_23\[16\] _11088_ _11912_ _11935_ VGND VGND VPWR
+ VPWR _11936_ sky130_fd_sc_hd__o22a_1
XFILLER_0_223_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14906_ _10938_ VGND VGND VPWR VPWR _10939_ sky130_fd_sc_hd__clkbuf_4
X_18674_ net208 net206 _09974_ _03879_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__o211ai_2
X_15886_ _11257_ VGND VGND VPWR VPWR _11869_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ net822 _12872_ _02996_ _03031_ _13219_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__o221a_1
X_14837_ _10763_ _10879_ VGND VGND VPWR VPWR _10880_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17556_ decode.regfile.registers_6\[19\] _10602_ _12626_ _12645_ VGND VGND VPWR VPWR
+ _02964_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_82_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14768_ _10810_ decode.id_ex_pc_reg\[13\] VGND VGND VPWR VPWR _10811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16507_ _11357_ _12471_ _12472_ VGND VGND VPWR VPWR _12473_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13719_ _10003_ memory.io_wb_aluresult\[17\] _10004_ memory.io_wb_readdata\[17\]
+ _09995_ VGND VGND VPWR VPWR _10067_ sky130_fd_sc_hd__a221oi_2
X_17487_ decode.regfile.registers_14\[17\] _12984_ _13420_ _13434_ _12874_ VGND VGND
+ VPWR VPWR _13435_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_15_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14699_ execute.io_target_pc\[20\] _10716_ execute.io_target_pc\[17\] _10736_ VGND
+ VGND VPWR VPWR _10742_ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19226_ _04519_ _04518_ _04039_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_229_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16438_ _11106_ _12404_ _12405_ VGND VGND VPWR VPWR _12406_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19157_ net213 VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__clkbuf_4
X_16369_ _11076_ _11090_ decode.regfile.registers_25\[27\] _12311_ _12338_ VGND VGND
+ VPWR VPWR _12339_ sky130_fd_sc_hd__o32a_1
XFILLER_0_6_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18108_ _03469_ _03480_ _03474_ decode.io_id_pc\[11\] VGND VGND VPWR VPWR _03481_
+ sky130_fd_sc_hd__and4bb_1
X_19088_ _04297_ decode.id_ex_imm_reg\[4\] _04035_ _04298_ _04306_ VGND VGND VPWR
+ VPWR _04386_ sky130_fd_sc_hd__a221o_4
XFILLER_0_48_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18039_ decode.regfile.registers_21\[31\] _12822_ _12909_ VGND VGND VPWR VPWR _03435_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21050_ execute.csr_read_data_out_reg\[14\] _06002_ _06010_ VGND VGND VPWR VPWR _06011_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_100_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20001_ _05222_ _05225_ _05227_ _00548_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__o22a_1
XFILLER_0_226_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24740_ _08554_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__clkbuf_1
X_21952_ net1913 _06574_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20903_ _05925_ _05921_ net37 VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__and3_1
X_24671_ net929 execute.io_target_pc\[24\] _07285_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21883_ _06527_ _06519_ _06520_ _06528_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23622_ _07957_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__clkbuf_1
X_26410_ _09389_ _09545_ VGND VGND VPWR VPWR _09546_ sky130_fd_sc_hd__nand2_1
X_20834_ _05893_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__clkbuf_1
X_27390_ clknet_leaf_9_clock _00419_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[31\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23553_ net2138 _07918_ _07915_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__or3b_1
XFILLER_0_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26341_ net727 _09505_ _09506_ _09499_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20765_ _05851_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22504_ _07066_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__buf_4
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29060_ clknet_leaf_223_clock _02073_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_26272_ net2264 _09462_ _09466_ _09458_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23484_ decode.control.io_funct7\[2\] _07876_ _07873_ VGND VGND VPWR VPWR _07881_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_169_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20696_ _05804_ _00695_ _05814_ net183 net700 VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25223_ _08062_ net1768 _08837_ VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__mux2_1
X_28011_ clknet_leaf_189_clock _01033_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22435_ fetch.bht.bhtTable_tag\[8\]\[12\] fetch.bht.bhtTable_tag\[9\]\[12\] net300
+ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25154_ _10573_ net2635 _08804_ VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22366_ fetch.bht.bhtTable_tag\[8\]\[2\] fetch.bht.bhtTable_tag\[9\]\[2\] fetch.bht.bhtTable_tag\[10\]\[2\]
+ fetch.bht.bhtTable_tag\[11\]\[2\] net303 _06620_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__mux4_1
X_24105_ _08225_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__clkbuf_1
X_21317_ net1655 _10868_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25085_ _08770_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__clkbuf_1
X_22297_ _06641_ _06838_ _06842_ _06848_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__o31a_1
XFILLER_0_130_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28913_ clknet_leaf_105_clock _01926_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_24036_ net1711 execute.io_target_pc\[6\] _08187_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21248_ net1043 _06124_ _06120_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold370 decode.regfile.registers_12\[8\] VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__dlygate4sd3_1
X_29893_ clknet_leaf_302_clock _02906_ VGND VGND VPWR VPWR decode.regfile.registers_20\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold381 decode.regfile.registers_28\[31\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold392 decode.regfile.registers_6\[9\] VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_225_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28844_ clknet_leaf_109_clock _01857_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_21179_ _06084_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_196_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28775_ clknet_leaf_119_clock _01788_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25987_ net2719 _09286_ _09289_ _09277_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_221_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27726_ clknet_leaf_69_clock _00755_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_15740_ decode.regfile.registers_19\[11\] _11271_ _11101_ VGND VGND VPWR VPWR _11726_
+ sky130_fd_sc_hd__a21o_1
X_24938_ csr._mcycle_T_3\[47\] csr._mcycle_T_3\[46\] _08668_ VGND VGND VPWR VPWR _08672_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_172_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1070 decode.regfile.registers_29\[29\] VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 fetch.bht.bhtTable_target_pc\[3\]\[31\] VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1092 fetch.bht.bhtTable_target_pc\[7\]\[3\] VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15671_ _11652_ _11658_ _11318_ _11084_ VGND VGND VPWR VPWR _11659_ sky130_fd_sc_hd__o2bb2a_1
X_27657_ clknet_leaf_38_clock _00686_ VGND VGND VPWR VPWR execute.io_mret_out sky130_fd_sc_hd__dfxtp_1
X_24869_ _08622_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_213_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ decode.regfile.registers_17\[15\] _12579_ _12565_ VGND VGND VPWR VPWR _13360_
+ sky130_fd_sc_hd__o21a_1
X_14622_ decode.control.io_opcode\[6\] _10578_ VGND VGND VPWR VPWR _10665_ sky130_fd_sc_hd__nor2_1
X_26608_ _09438_ _09621_ VGND VGND VPWR VPWR _09659_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _03688_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__buf_8
X_27588_ clknet_leaf_136_clock _00617_ VGND VGND VPWR VPWR csr.io_mem_pc\[29\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_157_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29327_ clknet_leaf_226_clock _02340_ VGND VGND VPWR VPWR decode.regfile.registers_2\[21\]
+ sky130_fd_sc_hd__dfxtp_2
X_17341_ _12516_ _13290_ _13291_ _13292_ VGND VGND VPWR VPWR _13293_ sky130_fd_sc_hd__a31o_1
X_26539_ net2203 _09579_ _09618_ _09619_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14553_ net2181 VGND VGND VPWR VPWR _10596_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13504_ csr.io_mem_pc\[2\] csr.io_mem_pc\[3\] VGND VGND VPWR VPWR _09886_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29258_ clknet_leaf_224_clock _02271_ VGND VGND VPWR VPWR decode.regfile.registers_0\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_17272_ decode.regfile.registers_9\[12\] _12603_ _12790_ VGND VGND VPWR VPWR _13225_
+ sky130_fd_sc_hd__o21ai_1
X_14484_ _10102_ _10530_ VGND VGND VPWR VPWR _10538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19011_ decode.id_ex_imm_reg\[0\] _03726_ _03669_ _04229_ _04309_ VGND VGND VPWR
+ VPWR _04310_ sky130_fd_sc_hd__o2111a_1
X_28209_ clknet_leaf_61_clock net1937 VGND VGND VPWR VPWR csr.mscratch\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16223_ decode.regfile.registers_25\[23\] _11483_ _11484_ decode.regfile.registers_24\[23\]
+ VGND VGND VPWR VPWR _12197_ sky130_fd_sc_hd__o22a_1
XFILLER_0_153_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29189_ clknet_leaf_164_clock _02202_ VGND VGND VPWR VPWR fetch.btb.btbTable\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer4 net228 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_1
X_16154_ _11489_ decode.regfile.registers_28\[21\] decode.regfile.registers_29\[21\]
+ _11063_ _11245_ VGND VGND VPWR VPWR _12130_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_185_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15105_ _11101_ VGND VGND VPWR VPWR _11102_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_185_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16085_ decode.regfile.registers_2\[20\] _10647_ _11148_ _11152_ _12061_ VGND VGND
+ VPWR VPWR _12062_ sky130_fd_sc_hd__o311a_1
XFILLER_0_107_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19913_ _04244_ _05008_ _05180_ _04305_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__o2bb2a_1
X_15036_ _10965_ _10964_ _10951_ VGND VGND VPWR VPWR _11034_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_220_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1096 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19844_ net188 net189 _04274_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19775_ _03849_ _05045_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_144_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16987_ decode.regfile.registers_14\[5\] _10603_ _10618_ _12722_ VGND VGND VPWR VPWR
+ _12947_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18726_ _04009_ _04024_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15938_ _11313_ decode.regfile.registers_4\[16\] _10647_ _10630_ _11462_ VGND VGND
+ VPWR VPWR _11919_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_140_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18657_ _10086_ _03771_ _03774_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_204_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15869_ decode.regfile.registers_8\[14\] _11175_ _11365_ _11851_ VGND VGND VPWR VPWR
+ _11852_ sky130_fd_sc_hd__o211a_1
X_17608_ decode.regfile.registers_16\[20\] _12575_ _02999_ _03014_ VGND VGND VPWR
+ VPWR _03015_ sky130_fd_sc_hd__o22a_1
XFILLER_0_171_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18588_ _03688_ decode.id_ex_rs1_data_reg\[22\] _03700_ _03883_ _03886_ VGND VGND
+ VPWR VPWR _03887_ sky130_fd_sc_hd__o221a_1
XFILLER_0_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17539_ _13183_ _13481_ _13483_ _13485_ VGND VGND VPWR VPWR _13486_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_43_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20550_ csr._csr_read_data_T_8\[15\] _05617_ _05693_ _05694_ VGND VGND VPWR VPWR
+ _05695_ sky130_fd_sc_hd__a211o_1
XFILLER_0_229_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19209_ _04504_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20481_ net2517 _05593_ _05625_ _05633_ _05634_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__o32a_1
XFILLER_0_73_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22220_ _06812_ _06813_ _06675_ _06814_ _06627_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_42_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22151_ _06661_ _06743_ _06629_ _06745_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_140_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21102_ execute.exception_out_reg _06033_ net329 net132 VGND VGND VPWR VPWR _06042_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_218_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22082_ _06620_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21033_ _06001_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
X_25910_ _08982_ _09243_ VGND VGND VPWR VPWR _09245_ sky130_fd_sc_hd__nand2_1
X_26890_ _09794_ VGND VGND VPWR VPWR _09822_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25841_ _08914_ _09200_ VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28560_ clknet_leaf_207_clock _01573_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_22984_ _07348_ _07431_ _10019_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__o21a_1
X_25772_ _08920_ _09157_ VGND VGND VPWR VPWR _09165_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27511_ clknet_leaf_15_clock _00540_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dfxtp_1
X_24723_ _08085_ net1884 _08542_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28491_ clknet_leaf_202_clock _01504_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_21935_ _06563_ _06543_ _06544_ _06564_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27442_ clknet_leaf_153_clock _00471_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_24654_ _08510_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21866_ csr.io_mret_vector\[9\] _10817_ _06515_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23605_ _07948_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20817_ net127 _05879_ _05875_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__and3_1
X_27373_ clknet_leaf_9_clock _00402_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_24585_ net1430 execute.io_target_pc\[14\] _08473_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__mux2_1
X_21797_ csr.io_csr_write_address\[1\] csr.io_csr_write_address\[3\] csr.io_csr_write_address\[2\]
+ csr.io_csr_write_enable VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29112_ clknet_leaf_17_clock _02125_ VGND VGND VPWR VPWR csr._mcycle_T_3\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26324_ net766 _09491_ _09496_ _09484_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23536_ net2305 _07904_ _07901_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_150_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20748_ _05818_ decode.id_ex_rs1_data_reg\[31\] _03585_ VGND VGND VPWR VPWR _05845_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_189_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_189_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29043_ clknet_leaf_133_clock _02056_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_23467_ net13 _07861_ _07870_ _07865_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__o211a_1
X_26255_ net718 _09447_ _09456_ _09440_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20679_ _00690_ _05803_ _05801_ _05802_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22418_ fetch.bht.bhtTable_tag\[14\]\[1\] fetch.bht.bhtTable_tag\[15\]\[1\] net298
+ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__mux2_1
X_25206_ _10568_ _10815_ VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23398_ fetch.bht.bhtTable_target_pc\[12\]\[30\] fetch.bht.bhtTable_target_pc\[13\]\[30\]
+ fetch.bht.bhtTable_target_pc\[14\]\[30\] fetch.bht.bhtTable_target_pc\[15\]\[30\]
+ _07106_ _07386_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__mux4_1
X_26186_ net2591 _09395_ _09409_ _09394_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_5_11__f_clock clknet_2_1_0_clock VGND VGND VPWR VPWR clknet_5_11__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_122_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22349_ net74 _06943_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__xnor2_1
X_25137_ _03526_ net214 _03524_ _07250_ VGND VGND VPWR VPWR _08797_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_227_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25068_ _06331_ _08758_ _08759_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__nor3_1
X_29945_ clknet_leaf_335_clock _02958_ VGND VGND VPWR VPWR decode.regfile.registers_21\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_223_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_223_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24019_ net1123 execute.io_target_pc\[30\] _07960_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__mux2_1
X_16910_ net918 _12709_ _12821_ _12871_ _12705_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__o221a_1
X_17890_ decode.regfile.registers_22\[27\] _13100_ _03289_ _13289_ VGND VGND VPWR
+ VPWR _03290_ sky130_fd_sc_hd__a211o_1
X_29876_ clknet_leaf_300_clock _02889_ VGND VGND VPWR VPWR decode.regfile.registers_19\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28827_ clknet_leaf_173_clock _01840_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_16841_ decode.regfile.registers_19\[2\] _11013_ _11012_ _12519_ _12545_ VGND VGND
+ VPWR VPWR _12804_ sky130_fd_sc_hd__o41a_1
XFILLER_0_219_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19560_ _04832_ _04833_ _04842_ _04505_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__o211a_1
X_28758_ clknet_leaf_126_clock _01771_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16772_ _12727_ _12734_ _12735_ VGND VGND VPWR VPWR _12736_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_107_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13984_ _09975_ _10244_ VGND VGND VPWR VPWR _10250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18511_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__inv_2
X_15723_ _11203_ _11708_ _11709_ VGND VGND VPWR VPWR _11710_ sky130_fd_sc_hd__o21ai_1
X_27709_ clknet_leaf_19_clock _00738_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_19491_ _04539_ _04775_ _04776_ _04492_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28689_ clknet_leaf_104_clock _01702_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ csr.io_csr_address\[2\] VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__inv_2
X_15654_ _11396_ decode.regfile.registers_28\[8\] decode.regfile.registers_29\[8\]
+ _11255_ VGND VGND VPWR VPWR _11643_ sky130_fd_sc_hd__o22a_1
XFILLER_0_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_90 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14605_ _10647_ VGND VGND VPWR VPWR _10648_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_174_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ decode.io_wb_rd\[2\] decode.io_wb_rd\[3\] VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nor2_8
XFILLER_0_84_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15585_ decode.regfile.registers_9\[7\] _11280_ _11281_ _11183_ VGND VGND VPWR VPWR
+ _11575_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17324_ decode.regfile.registers_9\[13\] _11018_ _12977_ _12510_ _12653_ VGND VGND
+ VPWR VPWR _13276_ sky130_fd_sc_hd__o41a_1
X_14536_ decode.control.io_opcode\[6\] VGND VGND VPWR VPWR _10579_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17255_ _10927_ decode.regfile.registers_24\[11\] _13170_ _13083_ _12862_ VGND VGND
+ VPWR VPWR _13209_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_4_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14467_ _10064_ _10517_ VGND VGND VPWR VPWR _10528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16206_ _12175_ _12178_ _12179_ VGND VGND VPWR VPWR _12180_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_948 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17186_ decode.regfile.registers_7\[10\] _12610_ _12622_ decode.regfile.registers_6\[10\]
+ VGND VGND VPWR VPWR _13141_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14398_ net1521 _10477_ _10488_ _10481_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_180_Right_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16137_ decode.regfile.registers_9\[21\] _11547_ _12111_ _12112_ _11509_ VGND VGND
+ VPWR VPWR _12113_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16068_ _10992_ _11066_ _11261_ _12045_ VGND VGND VPWR VPWR _12046_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15019_ _10998_ VGND VGND VPWR VPWR _11028_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2507 decode.regfile.registers_10\[25\] VGND VGND VPWR VPWR net2734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2518 decode.regfile.registers_2\[8\] VGND VGND VPWR VPWR net2745 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2529 decode.regfile.registers_7\[25\] VGND VGND VPWR VPWR net2756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1806 decode.regfile.registers_13\[17\] VGND VGND VPWR VPWR net2033 sky130_fd_sc_hd__dlygate4sd3_1
X_19827_ _05098_ _03639_ _04667_ _03829_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__a211o_1
Xhold1817 fetch.bht.bhtTable_tag\[7\]\[19\] VGND VGND VPWR VPWR net2044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1828 fetch.bht.bhtTable_tag\[5\]\[4\] VGND VGND VPWR VPWR net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1839 fetch.bht.bhtTable_tag\[5\]\[12\] VGND VGND VPWR VPWR net2066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_224_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19758_ _05029_ _05030_ _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_79_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18709_ _03972_ _03974_ _04007_ _03971_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19689_ _04546_ _04556_ _04879_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21720_ _03579_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21651_ csr.minstret\[14\] _06333_ _06355_ _06360_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__nand4_2
XFILLER_0_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20602_ _03555_ _05588_ _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24370_ net1037 execute.io_target_pc\[8\] _08356_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21582_ _06153_ net1706 _06306_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23321_ fetch.bht.bhtTable_target_pc\[12\]\[25\] fetch.bht.bhtTable_target_pc\[13\]\[25\]
+ fetch.bht.bhtTable_target_pc\[14\]\[25\] fetch.bht.bhtTable_target_pc\[15\]\[25\]
+ _07384_ _07386_ VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_25_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20533_ csr._minstret_T_3\[45\] _05577_ _05578_ _05552_ csr.mcycle\[13\] VGND VGND
+ VPWR VPWR _05680_ sky130_fd_sc_hd__a32o_1
XFILLER_0_145_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23252_ _07064_ _07676_ _07677_ _07684_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__a31o_1
X_26040_ net2627 _09313_ _09319_ _09318_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20464_ csr._minstret_T_3\[36\] _05616_ _05618_ csr._csr_read_data_T_8\[4\] _05619_
+ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22203_ fetch.bht.bhtTable_tag\[6\]\[24\] fetch.bht.bhtTable_tag\[7\]\[24\] _06700_
+ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23183_ _05864_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20395_ net294 _05525_ _05536_ _05540_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__and4_2
X_22134_ fetch.bht.bhtTable_tag\[6\]\[4\] fetch.bht.bhtTable_tag\[7\]\[4\] _06643_
+ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27991_ clknet_leaf_233_clock _01013_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29730_ clknet_leaf_291_clock _02743_ VGND VGND VPWR VPWR decode.regfile.registers_15\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_22065_ _06619_ fetch.bht.bhtTable_tag\[7\]\[18\] _06652_ VGND VGND VPWR VPWR _06660_
+ sky130_fd_sc_hd__a21bo_1
X_26942_ net2116 _09839_ _09851_ _09852_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21016_ _05992_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__clkbuf_1
X_29661_ clknet_leaf_287_clock _02674_ VGND VGND VPWR VPWR decode.regfile.registers_13\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26873_ _09400_ _09806_ VGND VGND VPWR VPWR _09813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28612_ clknet_leaf_132_clock _01625_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_25824_ net1597 _09183_ _09193_ _09194_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29592_ clknet_leaf_312_clock _02605_ VGND VGND VPWR VPWR decode.regfile.registers_10\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28543_ clknet_leaf_200_clock _01556_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_25755_ _09154_ VGND VGND VPWR VPWR _09155_ sky130_fd_sc_hd__clkbuf_4
X_22967_ net93 _07343_ _07344_ _07415_ _06566_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__o311a_1
XFILLER_0_134_1218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24706_ _08068_ net1081 _08531_ VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21918_ csr.io_mret_vector\[24\] _10772_ _06539_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__mux2_1
X_28474_ clknet_leaf_161_clock _01487_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25686_ _08910_ _09112_ VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22898_ _06820_ _07037_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27425_ clknet_leaf_53_clock _00454_ VGND VGND VPWR VPWR decode.id_ex_rdsel_reg sky130_fd_sc_hd__dfxtp_4
XFILLER_0_210_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24637_ _08501_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__clkbuf_1
X_21849_ _06503_ _06494_ _06495_ _06504_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_216_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_216_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_43_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27356_ clknet_leaf_47_clock _00385_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[29\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15370_ _11287_ VGND VGND VPWR VPWR _11365_ sky130_fd_sc_hd__clkbuf_4
X_24568_ net1170 execute.io_target_pc\[6\] _08462_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26307_ _09438_ _09446_ VGND VGND VPWR VPWR _09486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14321_ _10418_ VGND VGND VPWR VPWR _10444_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23519_ net2786 _07889_ _07900_ _07893_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27287_ clknet_leaf_8_clock _00316_ VGND VGND VPWR VPWR decode.regfile.registers_31\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24499_ _08430_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29026_ clknet_leaf_134_clock _02039_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_17040_ _12712_ decode.regfile.registers_24\[6\] _12997_ _12998_ _11025_ VGND VGND
+ VPWR VPWR _12999_ sky130_fd_sc_hd__o2111a_1
X_14252_ net1367 _10403_ _10404_ _10398_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__o211a_1
X_26238_ _09445_ VGND VGND VPWR VPWR _09446_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14183_ _10107_ _10355_ VGND VGND VPWR VPWR _10364_ sky130_fd_sc_hd__nand2_1
X_26169_ _10035_ VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__buf_4
XFILLER_0_221_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18991_ _04289_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17942_ decode.regfile.registers_10\[29\] _12790_ _12792_ VGND VGND VPWR VPWR _03340_
+ sky130_fd_sc_hd__o21ai_1
X_29928_ clknet_leaf_337_clock _02941_ VGND VGND VPWR VPWR decode.regfile.registers_21\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17873_ _12729_ _03270_ _03272_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__a21oi_1
X_29859_ clknet_leaf_307_clock _02872_ VGND VGND VPWR VPWR decode.regfile.registers_19\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16824_ _12612_ _12785_ _12786_ VGND VGND VPWR VPWR _12787_ sky130_fd_sc_hd__o21a_1
X_19612_ _04891_ _04892_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19543_ _04408_ _03929_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_176_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16755_ _12578_ VGND VGND VPWR VPWR _12719_ sky130_fd_sc_hd__clkbuf_4
Xmax_cap2 _04495_ VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_1
XFILLER_0_215_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13967_ _10142_ _10198_ VGND VGND VPWR VPWR _10238_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15706_ decode.regfile.registers_8\[10\] _11046_ _11175_ VGND VGND VPWR VPWR _11693_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19474_ net271 _04757_ _04758_ _04759_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__a31o_1
XFILLER_0_186_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16686_ _11016_ _10602_ _12508_ _12501_ VGND VGND VPWR VPWR _12651_ sky130_fd_sc_hd__or4_1
X_13898_ _10198_ VGND VGND VPWR VPWR _10199_ sky130_fd_sc_hd__clkbuf_4
XINSDIODE1_300 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_311 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_322 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18425_ _03716_ _03717_ _03720_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__nand4_4
X_15637_ _11382_ decode.regfile.registers_10\[8\] _11364_ _11625_ VGND VGND VPWR VPWR
+ _11626_ sky130_fd_sc_hd__o211a_1
XINSDIODE1_333 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_344 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_355 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_366 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_229_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_377 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18356_ _03644_ _03645_ _03649_ _03654_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__nand4_4
XFILLER_0_174_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15568_ decode.regfile.registers_20\[6\] _11102_ _11327_ _11558_ VGND VGND VPWR VPWR
+ _11559_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_352_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_352_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17307_ _13099_ _12768_ _13182_ decode.regfile.registers_29\[12\] _13259_ VGND VGND
+ VPWR VPWR _13260_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14519_ _10550_ _10554_ _10559_ _10563_ VGND VGND VPWR VPWR _10564_ sky130_fd_sc_hd__o22ai_4
X_18287_ _03608_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_25_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15499_ _11344_ net429 _11444_ _11491_ _11249_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__o221a_1
XFILLER_0_182_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17238_ decode.regfile.registers_1\[11\] _12778_ _12830_ _13191_ VGND VGND VPWR VPWR
+ _13192_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold903 fetch.bht.bhtTable_target_pc\[4\]\[19\] VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold914 fetch.bht.bhtTable_target_pc\[8\]\[0\] VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ decode.regfile.registers_20\[9\] _12771_ _13123_ _13124_ _12538_ VGND VGND
+ VPWR VPWR _13125_ sky130_fd_sc_hd__a221o_1
Xhold925 fetch.bht.bhtTable_tag\[10\]\[1\] VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold936 fetch.bht.bhtTable_tag\[2\]\[13\] VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold947 fetch.bht.bhtTable_target_pc\[4\]\[2\] VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold958 fetch.bht.bhtTable_tag\[12\]\[0\] VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__dlygate4sd3_1
X_20180_ decode.id_ex_imm_reg\[26\] decode.id_ex_pc_reg\[26\] VGND VGND VPWR VPWR
+ _05381_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold969 fetch.bht.bhtTable_tag\[10\]\[0\] VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2304 execute.csr_write_data_out_reg\[20\] VGND VGND VPWR VPWR net2531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2315 _08737_ VGND VGND VPWR VPWR net2542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2326 decode.regfile.registers_6\[19\] VGND VGND VPWR VPWR net2553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2337 fetch.btb.btbTable\[12\]\[1\] VGND VGND VPWR VPWR net2564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1603 fetch.bht.bhtTable_target_pc\[7\]\[4\] VGND VGND VPWR VPWR net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2348 csr._csr_read_data_T_8\[27\] VGND VGND VPWR VPWR net2575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1614 fetch.bht.bhtTable_tag\[15\]\[25\] VGND VGND VPWR VPWR net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2359 decode.regfile.registers_9\[23\] VGND VGND VPWR VPWR net2586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1625 fetch.bht.bhtTable_target_pc\[11\]\[17\] VGND VGND VPWR VPWR net1852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1636 decode.regfile.registers_4\[31\] VGND VGND VPWR VPWR net1863 sky130_fd_sc_hd__dlygate4sd3_1
X_23870_ execute.io_target_pc\[25\] VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1647 decode.regfile.registers_4\[15\] VGND VGND VPWR VPWR net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1658 fetch.bht.bhtTable_tag\[15\]\[19\] VGND VGND VPWR VPWR net1885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1669 fetch.bht.bhtTable_tag\[7\]\[4\] VGND VGND VPWR VPWR net1896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22821_ net1291 _10772_ _07297_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_305_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_305_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25540_ net2163 _09024_ _09031_ _09017_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22752_ _06126_ net1239 _07265_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21703_ csr.minstret\[25\] csr.minstret\[26\] _06392_ VGND VGND VPWR VPWR _06405_
+ sky130_fd_sc_hd__and3_1
X_22683_ csr._mcycle_T_2\[17\] _07223_ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__or2_1
X_25471_ net2191 _08979_ _08989_ _08991_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__o211a_1
X_27210_ clknet_leaf_363_clock _00239_ VGND VGND VPWR VPWR decode.regfile.registers_28\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_24422_ _08049_ net1843 _08389_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21634_ net606 _06350_ _06351_ _06352_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_133_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28190_ clknet_leaf_112_clock _01212_ VGND VGND VPWR VPWR csr.io_mret_vector\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27141_ clknet_leaf_359_clock _00170_ VGND VGND VPWR VPWR decode.regfile.registers_26\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_21565_ _06136_ net1487 _06295_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__mux2_1
X_24353_ net1141 execute.io_target_pc\[0\] _06141_ VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_211_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_211_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_209_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23304_ net222 _07706_ _07707_ _07733_ _07705_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__o311a_1
X_20516_ csr.meie _05517_ _05527_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24284_ _08317_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__clkbuf_1
X_27072_ clknet_leaf_347_clock _00101_ VGND VGND VPWR VPWR decode.regfile.registers_24\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_21496_ _06265_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23235_ _07066_ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26023_ net2321 _09300_ _09309_ _09305_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20447_ _05539_ _05522_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23166_ fetch.bht.bhtTable_target_pc\[0\]\[16\] fetch.bht.bhtTable_target_pc\[1\]\[16\]
+ fetch.bht.bhtTable_target_pc\[2\]\[16\] fetch.bht.bhtTable_target_pc\[3\]\[16\]
+ _07439_ _07112_ VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20378_ _05540_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22117_ fetch.bht.bhtTable_tag\[12\]\[3\] fetch.bht.bhtTable_tag\[13\]\[3\] _06644_
+ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__mux2_1
X_27974_ clknet_leaf_196_clock _00996_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_23097_ csr._csr_read_data_T_8\[12\] _06039_ csr.io_mret_vector\[12\] _06463_ VGND
+ VGND VPWR VPWR _07538_ sky130_fd_sc_hd__a22o_1
X_29713_ clknet_leaf_283_clock _02726_ VGND VGND VPWR VPWR decode.regfile.registers_14\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_22048_ _06615_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__clkbuf_8
X_26925_ _09969_ _09840_ VGND VGND VPWR VPWR _09843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_162_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29644_ clknet_leaf_277_clock _02657_ VGND VGND VPWR VPWR decode.regfile.registers_12\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14870_ _10575_ VGND VGND VPWR VPWR _10912_ sky130_fd_sc_hd__clkbuf_2
X_26856_ _09383_ _09796_ VGND VGND VPWR VPWR _09803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_215_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13821_ _10152_ VGND VGND VPWR VPWR _10154_ sky130_fd_sc_hd__buf_2
X_25807_ decode.regfile.registers_6\[21\] _09183_ _09185_ _09182_ VGND VGND VPWR VPWR
+ _02468_ sky130_fd_sc_hd__o211a_1
X_29575_ clknet_leaf_273_clock _02588_ VGND VGND VPWR VPWR decode.regfile.registers_10\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_26787_ _09751_ VGND VGND VPWR VPWR _09763_ sky130_fd_sc_hd__clkbuf_4
X_23999_ net1619 execute.io_target_pc\[20\] _08164_ VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_218_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28526_ clknet_leaf_214_clock _01539_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16540_ _12504_ VGND VGND VPWR VPWR _12505_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13752_ memory.io_wb_reg_pc\[22\] _09946_ _09947_ _10094_ VGND VGND VPWR VPWR _10095_
+ sky130_fd_sc_hd__a31o_1
X_25738_ net2003 _09139_ _09145_ _09142_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28457_ clknet_leaf_149_clock _01470_ VGND VGND VPWR VPWR decode.io_id_pc\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16471_ decode.regfile.registers_18\[30\] _11269_ _12436_ _12437_ _11271_ VGND VGND
+ VPWR VPWR _12438_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13683_ _10036_ _10016_ VGND VGND VPWR VPWR _10037_ sky130_fd_sc_hd__nand2_1
X_25669_ _08968_ _09067_ VGND VGND VPWR VPWR _09105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_214_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18210_ _12494_ _03518_ _03521_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__or3b_1
XFILLER_0_156_948 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27408_ clknet_leaf_10_clock _00437_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[17\]
+ sky130_fd_sc_hd__dfxtp_4
X_15422_ decode.regfile.registers_4\[3\] _11410_ _11097_ _10648_ _11415_ VGND VGND
+ VPWR VPWR _11416_ sky130_fd_sc_hd__o221a_1
X_19190_ _04274_ _04054_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__nor2_1
X_28388_ clknet_leaf_145_clock _01401_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18141_ _03499_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27339_ clknet_leaf_43_clock _00368_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_15353_ _11338_ VGND VGND VPWR VPWR _11348_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14304_ _10031_ _10431_ VGND VGND VPWR VPWR _10435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18072_ _03459_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15284_ _11192_ VGND VGND VPWR VPWR _11280_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_130_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29009_ clknet_leaf_103_clock _02022_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_169_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire174 net175 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
X_17023_ decode.regfile.registers_13\[6\] _12927_ _12588_ VGND VGND VPWR VPWR _12982_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_150_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire185 _00507_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
X_14235_ net1233 _10390_ _10394_ _10385_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_169_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14166_ _10069_ _10342_ VGND VGND VPWR VPWR _10354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18974_ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__clkbuf_4
X_14097_ net2559 _10302_ _10314_ _10304_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17925_ decode.regfile.registers_18\[28\] _10924_ _12568_ _12524_ _11008_ VGND VGND
+ VPWR VPWR _03324_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_128_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17856_ _02986_ decode.regfile.registers_26\[26\] _13002_ _13484_ _02987_ VGND VGND
+ VPWR VPWR _03257_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_179_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1083 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16807_ _12524_ _12551_ _12523_ VGND VGND VPWR VPWR _12770_ sky130_fd_sc_hd__and3_1
X_17787_ decode.regfile.registers_4\[25\] decode.regfile.registers_5\[25\] _10616_
+ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14999_ _11011_ _11004_ _11006_ _11007_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19526_ _04408_ _04508_ _04807_ _04415_ _04809_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__o311a_1
XFILLER_0_53_1212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16738_ net2489 _12491_ _12520_ net505 _12702_ VGND VGND VPWR VPWR _12703_ sky130_fd_sc_hd__o32a_1
XFILLER_0_159_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19457_ _04334_ _04152_ _04160_ _04164_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16669_ _12633_ VGND VGND VPWR VPWR _12634_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_291_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_291_clock
+ sky130_fd_sc_hd__clkbuf_8
XINSDIODE1_130 _11217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_141 _12412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_152 _12636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18408_ _03706_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__buf_4
XFILLER_0_173_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19388_ _04509_ _04369_ _04515_ _04633_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_163 decode.id_ex_rs1_data_reg\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_174 decode.id_ex_rs2_data_reg\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_185 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_196 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18339_ _03637_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_98_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21350_ _10556_ _10557_ _09885_ _09916_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__nand4_4
XFILLER_0_112_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20301_ _05340_ _05473_ _05411_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21281_ _10771_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__buf_2
XFILLER_0_163_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold700 decode.regfile.registers_26\[2\] VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 fetch.bht.bhtTable_target_pc\[8\]\[15\] VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23020_ _07391_ _07392_ _07464_ _07465_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold722 csr._mcycle_T_3\[57\] VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 fetch.bht.bhtTable_tag\[3\]\[2\] VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__dlygate4sd3_1
X_20232_ _05422_ _05423_ _05245_ _05411_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold744 fetch.bht.bhtTable_target_pc\[11\]\[13\] VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 decode.regfile.registers_28\[4\] VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold766 decode.regfile.registers_20\[2\] VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold777 fetch.bht.bhtTable_tag\[12\]\[15\] VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 fetch.bht.bhtTable_target_pc\[5\]\[4\] VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__dlygate4sd3_1
X_20163_ _05364_ _05366_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__xor2_1
Xhold799 fetch.bht.bhtTable_tag\[12\]\[16\] VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2101 decode.regfile.registers_4\[23\] VGND VGND VPWR VPWR net2328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2112 decode.regfile.registers_11\[10\] VGND VGND VPWR VPWR net2339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_200_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2123 decode.regfile.registers_8\[27\] VGND VGND VPWR VPWR net2350 sky130_fd_sc_hd__dlygate4sd3_1
X_20094_ _00561_ _05228_ _05307_ _05231_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__o22a_1
X_24971_ net2561 _08693_ _06318_ VGND VGND VPWR VPWR _08694_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_196_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2134 decode.regfile.registers_3\[19\] VGND VGND VPWR VPWR net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1400 fetch.bht.bhtTable_tag\[0\]\[9\] VGND VGND VPWR VPWR net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2145 decode.regfile.registers_20\[26\] VGND VGND VPWR VPWR net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2156 fetch.bht.bhtTable_tag\[15\]\[16\] VGND VGND VPWR VPWR net2383 sky130_fd_sc_hd__dlygate4sd3_1
X_26710_ _09387_ _09710_ VGND VGND VPWR VPWR _09719_ sky130_fd_sc_hd__nand2_1
Xhold1411 decode.regfile.registers_18\[2\] VGND VGND VPWR VPWR net1638 sky130_fd_sc_hd__dlygate4sd3_1
X_23922_ _08131_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__clkbuf_1
Xhold1422 fetch.bht.bhtTable_tag\[5\]\[1\] VGND VGND VPWR VPWR net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2167 decode.regfile.registers_3\[20\] VGND VGND VPWR VPWR net2394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 fetch.bht.bhtTable_target_pc\[0\]\[4\] VGND VGND VPWR VPWR net1660 sky130_fd_sc_hd__dlygate4sd3_1
X_27690_ clknet_leaf_25_clock _00719_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_244_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_244_clock
+ sky130_fd_sc_hd__clkbuf_8
Xhold2178 decode.regfile.registers_19\[28\] VGND VGND VPWR VPWR net2405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1444 fetch.bht.bhtTable_tag\[7\]\[5\] VGND VGND VPWR VPWR net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2189 decode.regfile.registers_25\[21\] VGND VGND VPWR VPWR net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 fetch.bht.bhtTable_target_pc\[10\]\[8\] VGND VGND VPWR VPWR net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1466 fetch.bht.bhtTable_tag\[13\]\[2\] VGND VGND VPWR VPWR net1693 sky130_fd_sc_hd__dlygate4sd3_1
X_26641_ _09664_ VGND VGND VPWR VPWR _09679_ sky130_fd_sc_hd__clkbuf_4
Xhold1477 fetch.bht.bhtTable_target_pc\[8\]\[6\] VGND VGND VPWR VPWR net1704 sky130_fd_sc_hd__dlygate4sd3_1
X_23853_ _08089_ net1892 _08079_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1488 fetch.bht.bhtTable_target_pc\[4\]\[8\] VGND VGND VPWR VPWR net1715 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 fetch.bht.bhtTable_tag\[5\]\[13\] VGND VGND VPWR VPWR net1726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22804_ _07285_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_169_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29360_ clknet_leaf_227_clock _02373_ VGND VGND VPWR VPWR decode.regfile.registers_3\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_26572_ net669 _09636_ _09639_ _09635_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__o211a_1
X_23784_ _08044_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20996_ _05981_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__clkbuf_1
X_28311_ clknet_leaf_165_clock _01324_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25523_ net2528 _08980_ _09020_ _09017_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22735_ _06109_ net1120 _09903_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__mux2_1
X_29291_ clknet_leaf_242_clock _02304_ VGND VGND VPWR VPWR decode.regfile.registers_1\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_259_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_259_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28242_ clknet_leaf_77_clock _01264_ VGND VGND VPWR VPWR csr._minstret_T_3\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_25454_ net2162 _08979_ _08981_ _08972_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__o211a_1
X_22666_ net2796 _07210_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24405_ net832 execute.io_target_pc\[25\] _09911_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21617_ _05613_ csr.minstret\[5\] _06338_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__and3_1
X_28173_ clknet_leaf_53_clock _01195_ VGND VGND VPWR VPWR csr.io_mret_vector\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25385_ _10041_ VGND VGND VPWR VPWR _08933_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_180_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22597_ csr._minstret_T_3\[47\] csr._minstret_T_3\[46\] _07172_ _06422_ VGND VGND
+ VPWR VPWR _07175_ sky130_fd_sc_hd__a31o_1
XFILLER_0_146_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27124_ clknet_leaf_329_clock _00153_ VGND VGND VPWR VPWR decode.regfile.registers_26\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_24336_ _08344_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21548_ _06119_ net2056 _06284_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27055_ clknet_leaf_330_clock _00084_ VGND VGND VPWR VPWR decode.regfile.registers_24\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_24267_ _08095_ net1971 _08300_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__mux2_1
X_21479_ _06256_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14020_ _10081_ _10268_ VGND VGND VPWR VPWR _10270_ sky130_fd_sc_hd__nand2_1
X_26006_ _09285_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__clkbuf_4
X_23218_ net76 _06887_ _07613_ net224 VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24198_ _08273_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23149_ _06025_ _07573_ _03546_ _07587_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_164_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27957_ clknet_leaf_195_clock _00979_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_15971_ decode.regfile.registers_5\[17\] _10636_ _11138_ VGND VGND VPWR VPWR _11951_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_160_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17710_ decode.regfile.registers_15\[23\] _10612_ _10619_ _12589_ _13031_ VGND VGND
+ VPWR VPWR _03114_ sky130_fd_sc_hd__a41o_1
X_14922_ _10579_ _10578_ VGND VGND VPWR VPWR _10951_ sky130_fd_sc_hd__or2_2
X_26908_ _09436_ _09794_ VGND VGND VPWR VPWR _09832_ sky130_fd_sc_hd__nand2_1
X_18690_ _03988_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__buf_4
X_27888_ clknet_leaf_22_clock _00917_ VGND VGND VPWR VPWR csr._mcycle_T_2\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17641_ decode.regfile.registers_10\[21\] _12654_ _03034_ _03046_ _12878_ VGND VGND
+ VPWR VPWR _03047_ sky130_fd_sc_hd__o221ai_4
X_14853_ _10894_ _10895_ VGND VGND VPWR VPWR _10896_ sky130_fd_sc_hd__nand2_1
X_29627_ clknet_leaf_271_clock _02640_ VGND VGND VPWR VPWR decode.regfile.registers_12\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_26839_ _09443_ _09751_ VGND VGND VPWR VPWR _09792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_216_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13804_ _10060_ _10138_ _09947_ memory.io_wb_aluresult\[30\] VGND VGND VPWR VPWR
+ _10139_ sky130_fd_sc_hd__o22a_1
X_17572_ decode.regfile.registers_21\[19\] _12682_ _12909_ VGND VGND VPWR VPWR _02980_
+ sky130_fd_sc_hd__o21a_1
X_29558_ clknet_leaf_266_clock _02571_ VGND VGND VPWR VPWR decode.regfile.registers_9\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14784_ _10684_ csr.io_mem_pc\[30\] _10826_ VGND VGND VPWR VPWR _10827_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_63_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_212_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19311_ _04435_ _04317_ _04294_ _04603_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__a211o_1
X_28509_ clknet_leaf_215_clock _01522_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16523_ _10598_ decode.immGen._imm_T_24\[17\] VGND VGND VPWR VPWR _12488_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_158_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13735_ net201 VGND VGND VPWR VPWR _10081_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29489_ clknet_leaf_264_clock _02502_ VGND VGND VPWR VPWR decode.regfile.registers_7\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19242_ _04243_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__clkbuf_4
X_16454_ _10647_ _11097_ decode.regfile.registers_5\[30\] VGND VGND VPWR VPWR _12421_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_156_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13666_ _10012_ _10021_ memory.io_wb_readdata\[9\] VGND VGND VPWR VPWR _10022_ sky130_fd_sc_hd__and3b_1
XFILLER_0_155_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15405_ _11397_ _11399_ VGND VGND VPWR VPWR _11400_ sky130_fd_sc_hd__nand2_1
X_19173_ _04363_ _04367_ _04246_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16385_ decode.regfile.registers_2\[28\] _11296_ VGND VGND VPWR VPWR _12354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ memory.io_wb_memtoreg\[1\] memory.io_wb_memtoreg\[0\] VGND VGND VPWR VPWR
+ _09961_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18124_ _03482_ _03480_ _03487_ decode.io_id_pc\[18\] VGND VGND VPWR VPWR _03490_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_143_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15336_ _11060_ _10977_ _11049_ _11072_ VGND VGND VPWR VPWR _11332_ sky130_fd_sc_hd__or4b_1
XFILLER_0_186_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18055_ _03448_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15267_ _10956_ VGND VGND VPWR VPWR _11263_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_93_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2 _00931_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17006_ _12492_ VGND VGND VPWR VPWR _12965_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_188_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14218_ _10290_ VGND VGND VPWR VPWR _10385_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15198_ _10648_ _10630_ _11044_ _11051_ VGND VGND VPWR VPWR _11195_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14149_ _10025_ _10342_ VGND VGND VPWR VPWR _10345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_892 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18957_ _03986_ _03985_ _03984_ _03987_ _04205_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__a311o_1
XFILLER_0_67_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ decode.regfile.registers_10\[28\] _10617_ _12776_ _10611_ _12604_ VGND VGND
+ VPWR VPWR _03307_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_94_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18888_ net284 _04103_ _04185_ _04186_ _04095_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_206_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17839_ decode.regfile.registers_10\[26\] _12654_ _12878_ VGND VGND VPWR VPWR _03240_
+ sky130_fd_sc_hd__o21ai_1
Xrebuffer14 net253 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer25 _03757_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_1
Xrebuffer36 net360 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_1
XFILLER_0_178_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20850_ net112 _05891_ _05899_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__and3_1
Xrebuffer47 _04106_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer58 net283 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__buf_1
XFILLER_0_117_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer69 net293 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_1
X_19509_ _04537_ _04792_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20781_ net99 _05859_ _05860_ _05862_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22520_ _07113_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22451_ _06645_ fetch.btb.btbTable\[3\]\[1\] fetch.bht.bhtTable_valid\[3\] _07045_
+ _06631_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_147_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer104 _09929_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_4
X_21402_ _06214_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer115 net341 VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22382_ _06928_ _06944_ _06965_ _06976_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__or4_1
X_25170_ _09880_ _09883_ _08813_ VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__or3_1
XFILLER_0_228_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24121_ net875 execute.io_target_pc\[15\] _08232_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__mux2_1
X_21333_ net1068 _10772_ _06168_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21264_ _06135_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__clkbuf_1
X_24052_ _07990_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold530 decode.regfile.registers_11\[5\] VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold541 decode.regfile.registers_25\[13\] VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 decode.regfile.registers_28\[25\] VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__dlygate4sd3_1
X_23003_ _07391_ _07392_ _07446_ _07449_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__a31o_1
X_20215_ _05410_ _05267_ _05200_ _05247_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__a22oi_2
Xhold563 csr._mcycle_T_3\[43\] VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28860_ clknet_leaf_183_clock _01873_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold574 decode.regfile.registers_31\[2\] VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd3_1
X_21195_ _06086_ _06082_ net1918 VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__and3_1
Xhold585 fetch.bht.bhtTable_tag\[2\]\[23\] VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold596 fetch.bht.bhtTable_tag\[2\]\[9\] VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27811_ clknet_leaf_35_clock _00840_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20146_ _05350_ _05351_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28791_ clknet_leaf_125_clock _01804_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_183_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_183_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_202_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27742_ clknet_leaf_37_clock _00771_ VGND VGND VPWR VPWR decode.io_wb_regwrite sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20077_ _05283_ _05292_ _05288_ _05289_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__a211o_1
X_24954_ csr._mcycle_T_3\[53\] _08682_ _06318_ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_198_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1230 fetch.bht.bhtTable_target_pc\[3\]\[9\] VGND VGND VPWR VPWR net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 fetch.bht.bhtTable_target_pc\[14\]\[11\] VGND VGND VPWR VPWR net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 fetch.bht.bhtTable_target_pc\[10\]\[27\] VGND VGND VPWR VPWR net1479 sky130_fd_sc_hd__dlygate4sd3_1
X_23905_ _08122_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27673_ clknet_leaf_28_clock _00702_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_24885_ _08634_ VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__clkbuf_2
Xhold1263 decode.regfile.registers_12\[31\] VGND VGND VPWR VPWR net1490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1274 fetch.bht.bhtTable_target_pc\[2\]\[2\] VGND VGND VPWR VPWR net1501 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 csr._minstret_T_3\[52\] VGND VGND VPWR VPWR net1512 sky130_fd_sc_hd__dlygate4sd3_1
X_29412_ clknet_leaf_257_clock _02425_ VGND VGND VPWR VPWR decode.regfile.registers_5\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1296 fetch.bht.bhtTable_target_pc\[13\]\[23\] VGND VGND VPWR VPWR net1523 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26624_ net2085 _09665_ _09669_ _09660_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__o211a_1
X_23836_ execute.io_target_pc\[14\] VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__buf_2
XFILLER_0_196_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_198_clock clknet_5_27__leaf_clock VGND VGND VPWR VPWR clknet_leaf_198_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29343_ clknet_leaf_230_clock _02356_ VGND VGND VPWR VPWR decode.regfile.registers_3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26555_ net2440 _09622_ _09629_ _09619_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23767_ _08035_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20979_ execute.io_reg_pc\[15\] _05965_ _05961_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13520_ net684 _09898_ VGND VGND VPWR VPWR _09899_ sky130_fd_sc_hd__or2_1
X_25506_ net2727 _09008_ _09011_ _09004_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__o211a_1
X_29274_ clknet_leaf_243_clock _02287_ VGND VGND VPWR VPWR decode.regfile.registers_1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_22718_ _10943_ _10941_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26486_ _09389_ _09589_ VGND VGND VPWR VPWR _09590_ sky130_fd_sc_hd__nand2_1
X_23698_ _07999_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_121_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_121_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28225_ clknet_leaf_87_clock net1958 VGND VGND VPWR VPWR csr.mscratch\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25437_ _08968_ _08905_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22649_ _07209_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28156_ clknet_leaf_66_clock _01178_ VGND VGND VPWR VPWR csr.mtie sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16170_ decode.regfile.registers_7\[22\] _11465_ _11466_ decode.regfile.registers_6\[22\]
+ _11166_ VGND VGND VPWR VPWR _12145_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25368_ _08920_ _08907_ VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27107_ clknet_leaf_357_clock _00136_ VGND VGND VPWR VPWR decode.regfile.registers_25\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_15121_ _11117_ VGND VGND VPWR VPWR _11118_ sky130_fd_sc_hd__clkbuf_4
X_24319_ _08081_ net1325 _08334_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28087_ clknet_leaf_199_clock _01109_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_136_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_136_clock
+ sky130_fd_sc_hd__clkbuf_8
X_25299_ _10018_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__buf_2
X_27038_ clknet_leaf_345_clock _00067_ VGND VGND VPWR VPWR decode.regfile.registers_23\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15052_ _11048_ VGND VGND VPWR VPWR _11049_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14003_ net731 _10258_ _10260_ _10249_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19860_ _05124_ _05125_ _05130_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_102_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput72 net72 VGND VGND VPWR VPWR io_fetch_address[14] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18811_ execute.io_reg_pc\[12\] _03662_ _03663_ net103 _04109_ VGND VGND VPWR VPWR
+ _04110_ sky130_fd_sc_hd__o221a_1
Xoutput83 net83 VGND VGND VPWR VPWR io_fetch_address[24] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput94 net94 VGND VGND VPWR VPWR io_fetch_address[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19791_ _04225_ _04424_ _05060_ _05063_ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__o32a_1
X_28989_ clknet_leaf_180_clock _02002_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15954_ decode.regfile.registers_21\[16\] _11061_ _11100_ _11229_ _11934_ VGND VGND
+ VPWR VPWR _11935_ sky130_fd_sc_hd__o311a_1
X_18742_ execute.io_reg_pc\[5\] _03776_ _03664_ net127 _04040_ VGND VGND VPWR VPWR
+ _04041_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14905_ _10595_ VGND VGND VPWR VPWR _10938_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_121_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18673_ _03967_ net241 net305 net359 decode.id_ex_immsrc_reg VGND VGND VPWR VPWR
+ _03972_ sky130_fd_sc_hd__a41o_4
X_15885_ _11260_ _11865_ _11866_ _11867_ VGND VGND VPWR VPWR _11868_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14836_ _10878_ _10812_ net268 csr.io_mem_pc\[12\] VGND VGND VPWR VPWR _10879_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_118_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17624_ _02997_ _13262_ _13182_ decode.regfile.registers_29\[20\] _03030_ VGND VGND
+ VPWR VPWR _03031_ sky130_fd_sc_hd__o221a_1
XFILLER_0_176_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17555_ _12838_ _02961_ _02962_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__o21ai_2
X_14767_ csr.io_mem_pc\[13\] _10763_ VGND VGND VPWR VPWR _10810_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16506_ _10640_ _11125_ _11104_ decode.regfile.registers_17\[31\] _11126_ VGND VGND
+ VPWR VPWR _12472_ sky130_fd_sc_hd__o32a_1
XFILLER_0_168_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13718_ _10012_ _10021_ memory.io_wb_reg_pc\[17\] VGND VGND VPWR VPWR _10066_ sky130_fd_sc_hd__or3b_1
X_17486_ decode.regfile.registers_12\[17\] _12542_ _12772_ _12658_ _13433_ VGND VGND
+ VPWR VPWR _13434_ sky130_fd_sc_hd__o311a_1
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14698_ _10731_ execute.io_target_pc\[7\] VGND VGND VPWR VPWR _10741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19225_ _04518_ _04039_ _04519_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__and3_1
X_16437_ decode.regfile.registers_18\[29\] _10956_ _11114_ _10989_ _10977_ VGND VGND
+ VPWR VPWR _12405_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13649_ memory.csr_read_data_out_reg\[7\] _09989_ _10002_ _10006_ VGND VGND VPWR
+ VPWR _10007_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_171_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19156_ _04024_ _04451_ _04452_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16368_ decode.regfile.registers_23\[27\] _11262_ _12312_ _12337_ _11335_ VGND VGND
+ VPWR VPWR _12338_ sky130_fd_sc_hd__o221a_1
XFILLER_0_186_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18107_ _10909_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__buf_2
XFILLER_0_26_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15319_ _10655_ _11313_ _11314_ _10660_ VGND VGND VPWR VPWR _11315_ sky130_fd_sc_hd__or4b_4
X_19087_ _04316_ _04374_ _04384_ _04243_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__a22o_1
X_16299_ _11756_ decode.regfile.registers_28\[25\] _11871_ _11681_ _11448_ VGND VGND
+ VPWR VPWR _12271_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_83_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18038_ decode.regfile.registers_20\[31\] _12771_ _03432_ _03433_ _12538_ VGND VGND
+ VPWR VPWR _03434_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20000_ _05226_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19989_ _05220_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1034 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21951_ net512 _06572_ _06576_ _10546_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ _05930_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__clkbuf_1
X_24670_ _08518_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21882_ net881 _06521_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23621_ _06151_ net2032 _07952_ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20833_ net103 _05891_ _05887_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26340_ _09396_ _09502_ VGND VGND VPWR VPWR _09506_ sky130_fd_sc_hd__nand2_1
X_23552_ net222 _07917_ _07920_ _05805_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_194_Right_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20764_ _03452_ _05425_ csr.io_csr_address\[9\] VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__and3b_1
XFILLER_0_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22503_ _06740_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__buf_4
XFILLER_0_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26271_ _09402_ _09459_ VGND VGND VPWR VPWR _09466_ sky130_fd_sc_hd__nand2_1
X_23483_ net19 _07875_ _07880_ _07879_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__o211a_1
X_20695_ decode.id_ex_funct3_reg\[0\] decode.id_ex_funct3_reg\[1\] _05056_ _10575_
+ _10909_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28010_ clknet_leaf_187_clock _01032_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25222_ _08840_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22434_ fetch.bht.bhtTable_tag\[10\]\[12\] fetch.bht.bhtTable_tag\[11\]\[12\] _06691_
+ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_53_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_53_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25153_ net406 _08804_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22365_ fetch.bht.bhtTable_tag\[12\]\[2\] fetch.bht.bhtTable_tag\[13\]\[2\] fetch.bht.bhtTable_tag\[14\]\[2\]
+ fetch.bht.bhtTable_tag\[15\]\[2\] net275 _06620_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24104_ net813 execute.io_target_pc\[7\] _08221_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__mux2_1
X_21316_ _06156_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__buf_4
X_25084_ _06101_ net1736 _08596_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__mux2_1
X_22296_ _06864_ _06888_ _06889_ _06890_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_103_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_68_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_68_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28912_ clknet_leaf_105_clock _01925_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_21247_ _10803_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__buf_2
X_24035_ _08189_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold360 decode.regfile.registers_12\[3\] VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 decode.regfile.registers_12\[9\] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__dlygate4sd3_1
X_29892_ clknet_leaf_302_clock _02905_ VGND VGND VPWR VPWR decode.regfile.registers_20\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold382 decode.regfile.registers_12\[2\] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 csr._mcycle_T_3\[33\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__dlygate4sd3_1
X_28843_ clknet_leaf_91_clock _01856_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_21178_ _06074_ _06082_ net1811 VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_225_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20129_ _05334_ _05337_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__xnor2_1
X_28774_ clknet_leaf_97_clock _01787_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_196_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25986_ _08982_ _09287_ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_221_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_221_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27725_ clknet_leaf_23_clock _00754_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_24937_ net2314 _08670_ _08671_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__o21ba_1
Xhold1060 fetch.bht.bhtTable_tag\[7\]\[9\] VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1071 decode.regfile.registers_9\[13\] VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1082 fetch.bht.bhtTable_target_pc\[6\]\[26\] VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__dlygate4sd3_1
X_27656_ clknet_leaf_65_clock _00685_ VGND VGND VPWR VPWR execute.io_wfi_out sky130_fd_sc_hd__dfxtp_1
X_15670_ _11375_ _11655_ _11656_ _11657_ _11138_ VGND VGND VPWR VPWR _11658_ sky130_fd_sc_hd__a32o_1
X_24868_ _06147_ net2303 _08388_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1093 fetch.bht.bhtTable_tag\[9\]\[14\] VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26607_ net2217 _09649_ _09658_ _09648_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__o211a_1
X_14621_ _10656_ _10658_ _10661_ _10663_ VGND VGND VPWR VPWR _10664_ sky130_fd_sc_hd__a2bb2o_1
X_23819_ _08066_ net1469 _08058_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27587_ clknet_leaf_150_clock _00616_ VGND VGND VPWR VPWR csr.io_mem_pc\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _08586_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_155_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29326_ clknet_leaf_226_clock _02339_ VGND VGND VPWR VPWR decode.regfile.registers_2\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17340_ _13250_ decode.regfile.registers_24\[13\] _13170_ _13083_ _12862_ VGND VGND
+ VPWR VPWR _13292_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_200_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26538_ _09566_ VGND VGND VPWR VPWR _09619_ sky130_fd_sc_hd__buf_2
X_14552_ _10594_ VGND VGND VPWR VPWR _10595_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13503_ fetch.bht.bhtTable_tag_MPORT_en VGND VGND VPWR VPWR _09885_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29257_ clknet_leaf_233_clock _02270_ VGND VGND VPWR VPWR decode.regfile.registers_0\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_17271_ decode.regfile.registers_12\[12\] _12551_ _12583_ _12775_ VGND VGND VPWR
+ VPWR _13224_ sky130_fd_sc_hd__a31o_1
X_26469_ net2180 _09578_ _09580_ _09567_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__o211a_1
X_14483_ net436 _10533_ _10537_ _10535_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19010_ _09949_ _04046_ _03985_ _03984_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__o211ai_1
X_28208_ clknet_leaf_62_clock net1591 VGND VGND VPWR VPWR csr.mscratch\[10\] sky130_fd_sc_hd__dfxtp_1
X_16222_ decode.regfile.registers_23\[23\] _11087_ _12171_ _12195_ VGND VGND VPWR
+ VPWR _12196_ sky130_fd_sc_hd__o22a_1
X_29188_ clknet_leaf_240_clock _02201_ VGND VGND VPWR VPWR fetch.btb.btbTable\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28139_ clknet_leaf_203_clock _01161_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16153_ _11251_ _11259_ decode.regfile.registers_27\[21\] _12099_ _12128_ VGND VGND
+ VPWR VPWR _12129_ sky130_fd_sc_hd__o32a_1
Xrebuffer5 net205 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15104_ _10625_ _11092_ _11048_ _10652_ VGND VGND VPWR VPWR _11101_ sky130_fd_sc_hd__and4_2
XFILLER_0_121_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16084_ _12059_ _12060_ _11369_ VGND VGND VPWR VPWR _12061_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15035_ decode.control.io_funct7\[5\] _10998_ _10969_ _11030_ VGND VGND VPWR VPWR
+ _00386_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19912_ _04325_ _05137_ _05179_ _04572_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_75_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19843_ _04805_ _04415_ _04751_ _04949_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__a31o_1
XFILLER_0_177_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19774_ _05026_ _03853_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16986_ decode.regfile.registers_12\[5\] _12745_ _12929_ _12945_ _12658_ VGND VGND
+ VPWR VPWR _12946_ sky130_fd_sc_hd__o221a_1
XFILLER_0_155_1305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18725_ _04022_ _04023_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__or2_2
XFILLER_0_218_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15937_ _11410_ _11192_ _11914_ _11917_ VGND VGND VPWR VPWR _11918_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_79_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15868_ _11849_ _11850_ VGND VGND VPWR VPWR _11851_ sky130_fd_sc_hd__nand2_1
X_18656_ net231 _03951_ decode.id_ex_rs1_data_reg\[20\] _03687_ VGND VGND VPWR VPWR
+ _03955_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_203_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14819_ _10769_ _10858_ decode.id_ex_pc_reg\[26\] VGND VGND VPWR VPWR _10862_ sky130_fd_sc_hd__o21ai_1
X_17607_ decode.regfile.registers_14\[20\] _12984_ _03000_ _03013_ _12874_ VGND VGND
+ VPWR VPWR _03014_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_47_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15799_ _11203_ _11782_ _11783_ VGND VGND VPWR VPWR _11784_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18587_ _03817_ _03885_ _03774_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17538_ _13087_ decode.regfile.registers_26\[18\] _13254_ _13484_ _13088_ VGND VGND
+ VPWR VPWR _13485_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17469_ decode.regfile.registers_20\[17\] _12525_ _12552_ _12523_ _12824_ VGND VGND
+ VPWR VPWR _13417_ sky130_fd_sc_hd__a41o_1
XFILLER_0_172_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19208_ _04311_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20480_ _05627_ csr.io_mret_vector\[6\] _05603_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19139_ _04280_ _04282_ _04289_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__o21ai_4
XPHY_EDGE_ROW_89_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22150_ _06652_ _06744_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__and2b_1
XFILLER_0_70_896 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21101_ _06040_ _06041_ _10577_ _09926_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__nor4_1
XFILLER_0_160_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22081_ fetch.bht.bhtTable_tag\[0\]\[7\] fetch.bht.bhtTable_tag\[1\]\[7\] fetch.bht.bhtTable_tag\[2\]\[7\]
+ fetch.bht.bhtTable_tag\[3\]\[7\] _06674_ _06675_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21032_ execute.csr_read_data_out_reg\[6\] _05989_ _05998_ VGND VGND VPWR VPWR _06001_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_100_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25840_ net672 _09199_ _09204_ _09194_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_214_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25771_ net1890 _09156_ _09164_ _09153_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_98_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22983_ execute.io_target_pc\[5\] _06032_ _07345_ _07418_ _07430_ VGND VGND VPWR
+ VPWR _07431_ sky130_fd_sc_hd__o311a_1
X_27510_ clknet_leaf_21_clock _00539_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dfxtp_1
X_24722_ _08545_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__clkbuf_1
X_28490_ clknet_leaf_200_clock _01503_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[15\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_21934_ csr._mcycle_T_2\[29\] _06545_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27441_ clknet_leaf_153_clock _00470_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_24653_ net1382 execute.io_target_pc\[15\] _08508_ VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21865_ _06039_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__clkbuf_4
X_23604_ _06134_ net2383 _07941_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20816_ _05883_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_1
X_27372_ clknet_leaf_9_clock _00401_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_24584_ net972 VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__clkbuf_1
X_21796_ _06460_ net590 _06396_ _06465_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29111_ clknet_leaf_18_clock _02124_ VGND VGND VPWR VPWR csr._mcycle_T_3\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26323_ _09379_ _09492_ VGND VGND VPWR VPWR _09496_ sky130_fd_sc_hd__nand2_1
X_23535_ net1384 _07903_ _07910_ _07907_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_150_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20747_ _05831_ _05813_ decode.id_ex_rs1_data_reg\[30\] _05844_ _00717_ VGND VGND
+ VPWR VPWR _00749_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_189_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_189_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29042_ clknet_leaf_101_clock _02055_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26254_ _09385_ _09448_ VGND VGND VPWR VPWR _09456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23466_ _10962_ _07862_ _07859_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__or3b_1
XFILLER_0_64_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20678_ _05798_ _05802_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__nor2_1
X_25205_ _08831_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22417_ fetch.bht.bhtTable_tag\[12\]\[1\] fetch.bht.bhtTable_tag\[13\]\[1\] _06691_
+ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26185_ _09408_ _09390_ VGND VGND VPWR VPWR _09409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23397_ net88 _06795_ _07783_ net90 VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25136_ _08796_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__clkbuf_1
X_22348_ _06641_ _06932_ _06936_ _06942_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__o31a_2
XFILLER_0_131_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25067_ csr.mcycle\[26\] csr.mcycle\[25\] _08754_ VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_148_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29944_ clknet_leaf_334_clock _02957_ VGND VGND VPWR VPWR decode.regfile.registers_21\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_22279_ fetch.bht.bhtTable_tag\[6\]\[6\] fetch.bht.bhtTable_tag\[7\]\[6\] _06700_
+ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_223_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24018_ _08180_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_180_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold190 execute.io_mem_isjump VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
X_29875_ clknet_leaf_300_clock _02888_ VGND VGND VPWR VPWR decode.regfile.registers_19\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28826_ clknet_leaf_179_clock _01839_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16840_ decode.regfile.registers_18\[2\] _12572_ _12562_ _12802_ VGND VGND VPWR VPWR
+ _12803_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_70_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16771_ _11016_ _10597_ _10935_ _10602_ VGND VGND VPWR VPWR _12735_ sky130_fd_sc_hd__or4_4
X_28757_ clknet_leaf_116_clock _01770_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_13983_ net2004 _10243_ _10248_ _10249_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__o211a_1
X_25969_ net2389 _09270_ _09278_ _09277_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15722_ decode.regfile.registers_16\[10\] _11203_ _11357_ VGND VGND VPWR VPWR _11709_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18510_ _03709_ decode.id_ex_imm_reg\[26\] _03807_ _03808_ VGND VGND VPWR VPWR _03809_
+ sky130_fd_sc_hd__a22oi_4
X_27708_ clknet_leaf_20_clock _00737_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_19490_ _04537_ _04572_ _04573_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__or3_1
X_28688_ clknet_leaf_120_clock _01701_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _11251_ _11259_ decode.regfile.registers_27\[8\] _11611_ _11641_ VGND VGND
+ VPWR VPWR _11642_ sky130_fd_sc_hd__o32a_1
XFILLER_0_34_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18441_ decode.io_wb_rd\[2\] csr.io_csr_address\[2\] VGND VGND VPWR VPWR _03740_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_201_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27639_ clknet_leaf_155_clock _00668_ VGND VGND VPWR VPWR execute.io_reg_pc\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XINSDIODE1_80 _10588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_91 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14604_ _10646_ VGND VGND VPWR VPWR _10647_ sky130_fd_sc_hd__buf_4
X_18372_ _09929_ decode.id_ex_ex_rs1_reg\[2\] VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__or2b_4
XFILLER_0_201_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15584_ decode.regfile.registers_14\[7\] _11360_ _11274_ decode.regfile.registers_15\[7\]
+ _11202_ VGND VGND VPWR VPWR _11574_ sky130_fd_sc_hd__a221o_1
XFILLER_0_205_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17323_ _12603_ _13274_ VGND VGND VPWR VPWR _13275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29309_ clknet_leaf_244_clock _02322_ VGND VGND VPWR VPWR decode.regfile.registers_2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14535_ decode.control.io_opcode\[3\] decode.control.io_opcode\[2\] decode.control.io_opcode\[1\]
+ decode.control.io_opcode\[0\] VGND VGND VPWR VPWR _10578_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_200_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17254_ _13081_ _13168_ decode.regfile.registers_23\[11\] _13041_ VGND VGND VPWR
+ VPWR _13208_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14466_ net438 _10520_ _10527_ _10522_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_137_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16205_ _11044_ decode.regfile.registers_4\[23\] _11191_ _10630_ _11084_ VGND VGND
+ VPWR VPWR _12179_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_226_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17185_ decode.regfile.registers_15\[10\] _10611_ _10618_ _12583_ _12672_ VGND VGND
+ VPWR VPWR _13140_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_77_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14397_ _10074_ _10487_ VGND VGND VPWR VPWR _10488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16136_ decode.regfile.registers_8\[21\] _11045_ _11175_ VGND VGND VPWR VPWR _12112_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_133_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_1174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_228_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16067_ decode.regfile.registers_23\[19\] _11087_ _12016_ _12044_ VGND VGND VPWR
+ VPWR _12045_ sky130_fd_sc_hd__o22a_1
XFILLER_0_224_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15018_ _11027_ _11004_ _11006_ _11007_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__a31o_1
XFILLER_0_209_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2508 _10693_ VGND VGND VPWR VPWR net2735 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2519 csr._csr_read_data_T_8\[5\] VGND VGND VPWR VPWR net2746 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19826_ _03825_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1807 decode.regfile.registers_19\[30\] VGND VGND VPWR VPWR net2034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1818 fetch.bht.bhtTable_tag\[9\]\[0\] VGND VGND VPWR VPWR net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1829 fetch.bht.bhtTable_tag\[13\]\[9\] VGND VGND VPWR VPWR net2056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19757_ _04503_ _05031_ _04589_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16969_ decode.regfile.registers_11\[5\] _12594_ _12582_ _12550_ VGND VGND VPWR VPWR
+ _12929_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18708_ _03889_ decode.id_ex_imm_reg\[3\] VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__nand2_4
XFILLER_0_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19688_ _04965_ _04876_ _04268_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18639_ _03918_ _03923_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_101_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21650_ net1048 _06363_ _06364_ _06352_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_192_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20601_ csr.minstret\[22\] _05658_ _05735_ _05738_ _05537_ VGND VGND VPWR VPWR _05739_
+ sky130_fd_sc_hd__o221a_1
X_21581_ _06311_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23320_ net221 net222 net223 _07716_ net220 VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__a41o_1
XFILLER_0_156_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20532_ _05679_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23251_ _07088_ _07682_ _07683_ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__a21o_1
X_20463_ csr.mcycle\[4\] _05587_ _05594_ _05613_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22202_ fetch.bht.bhtTable_tag\[4\]\[24\] fetch.bht.bhtTable_tag\[5\]\[24\] _06618_
+ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__mux2_1
X_23182_ net74 _07536_ _07537_ _07618_ _07535_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__o311a_1
X_20394_ net295 _05516_ net358 _05522_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__or4_4
XFILLER_0_127_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22133_ _06685_ _06725_ _06627_ _06727_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_100_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27990_ clknet_leaf_223_clock _01012_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_26941_ _09956_ VGND VGND VPWR VPWR _09852_ sky130_fd_sc_hd__clkbuf_4
X_22064_ _06619_ fetch.bht.bhtTable_tag\[6\]\[18\] VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__and2b_1
XFILLER_0_199_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21015_ execute.io_reg_pc\[31\] _05989_ _05985_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26872_ net2084 _09809_ _09811_ _09812_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__o211a_1
X_29660_ clknet_leaf_288_clock _02673_ VGND VGND VPWR VPWR decode.regfile.registers_13\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28611_ clknet_leaf_132_clock _01624_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_25823_ _09128_ VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29591_ clknet_leaf_275_clock _02604_ VGND VGND VPWR VPWR decode.regfile.registers_10\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28542_ clknet_leaf_197_clock _01555_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_25754_ _10373_ _09932_ _08903_ _09935_ VGND VGND VPWR VPWR _09154_ sky130_fd_sc_hd__and4_1
X_22966_ execute.io_target_pc\[4\] _07346_ _07400_ _07414_ _07348_ VGND VGND VPWR
+ VPWR _07415_ sky130_fd_sc_hd__a2111o_1
X_24705_ _08536_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__clkbuf_1
X_21917_ _06551_ _06543_ _06544_ _06552_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__o211a_1
X_28473_ clknet_leaf_148_clock _01486_ VGND VGND VPWR VPWR decode.io_id_pc\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25685_ net2429 _09111_ _09114_ _09115_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22897_ _07347_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27424_ clknet_leaf_52_clock _00453_ VGND VGND VPWR VPWR decode.id_ex_isjump_reg
+ sky130_fd_sc_hd__dfxtp_1
X_24636_ net992 execute.io_target_pc\[7\] _08497_ VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21848_ net590 _06497_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27355_ clknet_leaf_47_clock _00384_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[28\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_194_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24567_ _08465_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21779_ net1347 _10771_ _06450_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26306_ net1593 _09475_ _09485_ _09484_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__o211a_1
X_14320_ net440 _10434_ _10443_ _10440_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23518_ net2300 _07890_ _07887_ VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__or3b_1
XFILLER_0_81_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27286_ clknet_leaf_7_clock _00315_ VGND VGND VPWR VPWR decode.regfile.registers_31\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24498_ _08057_ net2231 _08428_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__mux2_1
X_29025_ clknet_leaf_169_clock _02038_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14251_ _10087_ _10400_ VGND VGND VPWR VPWR _10404_ sky130_fd_sc_hd__nand2_1
X_26237_ _10373_ _10195_ _10196_ _08903_ VGND VGND VPWR VPWR _09445_ sky130_fd_sc_hd__and4_1
X_23449_ _10944_ _07847_ _07859_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__or3b_1
XFILLER_0_145_1315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14182_ net2611 _10359_ _10363_ _10357_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__o211a_1
X_26168_ net2339 _09395_ _09397_ _09394_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25119_ _06136_ net1692 _08778_ VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18990_ _03975_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__buf_6
X_26099_ _09328_ VGND VGND VPWR VPWR _09353_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17941_ decode.regfile.registers_17\[29\] _11022_ _12567_ _12586_ _12570_ VGND VGND
+ VPWR VPWR _03339_ sky130_fd_sc_hd__a41o_1
X_29927_ clknet_leaf_337_clock _02940_ VGND VGND VPWR VPWR decode.regfile.registers_21\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17872_ _12315_ _12630_ _12829_ _10614_ _03271_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__o221a_1
X_29858_ clknet_leaf_306_clock _02871_ VGND VGND VPWR VPWR decode.regfile.registers_19\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19611_ _03923_ _04443_ _04446_ _04202_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28809_ clknet_leaf_95_clock _01822_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16823_ _12497_ _12539_ _12503_ decode.regfile.registers_7\[2\] _12645_ VGND VGND
+ VPWR VPWR _12786_ sky130_fd_sc_hd__o32a_1
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29789_ clknet_leaf_309_clock _02802_ VGND VGND VPWR VPWR decode.regfile.registers_17\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19542_ _04805_ _04806_ _04810_ _04825_ _04729_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_176_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13966_ net2403 _10226_ _10237_ _10232_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__o211a_1
X_16754_ decode.regfile.registers_18\[1\] _10924_ _12568_ _12524_ _11008_ VGND VGND
+ VPWR VPWR _12718_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_191_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap3 _04400_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__buf_1
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15705_ _11046_ decode.regfile.registers_10\[10\] VGND VGND VPWR VPWR _11692_ sky130_fd_sc_hd__and2_1
XFILLER_0_216_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16685_ _12649_ VGND VGND VPWR VPWR _12650_ sky130_fd_sc_hd__buf_4
X_19473_ _04104_ _04112_ _04118_ net274 _04525_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__a41o_1
X_13897_ _10197_ VGND VGND VPWR VPWR _10198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_301 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_312 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18424_ _03721_ execute.io_mem_rd\[0\] _03722_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__a21oi_2
XINSDIODE1_323 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15636_ decode.regfile.registers_9\[8\] _11547_ _11623_ _11624_ _11184_ VGND VGND
+ VPWR VPWR _11625_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_334 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_345 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_356 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ decode.regfile.registers_19\[6\] _11354_ _11325_ _11557_ VGND VGND VPWR VPWR
+ _11558_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_367 decode.id_ex_imm_reg\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18355_ _03640_ decode.id_ex_ex_rs1_reg\[3\] _03650_ _03651_ _03653_ VGND VGND VPWR
+ VPWR _03654_ sky130_fd_sc_hd__o2111a_2
XINSDIODE1_378 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14518_ _09879_ _09882_ _10560_ _10562_ VGND VGND VPWR VPWR _10563_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_135_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17306_ _13221_ _13256_ _13257_ _13258_ VGND VGND VPWR VPWR _13259_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15498_ _11445_ _11488_ _11490_ VGND VGND VPWR VPWR _11491_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18286_ decode.id_ex_rs2_data_reg\[9\] _03605_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17237_ _12934_ _10592_ _12558_ decode.regfile.registers_0\[11\] VGND VGND VPWR VPWR
+ _13191_ sky130_fd_sc_hd__a31o_1
X_14449_ _10015_ _10517_ VGND VGND VPWR VPWR _10518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold904 fetch.bht.bhtTable_tag\[3\]\[21\] VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17168_ decode.regfile.registers_19\[9\] _11013_ _11012_ _12519_ _12545_ VGND VGND
+ VPWR VPWR _13124_ sky130_fd_sc_hd__o41a_1
XFILLER_0_40_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold915 decode.regfile.registers_3\[29\] VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold926 decode.io_id_pc\[2\] VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold937 fetch.bht.bhtTable_target_pc\[8\]\[30\] VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16119_ _11038_ VGND VGND VPWR VPWR _12095_ sky130_fd_sc_hd__buf_2
Xhold948 fetch.bht.bhtTable_target_pc\[7\]\[27\] VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold959 fetch.bht.bhtTable_tag\[3\]\[7\] VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__dlygate4sd3_1
X_17099_ _13055_ decode.regfile.registers_30\[8\] _12487_ VGND VGND VPWR VPWR _13056_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_1112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2305 decode.regfile.registers_26\[14\] VGND VGND VPWR VPWR net2532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2316 decode.regfile.registers_12\[20\] VGND VGND VPWR VPWR net2543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2327 decode.regfile.registers_23\[27\] VGND VGND VPWR VPWR net2554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2338 decode.regfile.registers_25\[24\] VGND VGND VPWR VPWR net2565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1604 fetch.bht.bhtTable_tag\[7\]\[6\] VGND VGND VPWR VPWR net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2349 decode.regfile.registers_8\[23\] VGND VGND VPWR VPWR net2576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1615 decode.regfile.registers_1\[4\] VGND VGND VPWR VPWR net1842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1626 _08478_ VGND VGND VPWR VPWR net1853 sky130_fd_sc_hd__dlygate4sd3_1
X_19809_ _05077_ _05078_ _04445_ _05081_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__a211o_1
Xhold1637 fetch.bht.bhtTable_target_pc\[14\]\[29\] VGND VGND VPWR VPWR net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 fetch.bht.bhtTable_tag\[0\]\[12\] VGND VGND VPWR VPWR net1875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1659 fetch.bht.bhtTable_tag\[9\]\[2\] VGND VGND VPWR VPWR net1886 sky130_fd_sc_hd__dlygate4sd3_1
X_22820_ _07305_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22751_ _07268_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21702_ _06363_ _06402_ _06403_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25470_ _08990_ VGND VGND VPWR VPWR _08991_ sky130_fd_sc_hd__clkbuf_4
X_22682_ net2551 _07222_ _07228_ _07221_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24421_ _08388_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21633_ _03579_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_191_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27140_ clknet_leaf_359_clock _00169_ VGND VGND VPWR VPWR decode.regfile.registers_26\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24352_ _08352_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__clkbuf_1
X_21564_ _06302_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23303_ _07619_ _07573_ _07620_ _07732_ VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20515_ _05664_ _03587_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__nor2_1
X_27071_ clknet_leaf_345_clock _00100_ VGND VGND VPWR VPWR decode.regfile.registers_24\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_24283_ _08111_ net1829 _06218_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21495_ _06124_ net2262 _06263_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26022_ _08943_ _09297_ VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__nand2_1
X_23234_ _07110_ _07667_ _07080_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__o21a_1
X_20446_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23165_ fetch.bht.bhtTable_target_pc\[4\]\[16\] fetch.bht.bhtTable_target_pc\[5\]\[16\]
+ fetch.bht.bhtTable_target_pc\[6\]\[16\] fetch.bht.bhtTable_target_pc\[7\]\[16\]
+ _07439_ _07112_ VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__mux4_1
X_20377_ _03721_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__buf_2
XFILLER_0_24_1006 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22116_ fetch.bht.bhtTable_tag\[8\]\[3\] fetch.bht.bhtTable_tag\[9\]\[3\] fetch.bht.bhtTable_tag\[10\]\[3\]
+ fetch.bht.bhtTable_tag\[11\]\[3\] _06617_ _06690_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27973_ clknet_leaf_200_clock _00995_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_23096_ _03500_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_228_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29712_ clknet_leaf_284_clock _02725_ VGND VGND VPWR VPWR decode.regfile.registers_14\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22047_ _06641_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__buf_4
X_26924_ net1125 _09839_ _09842_ _09836_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_162_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29643_ clknet_leaf_278_clock _02656_ VGND VGND VPWR VPWR decode.regfile.registers_12\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26855_ net1027 _09795_ _09802_ _09799_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13820_ _10152_ VGND VGND VPWR VPWR _10153_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25806_ _08954_ _09179_ VGND VGND VPWR VPWR _09185_ sky130_fd_sc_hd__nand2_1
X_29574_ clknet_leaf_273_clock _02587_ VGND VGND VPWR VPWR decode.regfile.registers_10\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_26786_ net1025 _09752_ _09762_ _09758_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23998_ _08170_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_218_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_218_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28525_ clknet_leaf_182_clock _01538_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13751_ _10003_ memory.io_wb_aluresult\[22\] _09981_ memory.io_wb_readdata\[22\]
+ _09995_ VGND VGND VPWR VPWR _10094_ sky130_fd_sc_hd__a221o_1
X_25737_ _08960_ _09136_ VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__nand2_1
X_22949_ _06032_ _07091_ _10915_ _07398_ VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__o31a_1
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16470_ _10642_ _11125_ _11104_ decode.regfile.registers_17\[30\] _11127_ VGND VGND
+ VPWR VPWR _12437_ sky130_fd_sc_hd__o32a_1
XFILLER_0_195_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28456_ clknet_leaf_148_clock _01469_ VGND VGND VPWR VPWR decode.io_id_pc\[14\] sky130_fd_sc_hd__dfxtp_1
X_25668_ net2529 _09095_ _09104_ _09100_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__o211a_1
X_13682_ _10035_ VGND VGND VPWR VPWR _10036_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15421_ _11152_ _11412_ _11413_ _11414_ VGND VGND VPWR VPWR _11415_ sky130_fd_sc_hd__a31o_1
X_24619_ net1193 execute.io_target_pc\[31\] _09897_ VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__mux2_1
X_27407_ clknet_leaf_9_clock _00436_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[16\]
+ sky130_fd_sc_hd__dfxtp_4
X_28387_ clknet_leaf_56_clock _01400_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_66_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25599_ net1961 _09026_ _09064_ _09059_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18140_ _03495_ _03493_ _03487_ net2298 VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__and4bb_1
X_27338_ clknet_leaf_155_clock _00367_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_15352_ _11079_ VGND VGND VPWR VPWR _11347_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_947 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14303_ _10418_ VGND VGND VPWR VPWR _10434_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_170_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18071_ _10972_ _10579_ _10948_ _10018_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15283_ decode.regfile.registers_13\[1\] _11276_ _11278_ decode.regfile.registers_12\[1\]
+ VGND VGND VPWR VPWR _11279_ sky130_fd_sc_hd__a22oi_1
X_27269_ clknet_leaf_14_clock _00298_ VGND VGND VPWR VPWR decode.regfile.registers_30\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17022_ decode.regfile.registers_12\[6\] _12551_ _12588_ _12979_ _12980_ VGND VGND
+ VPWR VPWR _12981_ sky130_fd_sc_hd__a32o_1
X_29008_ clknet_leaf_105_clock _02021_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire175 _00667_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14234_ _10048_ _10387_ VGND VGND VPWR VPWR _10394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_169_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire186 _07354_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_169_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire197 _10106_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_4
XFILLER_0_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14165_ net2478 _10346_ _10353_ _10344_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ net242 VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__clkbuf_4
X_14096_ _10081_ _10312_ VGND VGND VPWR VPWR _10314_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17924_ decode.regfile.registers_17\[28\] _12524_ _12568_ _12535_ _03322_ VGND VGND
+ VPWR VPWR _03323_ sky130_fd_sc_hd__a41o_1
XFILLER_0_219_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17855_ _10938_ decode.regfile.registers_25\[26\] _13482_ _12811_ VGND VGND VPWR
+ VPWR _03256_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16806_ decode.regfile.registers_23\[2\] _12714_ _12515_ VGND VGND VPWR VPWR _12769_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17786_ decode.regfile.registers_17\[25\] _12524_ _12568_ _12535_ _12571_ VGND VGND
+ VPWR VPWR _03188_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_50_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14998_ _11010_ VGND VGND VPWR VPWR _11011_ sky130_fd_sc_hd__buf_4
XFILLER_0_178_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19525_ _04245_ _04627_ _04294_ _04808_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__a211o_1
X_16737_ _12701_ _12500_ _10606_ _10937_ VGND VGND VPWR VPWR _12702_ sky130_fd_sc_hd__or4_4
XFILLER_0_53_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13949_ net2392 _10226_ _10228_ _10219_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19456_ net266 _04741_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__nor2_1
XFILLER_0_220_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16668_ _12597_ _10934_ _10605_ _10607_ VGND VGND VPWR VPWR _12633_ sky130_fd_sc_hd__nand4_2
XINSDIODE1_120 _11058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XINSDIODE1_131 _11318_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_142 _12504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18407_ decode.id_ex_immsrc_reg VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__buf_4
XFILLER_0_201_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_153 _12690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15619_ _11346_ _11253_ _11064_ decode.regfile.registers_29\[7\] _11608_ VGND VGND
+ VPWR VPWR _11609_ sky130_fd_sc_hd__o221a_1
X_19387_ _04357_ _04384_ _04349_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_164 decode.id_ex_rs1_data_reg\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16599_ _10598_ _10588_ _10618_ _12500_ VGND VGND VPWR VPWR _12564_ sky130_fd_sc_hd__or4_2
XINSDIODE1_175 decode.id_ex_rs2_data_reg\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINSDIODE1_186 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_197 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18338_ decode.id_ex_aluop_reg\[0\] VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18269_ _03588_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20300_ _10806_ decode.id_ex_pc_reg\[18\] _05468_ _05340_ VGND VGND VPWR VPWR _05476_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21280_ _06146_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__clkbuf_1
Xhold701 fetch.bht.bhtTable_target_pc\[4\]\[3\] VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold712 decode.regfile.registers_15\[11\] VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 fetch.bht.bhtTable_target_pc\[11\]\[26\] VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout5 _03773_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_4
X_20231_ _10834_ _10747_ _05415_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold734 fetch.bht.bhtTable_target_pc\[2\]\[24\] VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_203_Left_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold745 _08474_ VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold756 fetch.bht.bhtTable_target_pc\[6\]\[29\] VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold767 fetch.bht.bhtTable_tag\[8\]\[23\] VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20162_ decode.id_ex_imm_reg\[22\] _10864_ _05365_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__a21o_1
Xhold778 decode.regfile.registers_26\[5\] VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold789 fetch.bht.bhtTable_tag\[4\]\[20\] VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2102 decode.regfile.registers_19\[21\] VGND VGND VPWR VPWR net2329 sky130_fd_sc_hd__dlygate4sd3_1
X_20093_ _05303_ _05306_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__and2_1
Xhold2113 decode.regfile.registers_1\[6\] VGND VGND VPWR VPWR net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24970_ _07199_ _08691_ _08693_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__nor3_1
Xhold2124 decode.regfile.registers_9\[21\] VGND VGND VPWR VPWR net2351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2135 decode.regfile.registers_7\[5\] VGND VGND VPWR VPWR net2362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1401 fetch.bht.bhtTable_target_pc\[8\]\[4\] VGND VGND VPWR VPWR net1628 sky130_fd_sc_hd__dlygate4sd3_1
X_23921_ net895 _08078_ _08130_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__mux2_1
Xhold2146 decode.regfile.registers_5\[5\] VGND VGND VPWR VPWR net2373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2157 decode.regfile.registers_8\[6\] VGND VGND VPWR VPWR net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 execute.csr_write_data_out_reg\[26\] VGND VGND VPWR VPWR net1639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1423 decode.regfile.registers_7\[4\] VGND VGND VPWR VPWR net1650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2168 execute.csr_write_data_out_reg\[15\] VGND VGND VPWR VPWR net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 fetch.bht.bhtTable_tag\[1\]\[0\] VGND VGND VPWR VPWR net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2179 decode.regfile.registers_14\[22\] VGND VGND VPWR VPWR net2406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1445 fetch.bht.bhtTable_target_pc\[2\]\[12\] VGND VGND VPWR VPWR net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 fetch.bht.bhtTable_tag\[6\]\[7\] VGND VGND VPWR VPWR net1683 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26640_ net1988 _09665_ _09678_ _09675_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__o211a_1
X_23852_ execute.io_target_pc\[19\] VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__buf_2
Xhold1467 fetch.bht.bhtTable_tag\[2\]\[7\] VGND VGND VPWR VPWR net1694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1478 fetch.bht.bhtTable_tag\[10\]\[16\] VGND VGND VPWR VPWR net1705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1489 fetch.bht.bhtTable_tag\[13\]\[11\] VGND VGND VPWR VPWR net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22803_ _07296_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__clkbuf_1
X_26571_ _09400_ _09632_ VGND VGND VPWR VPWR _09639_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_212_Left_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23783_ _06145_ net1573 _08041_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20995_ execute.io_reg_pc\[22\] _05977_ _05973_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__and3_1
X_28310_ clknet_leaf_238_clock _01323_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_25522_ _08973_ _08978_ VGND VGND VPWR VPWR _09020_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22734_ _07259_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__clkbuf_1
X_29290_ clknet_leaf_231_clock _02303_ VGND VGND VPWR VPWR decode.regfile.registers_1\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28241_ clknet_leaf_76_clock _01263_ VGND VGND VPWR VPWR csr._minstret_T_3\[41\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_48_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25453_ _09950_ _08980_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__nand2_1
X_22665_ net2341 _07208_ _07218_ _07164_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24404_ _08379_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21616_ _05613_ csr.minstret\[5\] _06338_ _06339_ _06336_ VGND VGND VPWR VPWR _01122_
+ sky130_fd_sc_hd__a311oi_1
X_28172_ clknet_leaf_53_clock _01194_ VGND VGND VPWR VPWR csr.io_mret_vector\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25384_ net2382 _08928_ _08932_ _08927_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__o211a_1
X_22596_ csr._minstret_T_3\[46\] csr._minstret_T_3\[45\] csr._minstret_T_3\[44\] _07168_
+ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__and4_1
XFILLER_0_146_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27123_ clknet_leaf_354_clock _00152_ VGND VGND VPWR VPWR decode.regfile.registers_26\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_24335_ _08097_ net1727 _08334_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21547_ _06293_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27054_ clknet_leaf_333_clock _00083_ VGND VGND VPWR VPWR decode.regfile.registers_23\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_24266_ _08308_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_221_Left_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21478_ _06107_ net2193 _06252_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26005_ net2167 _09286_ _09299_ _09292_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__o211a_1
X_23217_ net224 net76 net75 _07613_ VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20429_ _05551_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24197_ _08091_ net1338 _08266_ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23148_ _07581_ _05246_ _07584_ _07586_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_164_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_219_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27956_ clknet_leaf_192_clock _00978_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_23079_ csr._csr_read_data_T_8\[11\] _06039_ csr.io_mret_vector\[11\] _06463_ VGND
+ VGND VPWR VPWR _07521_ sky130_fd_sc_hd__a22o_1
X_15970_ decode.regfile.registers_7\[17\] _11092_ _11142_ _11169_ decode.regfile.registers_6\[17\]
+ VGND VGND VPWR VPWR _11950_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_160_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_351_clock clknet_5_4__leaf_clock VGND VGND VPWR VPWR clknet_leaf_351_clock
+ sky130_fd_sc_hd__clkbuf_8
X_14921_ decode.control.io_opcode\[3\] _10585_ VGND VGND VPWR VPWR _10950_ sky130_fd_sc_hd__nor2_2
X_26907_ net2486 _09822_ _09831_ _09825_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27887_ clknet_leaf_23_clock _00916_ VGND VGND VPWR VPWR csr._mcycle_T_2\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29626_ clknet_leaf_288_clock _02639_ VGND VGND VPWR VPWR decode.regfile.registers_12\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _03043_ _03044_ _03045_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__a21oi_2
X_14852_ _10884_ _10885_ _10680_ VGND VGND VPWR VPWR _10895_ sky130_fd_sc_hd__a21o_1
X_26838_ net2034 _09753_ _09791_ _09784_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1990 decode.regfile.registers_16\[28\] VGND VGND VPWR VPWR net2217 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ _10021_ memory.io_wb_reg_pc\[30\] VGND VGND VPWR VPWR _10138_ sky130_fd_sc_hd__and2b_1
X_14783_ decode.id_ex_pc_reg\[31\] csr.io_mem_pc\[31\] VGND VGND VPWR VPWR _10826_
+ sky130_fd_sc_hd__xnor2_1
X_17571_ decode.regfile.registers_20\[19\] _12771_ _02977_ _02978_ _12538_ VGND VGND
+ VPWR VPWR _02979_ sky130_fd_sc_hd__a221o_1
X_29557_ clknet_leaf_274_clock _02570_ VGND VGND VPWR VPWR decode.regfile.registers_9\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26769_ _09751_ VGND VGND VPWR VPWR _09753_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_63_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19310_ _04436_ _04432_ _04371_ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__o22ai_1
X_28508_ clknet_leaf_212_clock _01521_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_16522_ _12486_ VGND VGND VPWR VPWR _12487_ sky130_fd_sc_hd__clkbuf_4
X_13734_ memory.csr_read_data_out_reg\[19\] _09986_ _10078_ _10079_ VGND VGND VPWR
+ VPWR _10080_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_98_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29488_ clknet_leaf_264_clock _02501_ VGND VGND VPWR VPWR decode.regfile.registers_7\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19241_ _04287_ _04533_ _04534_ _04535_ _04289_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28439_ clknet_leaf_49_clock _01452_ VGND VGND VPWR VPWR decode.control.io_funct7\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13665_ _09940_ VGND VGND VPWR VPWR _10021_ sky130_fd_sc_hd__clkbuf_4
X_16453_ decode.regfile.registers_7\[30\] _11308_ _11169_ decode.regfile.registers_6\[30\]
+ _11133_ VGND VGND VPWR VPWR _12420_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15404_ _10960_ decode.regfile.registers_28\[2\] _11398_ VGND VGND VPWR VPWR _11399_
+ sky130_fd_sc_hd__o21ai_1
X_16384_ decode.regfile.registers_0\[28\] _11154_ _12352_ VGND VGND VPWR VPWR _12353_
+ sky130_fd_sc_hd__a21oi_1
X_19172_ _03703_ _04324_ _04274_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__and3_2
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13596_ memory.io_wb_memtoreg\[1\] memory.io_wb_memtoreg\[0\] VGND VGND VPWR VPWR
+ _09960_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_22_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18123_ _03489_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_22_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15335_ _10992_ _11244_ _11261_ _11330_ VGND VGND VPWR VPWR _11331_ sky130_fd_sc_hd__a31o_1
XFILLER_0_170_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18054_ _10583_ _10584_ _10998_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__and3_1
X_15266_ _11086_ VGND VGND VPWR VPWR _11262_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_93_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_3 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_304_clock clknet_5_16__leaf_clock VGND VGND VPWR VPWR clknet_leaf_304_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14217_ _09999_ _10377_ VGND VGND VPWR VPWR _10384_ sky130_fd_sc_hd__nand2_1
X_17005_ _12708_ net582 _12923_ _12964_ _12705_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_188_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15197_ _11193_ VGND VGND VPWR VPWR _11194_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14148_ net1033 _10332_ _10343_ _10344_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14079_ _10036_ _10299_ VGND VGND VPWR VPWR _10305_ sky130_fd_sc_hd__nand2_1
X_18956_ _04254_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_52_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17907_ decode.regfile.registers_13\[28\] _12927_ _12583_ _12663_ VGND VGND VPWR
+ VPWR _03306_ sky130_fd_sc_hd__a31o_1
XFILLER_0_218_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18887_ _04086_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_175_Right_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17838_ decode.regfile.registers_9\[26\] _12603_ _03230_ _03238_ VGND VGND VPWR VPWR
+ _03239_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer15 _04021_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_2
Xrebuffer26 _03757_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_1
Xrebuffer37 net263 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_1
Xrebuffer48 _06615_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_2
X_17769_ _03149_ _03171_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__nor2_1
Xrebuffer59 net285 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19508_ _04289_ _04594_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__or2_1
X_20780_ net133 execute.io_mem_zero net99 _05861_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_187_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19439_ _04539_ _04709_ _04713_ _04726_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22450_ _06674_ fetch.btb.btbTable\[2\]\[1\] fetch.bht.bhtTable_valid\[2\] VGND VGND
+ VPWR VPWR _07045_ sky130_fd_sc_hd__and3b_1
XFILLER_0_85_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21401_ _06149_ net1578 _06210_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer105 net331 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_1
X_22381_ net223 _06975_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__xnor2_1
Xrebuffer116 _11150_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_1
X_24120_ net1380 VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21332_ _06176_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24051_ net1412 VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21263_ net945 _06134_ _06120_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__mux2_1
Xhold520 fetch.bht.bhtTable_tag\[11\]\[16\] VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 decode.regfile.registers_13\[4\] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 fetch.bht.bhtTable_tag\[12\]\[9\] VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__dlygate4sd3_1
X_23002_ _07447_ _07448_ _07368_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20214_ _05408_ _05409_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__xnor2_1
Xhold553 decode.regfile.registers_25\[15\] VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold564 csr._mcycle_T_3\[62\] VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__dlygate4sd3_1
X_21194_ _06092_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__clkbuf_1
Xhold575 decode.regfile.registers_21\[16\] VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 fetch.bht.bhtTable_target_pc\[4\]\[7\] VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold597 fetch.bht.bhtTable_tag\[4\]\[8\] VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1058 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27810_ clknet_leaf_35_clock _00839_ VGND VGND VPWR VPWR memory.io_wb_reg_pc\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20145_ decode.id_ex_imm_reg\[21\] _10798_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__nand2_1
X_28790_ clknet_leaf_126_clock _01803_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_202_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24953_ _07199_ _08680_ _08682_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__nor3_1
X_27741_ clknet_leaf_26_clock _00770_ VGND VGND VPWR VPWR decode.io_wb_rd\[4\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_198_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ decode.id_ex_imm_reg\[9\] _10706_ _05284_ _05291_ VGND VGND VPWR VPWR _05292_
+ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_198_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 fetch.bht.bhtTable_target_pc\[9\]\[25\] VGND VGND VPWR VPWR net1447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 fetch.bht.bhtTable_target_pc\[14\]\[0\] VGND VGND VPWR VPWR net1458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 fetch.bht.bhtTable_target_pc\[15\]\[8\] VGND VGND VPWR VPWR net1469 sky130_fd_sc_hd__dlygate4sd3_1
X_23904_ net1139 _08062_ _08119_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1253 fetch.bht.bhtTable_target_pc\[15\]\[17\] VGND VGND VPWR VPWR net1480 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24884_ _08633_ _03558_ csr.mcycle\[7\] csr.mcycle\[6\] VGND VGND VPWR VPWR _08634_
+ sky130_fd_sc_hd__and4_1
X_27672_ clknet_leaf_28_clock _00701_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[14\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold1264 decode.regfile.registers_14\[0\] VGND VGND VPWR VPWR net1491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1275 decode.regfile.registers_10\[27\] VGND VGND VPWR VPWR net1502 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_194_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29411_ clknet_leaf_247_clock _02424_ VGND VGND VPWR VPWR decode.regfile.registers_5\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_23835_ _08077_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_194_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 decode.regfile.registers_4\[11\] VGND VGND VPWR VPWR net1513 sky130_fd_sc_hd__dlygate4sd3_1
X_26623_ _09377_ _09666_ VGND VGND VPWR VPWR _09669_ sky130_fd_sc_hd__nand2_1
Xhold1297 csr._minstret_T_3\[58\] VGND VGND VPWR VPWR net1524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29342_ clknet_leaf_256_clock _02355_ VGND VGND VPWR VPWR decode.regfile.registers_3\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26554_ _09383_ _09623_ VGND VGND VPWR VPWR _09629_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23766_ _06128_ net1485 _08030_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20978_ _05971_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25505_ _08956_ _09005_ VGND VGND VPWR VPWR _09011_ sky130_fd_sc_hd__nand2_1
X_22717_ _10575_ _11000_ _11006_ _10586_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__or4b_1
X_29273_ clknet_leaf_235_clock _02286_ VGND VGND VPWR VPWR decode.regfile.registers_0\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_26485_ _09577_ VGND VGND VPWR VPWR _09589_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23697_ net840 csr.io_mem_pc\[12\] _07992_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_211_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_109_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28224_ clknet_leaf_86_clock net2015 VGND VGND VPWR VPWR csr.mscratch\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25436_ net191 VGND VGND VPWR VPWR _08968_ sky130_fd_sc_hd__clkbuf_8
X_22648_ _06457_ net217 _06458_ _06466_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__nand4_2
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28155_ clknet_leaf_64_clock _01177_ VGND VGND VPWR VPWR csr.ie sky130_fd_sc_hd__dfxtp_2
X_25367_ _10007_ VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__buf_4
X_22579_ net2712 _07162_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15120_ _11116_ VGND VGND VPWR VPWR _11117_ sky130_fd_sc_hd__buf_4
XFILLER_0_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24318_ _08335_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__clkbuf_1
X_27106_ clknet_leaf_357_clock _00135_ VGND VGND VPWR VPWR decode.regfile.registers_25\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_28086_ clknet_leaf_201_clock _01108_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25298_ _08879_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__clkbuf_1
X_15051_ _11047_ VGND VGND VPWR VPWR _11048_ sky130_fd_sc_hd__buf_4
X_27037_ clknet_leaf_338_clock _00066_ VGND VGND VPWR VPWR decode.regfile.registers_23\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_24249_ _08299_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14002_ _10036_ _10255_ VGND VGND VPWR VPWR _10260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Left_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18810_ execute.csr_read_data_out_reg\[12\] _03661_ _03660_ VGND VGND VPWR VPWR _04109_
+ sky130_fd_sc_hd__or3_1
Xoutput73 net73 VGND VGND VPWR VPWR io_fetch_address[15] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_290_clock clknet_5_17__leaf_clock VGND VGND VPWR VPWR clknet_leaf_290_clock
+ sky130_fd_sc_hd__clkbuf_8
Xoutput84 net84 VGND VGND VPWR VPWR io_fetch_address[25] sky130_fd_sc_hd__clkbuf_4
X_19790_ _04330_ _04965_ _04877_ _04537_ _04302_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28988_ clknet_leaf_184_clock _02001_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_183_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput95 net95 VGND VGND VPWR VPWR io_fetch_address[6] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_125_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18741_ execute.csr_read_data_out_reg\[5\] _03661_ _03660_ VGND VGND VPWR VPWR _04040_
+ sky130_fd_sc_hd__or3_1
X_27939_ clknet_leaf_217_clock _00961_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_15953_ decode.regfile.registers_20\[16\] _11452_ _11222_ _11933_ VGND VGND VPWR
+ VPWR _11934_ sky130_fd_sc_hd__a211o_1
XFILLER_0_216_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14904_ _10606_ _10577_ _10673_ _10911_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__nor4_1
X_18672_ _09974_ _03771_ _03969_ _03970_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__a211oi_4
XTAP_TAPCELL_ROW_121_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _11436_ decode.regfile.registers_26\[14\] _11676_ _11338_ _11564_ VGND VGND
+ VPWR VPWR _11867_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_188_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _13221_ _03027_ _03028_ _03029_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__a31o_1
X_29609_ clknet_leaf_275_clock _02622_ VGND VGND VPWR VPWR decode.regfile.registers_11\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ csr.io_mem_pc\[10\] VGND VGND VPWR VPWR _10878_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_2__f_clock clknet_2_0_0_clock VGND VGND VPWR VPWR clknet_5_2__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17554_ decode.regfile.registers_4\[19\] _12618_ _12620_ decode.regfile.registers_5\[19\]
+ _12737_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_203_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14766_ _10807_ _10808_ VGND VGND VPWR VPWR _10809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_127_Left_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16505_ decode.regfile.registers_16\[31\] _11359_ _12454_ _12470_ VGND VGND VPWR
+ VPWR _12471_ sky130_fd_sc_hd__o22a_1
X_13717_ net1824 _10027_ _10065_ _10020_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__o211a_1
X_14697_ _10719_ _10724_ _10727_ _10739_ VGND VGND VPWR VPWR _10740_ sky130_fd_sc_hd__nand4b_1
X_17485_ decode.regfile.registers_11\[17\] _12724_ _12587_ _12550_ _13432_ VGND VGND
+ VPWR VPWR _13433_ sky130_fd_sc_hd__a221o_2
XFILLER_0_85_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19224_ _04027_ _04028_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16436_ decode.regfile.registers_17\[29\] _10989_ _11114_ _11119_ _12403_ VGND VGND
+ VPWR VPWR _12404_ sky130_fd_sc_hd__a41o_1
XFILLER_0_67_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13648_ _10003_ memory.io_wb_aluresult\[7\] _10004_ memory.io_wb_readdata\[7\] _10005_
+ VGND VGND VPWR VPWR _10006_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19155_ _04401_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__buf_4
X_16367_ decode.regfile.registers_21\[27\] _11267_ _11098_ _11227_ _12336_ VGND VGND
+ VPWR VPWR _12337_ sky130_fd_sc_hd__o311a_1
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13579_ _09939_ memory.io_wb_aluresult\[0\] _09940_ VGND VGND VPWR VPWR _09944_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18106_ _03479_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_243_clock clknet_5_28__leaf_clock VGND VGND VPWR VPWR clknet_leaf_243_clock
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_41_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15318_ _11057_ _10628_ VGND VGND VPWR VPWR _11314_ sky130_fd_sc_hd__nand2_1
X_19086_ _04269_ _04378_ _04383_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__o21ai_1
X_16298_ _11679_ decode.regfile.registers_27\[25\] _11869_ VGND VGND VPWR VPWR _12270_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_14_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18037_ decode.regfile.registers_19\[31\] _11013_ _10589_ _12519_ _12544_ VGND VGND
+ VPWR VPWR _03433_ sky130_fd_sc_hd__o41a_1
XFILLER_0_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15249_ _11245_ VGND VGND VPWR VPWR _11246_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_258_clock clknet_5_23__leaf_clock VGND VGND VPWR VPWR clknet_leaf_258_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19988_ _10854_ _05214_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__and2_1
XFILLER_0_226_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18939_ _03867_ _04213_ _04170_ _04237_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__or4b_4
XFILLER_0_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21950_ net795 _06574_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20901_ _05925_ _05921_ net36 VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21881_ csr.io_mret_vector\[13\] _10871_ _06515_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23620_ _07956_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_145_Left_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20832_ _05892_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23551_ net2190 _07918_ _07915_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__or3b_1
X_20763_ _05850_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22502_ _03580_ _07096_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26270_ net2214 _09462_ _09465_ _09458_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23482_ decode.control.io_funct7\[1\] _07876_ _07873_ VGND VGND VPWR VPWR _07880_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_64_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20694_ _05813_ net700 VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25221_ _08060_ net963 _08837_ VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22433_ _06675_ _07027_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25152_ _06281_ _10569_ VGND VGND VPWR VPWR _08804_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22364_ _06957_ _06958_ _00002_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24103_ _08224_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21315_ _06167_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_154_Left_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25083_ net546 _08646_ _08769_ _06327_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22295_ _06887_ _06886_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_211_Right_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28911_ clknet_leaf_107_clock _01924_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[10\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_24034_ net999 execute.io_target_pc\[5\] _08187_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__mux2_1
X_21246_ _06123_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__clkbuf_1
Xhold350 decode.regfile.registers_1\[26\] VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29891_ clknet_leaf_303_clock _02904_ VGND VGND VPWR VPWR decode.regfile.registers_20\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold361 decode.regfile.registers_22\[9\] VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 decode.regfile.registers_5\[10\] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold383 decode.regfile.registers_30\[25\] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__dlygate4sd3_1
X_28842_ clknet_leaf_97_clock _01855_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold394 _08638_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21177_ _06083_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_225_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20128_ decode.id_ex_imm_reg\[17\] _10806_ _05336_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__o21ai_1
X_28773_ clknet_leaf_136_clock _01786_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_25985_ net2399 _09286_ _09288_ _09277_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_221_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27724_ clknet_leaf_24_clock _00753_ VGND VGND VPWR VPWR execute.csr_write_address_out_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20059_ _00556_ _05228_ _05277_ _05231_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__o22a_1
X_24936_ csr._mcycle_T_3\[47\] csr._mcycle_T_3\[46\] _08668_ _06422_ VGND VGND VPWR
+ VPWR _08671_ sky130_fd_sc_hd__a31o_1
Xhold1050 _08169_ VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 fetch.bht.bhtTable_target_pc\[1\]\[13\] VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_163_Left_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1072 fetch.bht.bhtTable_tag\[12\]\[19\] VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27655_ clknet_leaf_65_clock _00684_ VGND VGND VPWR VPWR execute.exception_out_reg
+ sky130_fd_sc_hd__dfxtp_1
Xhold1083 decode.regfile.registers_25\[0\] VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 fetch.bht.bhtTable_tag\[10\]\[20\] VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__dlygate4sd3_1
X_24867_ _08621_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26606_ _09436_ _09621_ VGND VGND VPWR VPWR _09658_ sky130_fd_sc_hd__nand2_1
X_14620_ _10662_ decode.id_ex_ex_rd_reg\[3\] VGND VGND VPWR VPWR _10663_ sky130_fd_sc_hd__nand2_1
X_23818_ execute.io_target_pc\[8\] VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__buf_2
X_24798_ _08091_ net1115 _08585_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27586_ clknet_leaf_136_clock _00615_ VGND VGND VPWR VPWR csr.io_mem_pc\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29325_ clknet_leaf_226_clock _02338_ VGND VGND VPWR VPWR decode.regfile.registers_2\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_14551_ _10593_ VGND VGND VPWR VPWR _10594_ sky130_fd_sc_hd__clkbuf_8
X_23749_ _06111_ net1583 _09907_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__mux2_1
X_26537_ _09443_ _09577_ VGND VGND VPWR VPWR _09618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13502_ _09883_ VGND VGND VPWR VPWR _09884_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29256_ clknet_leaf_231_clock _02269_ VGND VGND VPWR VPWR decode.regfile.registers_0\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_17270_ _10923_ _12876_ decode.regfile.registers_14\[12\] _12555_ VGND VGND VPWR
+ VPWR _13223_ sky130_fd_sc_hd__and4b_1
X_14482_ _10097_ _10530_ VGND VGND VPWR VPWR _10537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26468_ _10245_ _09579_ VGND VGND VPWR VPWR _09580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28207_ clknet_leaf_62_clock net885 VGND VGND VPWR VPWR csr.mscratch\[9\] sky130_fd_sc_hd__dfxtp_1
X_16221_ decode.regfile.registers_21\[23\] _11061_ _11099_ _11228_ _12194_ VGND VGND
+ VPWR VPWR _12195_ sky130_fd_sc_hd__o311a_1
X_25419_ _08956_ _08946_ VGND VGND VPWR VPWR _08957_ sky130_fd_sc_hd__nand2_1
X_29187_ clknet_leaf_240_clock _02200_ VGND VGND VPWR VPWR fetch.btb.btbTable\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_26399_ _09417_ VGND VGND VPWR VPWR _09540_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_114_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16152_ _11075_ _12126_ _12127_ _11486_ VGND VGND VPWR VPWR _12128_ sky130_fd_sc_hd__o211a_1
X_28138_ clknet_leaf_210_clock _01160_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer6 net232 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15103_ _11099_ VGND VGND VPWR VPWR _11100_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_185_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16083_ decode.regfile.registers_1\[20\] _11117_ _11057_ _11109_ VGND VGND VPWR VPWR
+ _12060_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_185_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28069_ clknet_leaf_166_clock _01091_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_185_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15034_ net433 _11028_ _11029_ _11031_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__a31o_1
X_19911_ _03704_ _04338_ _04320_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_75_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_208_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19842_ _04508_ _04728_ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19773_ _03849_ _05045_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_88_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16985_ decode.regfile.registers_10\[5\] _12653_ _12930_ _12944_ _12792_ VGND VGND
+ VPWR VPWR _12945_ sky130_fd_sc_hd__o221a_1
XFILLER_0_219_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18724_ _04014_ _04020_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15936_ decode.regfile.registers_2\[16\] _11369_ _11297_ _11121_ _11916_ VGND VGND
+ VPWR VPWR _11917_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_155_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18655_ _03707_ decode.id_ex_imm_reg\[20\] VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__nand2_2
XFILLER_0_204_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15867_ decode.regfile.registers_7\[14\] _11465_ _11169_ decode.regfile.registers_6\[14\]
+ _11165_ VGND VGND VPWR VPWR _11850_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17606_ decode.regfile.registers_12\[20\] _12541_ _12772_ _12658_ _03012_ VGND VGND
+ VPWR VPWR _03013_ sky130_fd_sc_hd__o311a_1
X_14818_ csr.io_mem_pc\[24\] _10768_ VGND VGND VPWR VPWR _10861_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_47_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18586_ net114 _03666_ _03884_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_176_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15798_ decode.regfile.registers_16\[12\] _11203_ _11357_ VGND VGND VPWR VPWR _11783_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_47_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17537_ _11010_ VGND VGND VPWR VPWR _13484_ sky130_fd_sc_hd__buf_2
XFILLER_0_86_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14749_ csr.io_mem_pc\[24\] csr.io_mem_pc\[25\] _10768_ VGND VGND VPWR VPWR _10792_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_103_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17468_ _10926_ decode.regfile.registers_22\[17\] _12554_ _11009_ _12546_ VGND VGND
+ VPWR VPWR _13416_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19207_ _03638_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__buf_4
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_182_clock clknet_5_26__leaf_clock VGND VGND VPWR VPWR clknet_leaf_182_clock
+ sky130_fd_sc_hd__clkbuf_8
X_16419_ decode.regfile.registers_1\[29\] VGND VGND VPWR VPWR _12387_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17399_ decode.regfile.registers_7\[15\] _12611_ _12888_ VGND VGND VPWR VPWR _13349_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19138_ _04249_ _04333_ _04434_ _04327_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_225_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19069_ _03863_ _04233_ net187 VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_197_clock clknet_5_30__leaf_clock VGND VGND VPWR VPWR clknet_leaf_197_clock
+ sky130_fd_sc_hd__clkbuf_8
X_21100_ _10970_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__buf_4
X_22080_ _06649_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21031_ _06000_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_120_clock clknet_5_14__leaf_clock VGND VGND VPWR VPWR clknet_leaf_120_clock
+ sky130_fd_sc_hd__clkbuf_8
X_22982_ _07426_ _10758_ _07429_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__or3b_1
X_25770_ _08918_ _09157_ VGND VGND VPWR VPWR _09164_ sky130_fd_sc_hd__nand2_1
X_24721_ _08083_ net1772 _08542_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__mux2_1
X_21933_ csr.io_mret_vector\[29\] csr.io_mem_pc\[29\] _06481_ VGND VGND VPWR VPWR
+ _06563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_135_clock clknet_5_15__leaf_clock VGND VGND VPWR VPWR clknet_leaf_135_clock
+ sky130_fd_sc_hd__clkbuf_8
X_24652_ _08509_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27440_ clknet_leaf_146_clock _00469_ VGND VGND VPWR VPWR decode.id_ex_pc_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21864_ _06513_ _06494_ _06495_ _06514_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23603_ _07947_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20815_ net126 _05879_ _05875_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__and3_1
X_24583_ net971 execute.io_target_pc\[13\] _08473_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__mux2_1
X_27371_ clknet_leaf_9_clock _00400_ VGND VGND VPWR VPWR decode.id_ex_rs2_data_reg\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_194_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21795_ csr.ie _05857_ _06463_ csr.pie _06464_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29110_ clknet_leaf_18_clock _02123_ VGND VGND VPWR VPWR csr._mcycle_T_3\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23534_ net2771 _07904_ _07901_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__or3b_1
X_26322_ net632 _09491_ _09495_ _09484_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__o211a_1
X_20746_ _05818_ decode.id_ex_rs1_data_reg\[30\] _03585_ VGND VGND VPWR VPWR _05844_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29041_ clknet_leaf_103_clock _02054_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[14\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_189_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26253_ net538 _09447_ _09455_ _09440_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23465_ net11 _07861_ _07869_ _07865_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20677_ decode.id_ex_rs1_data_reg\[3\] decode.id_ex_ex_rs1_reg\[3\] _05056_ VGND
+ VGND VPWR VPWR _05802_ sky130_fd_sc_hd__mux2_1
X_25204_ _10572_ fetch.btb.btbTable\[1\]\[1\] _08830_ VGND VGND VPWR VPWR _08831_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22416_ fetch.bht.bhtTable_tag\[8\]\[1\] fetch.bht.bhtTable_tag\[9\]\[1\] fetch.bht.bhtTable_tag\[10\]\[1\]
+ fetch.bht.bhtTable_tag\[11\]\[1\] _06674_ _06650_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__mux4_1
XFILLER_0_150_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26184_ _10063_ VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23396_ net90 net88 _06795_ _07783_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__nand4_2
XFILLER_0_116_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25135_ _06153_ net1505 _08562_ VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__mux2_1
X_22347_ _06790_ _06937_ _06939_ _06941_ _06640_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_143_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_227_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_227_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_227_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25066_ csr._mcycle_T_2\[26\] _08712_ _08757_ csr.mcycle\[25\] csr.mcycle\[26\] VGND
+ VGND VPWR VPWR _08758_ sky130_fd_sc_hd__a221oi_1
X_29943_ clknet_leaf_339_clock _02956_ VGND VGND VPWR VPWR decode.regfile.registers_21\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22278_ _06651_ _06872_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_148_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_148_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24017_ net886 execute.io_target_pc\[29\] _07960_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21229_ net2150 _06111_ _09912_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__mux2_1
Xhold180 fetch.btb.btbTable\[7\]\[0\] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold191 _00765_ VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
X_29874_ clknet_leaf_300_clock _02887_ VGND VGND VPWR VPWR decode.regfile.registers_19\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_217_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28825_ clknet_leaf_127_clock _01838_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_171_Left_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_219_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28756_ clknet_leaf_124_clock _01769_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_16770_ _12729_ _12730_ _12733_ VGND VGND VPWR VPWR _12734_ sky130_fd_sc_hd__o21a_1
X_13982_ _10131_ VGND VGND VPWR VPWR _10249_ sky130_fd_sc_hd__clkbuf_4
X_25968_ _08964_ _09267_ VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_107_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _11199_ _11706_ _11707_ VGND VGND VPWR VPWR _11708_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_5_20__f_clock clknet_2_2_0_clock VGND VGND VPWR VPWR clknet_5_20__leaf_clock
+ sky130_fd_sc_hd__clkbuf_16
X_27707_ clknet_leaf_20_clock _00736_ VGND VGND VPWR VPWR execute.csr_write_data_out_reg\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_24919_ csr._mcycle_T_3\[41\] csr._mcycle_T_3\[40\] csr._mcycle_T_3\[39\] _08656_
+ _07148_ VGND VGND VPWR VPWR _08660_ sky130_fd_sc_hd__a41o_1
X_28687_ clknet_leaf_112_clock _01700_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_25899_ decode.regfile.registers_7\[29\] _09226_ _09237_ _09235_ VGND VGND VPWR VPWR
+ _02508_ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ decode.io_wb_rd\[3\] _03719_ _03735_ _03736_ _03738_ VGND VGND VPWR VPWR
+ _03739_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_178_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27638_ clknet_leaf_45_clock net173 VGND VGND VPWR VPWR execute.io_reg_pc\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _11075_ _11639_ _11640_ _11236_ VGND VGND VPWR VPWR _11641_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_70 _10130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_198_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XINSDIODE1_81 _10588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_92 _10606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14603_ _10645_ VGND VGND VPWR VPWR _10646_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18371_ _03669_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__buf_4
X_27569_ clknet_leaf_159_clock _00598_ VGND VGND VPWR VPWR csr.io_mem_pc\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15583_ _11263_ decode.regfile.registers_22\[7\] _11404_ _10978_ _10990_ VGND VGND
+ VPWR VPWR _11573_ sky130_fd_sc_hd__o2111a_1
X_29308_ clknet_leaf_244_clock _02321_ VGND VGND VPWR VPWR decode.regfile.registers_2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17322_ _13267_ _13273_ _12892_ decode.regfile.registers_8\[13\] VGND VGND VPWR VPWR
+ _13274_ sky130_fd_sc_hd__o2bb2ai_1
X_14534_ _10576_ VGND VGND VPWR VPWR _10577_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_180_Left_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29239_ clknet_leaf_181_clock _02252_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[9\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17253_ decode.regfile.registers_22\[11\] _12528_ _13206_ _12687_ VGND VGND VPWR
+ VPWR _13207_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14465_ _10058_ _10517_ VGND VGND VPWR VPWR _10527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16204_ decode.regfile.registers_2\[23\] _11191_ _11149_ _11152_ _12177_ VGND VGND
+ VPWR VPWR _12178_ sky130_fd_sc_hd__o311a_1
XFILLER_0_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_226_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17184_ decode.regfile.registers_20\[10\] _11024_ _12553_ _12554_ _12537_ VGND VGND
+ VPWR VPWR _13139_ sky130_fd_sc_hd__a41o_1
X_14396_ _10462_ VGND VGND VPWR VPWR _10487_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_77_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16135_ _11289_ _12109_ _12110_ VGND VGND VPWR VPWR _12111_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_133_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_1186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16066_ decode.regfile.registers_21\[19\] _11267_ _11099_ _11228_ _12043_ VGND VGND
+ VPWR VPWR _12044_ sky130_fd_sc_hd__o311a_1
X_15017_ _11026_ VGND VGND VPWR VPWR _11027_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2509 csr._csr_read_data_T_8\[24\] VGND VGND VPWR VPWR net2736 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_36_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19825_ _04708_ _04924_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1808 fetch.bht.bhtTable_target_pc\[7\]\[6\] VGND VGND VPWR VPWR net2035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1819 fetch.bht.bhtTable_tag\[6\]\[0\] VGND VGND VPWR VPWR net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19756_ _03847_ _03844_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__and2b_1
X_16968_ decode.regfile.registers_13\[5\] _12927_ _12587_ _12663_ VGND VGND VPWR VPWR
+ _12928_ sky130_fd_sc_hd__a31o_1
XFILLER_0_223_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_52_clock clknet_5_12__leaf_clock VGND VGND VPWR VPWR clknet_leaf_52_clock
+ sky130_fd_sc_hd__clkbuf_8
X_18707_ _04004_ _04005_ _03997_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__nand3_2
XFILLER_0_155_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15919_ decode.regfile.registers_19\[15\] _11453_ _11454_ _11900_ VGND VGND VPWR
+ VPWR _11901_ sky130_fd_sc_hd__o211a_1
X_19687_ _04964_ _04918_ _04247_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16899_ _11015_ _10937_ decode.regfile.registers_23\[3\] _12520_ VGND VGND VPWR VPWR
+ _12861_ sky130_fd_sc_hd__or4_1
XFILLER_0_91_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18638_ _03898_ _03899_ _03902_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18569_ memory.csr_read_data_out_reg\[23\] _09987_ _10099_ _10100_ VGND VGND VPWR
+ VPWR _03868_ sky130_fd_sc_hd__o22a_2
Xclkbuf_leaf_67_clock clknet_5_9__leaf_clock VGND VGND VPWR VPWR clknet_leaf_67_clock
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20600_ csr.mscratch\[22\] _05591_ _05611_ _05736_ _05737_ VGND VGND VPWR VPWR _05738_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_47_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21580_ _06151_ net1805 _06306_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20531_ _10909_ _05678_ _09954_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23250_ execute.io_target_pc\[20\] _10757_ _10970_ _06037_ VGND VGND VPWR VPWR _07683_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_172_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20462_ _05617_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22201_ fetch.bht.bhtTable_tag\[0\]\[24\] fetch.bht.bhtTable_tag\[1\]\[24\] fetch.bht.bhtTable_tag\[2\]\[24\]
+ fetch.bht.bhtTable_tag\[3\]\[24\] _06646_ _06652_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23181_ _07611_ _07615_ _07617_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__a21o_1
XFILLER_0_160_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20393_ _05534_ csr.minstret\[0\] _05538_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22132_ _06684_ _06726_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22063_ _06657_ _06629_ _06642_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__a21o_1
X_26940_ _10024_ _09849_ VGND VGND VPWR VPWR _09851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21014_ _05991_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26871_ _09701_ VGND VGND VPWR VPWR _09812_ sky130_fd_sc_hd__buf_2
XFILLER_0_226_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28610_ clknet_leaf_133_clock _01623_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25822_ _08970_ _09155_ VGND VGND VPWR VPWR _09193_ sky130_fd_sc_hd__nand2_1
X_29590_ clknet_leaf_275_clock _02603_ VGND VGND VPWR VPWR decode.regfile.registers_10\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_28541_ clknet_leaf_192_clock _01554_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_22965_ _07368_ _07410_ _05246_ _07413_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__a211oi_1
X_25753_ net1987 _09112_ _09152_ _09153_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__o211a_1
X_24704_ _08066_ net1551 _08531_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21916_ net723 _06545_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__or2_1
X_28472_ clknet_leaf_138_clock _01485_ VGND VGND VPWR VPWR decode.io_id_pc\[30\] sky130_fd_sc_hd__dfxtp_1
X_22896_ _03592_ _10672_ _03590_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__and3_2
X_25684_ _08990_ VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_1208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27423_ clknet_leaf_41_clock _00452_ VGND VGND VPWR VPWR decode.id_ex_islui_reg sky130_fd_sc_hd__dfxtp_1
X_24635_ _08500_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__clkbuf_1
X_21847_ csr.io_mret_vector\[3\] _10557_ _06040_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_216_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24566_ net1161 execute.io_target_pc\[5\] _08462_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__mux2_1
X_27354_ clknet_leaf_47_clock _00383_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[27\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21778_ _06452_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26305_ _09436_ _09446_ VGND VGND VPWR VPWR _09485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_915 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23517_ _06718_ _07889_ _07899_ _07893_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__o211a_1
X_20729_ decode.id_ex_funct3_reg\[0\] _05804_ _05834_ _03517_ _03581_ VGND VGND VPWR
+ VPWR _05835_ sky130_fd_sc_hd__a2111oi_1
X_24497_ _08429_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__clkbuf_1
X_27285_ clknet_leaf_30_clock _00314_ VGND VGND VPWR VPWR decode.regfile.registers_31\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29024_ clknet_leaf_170_clock _02037_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14250_ _10375_ VGND VGND VPWR VPWR _10403_ sky130_fd_sc_hd__buf_2
X_23448_ decode.id_ex_memread_reg VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__clkbuf_2
X_26236_ net872 _09374_ _09444_ _09440_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14181_ _10102_ _10355_ VGND VGND VPWR VPWR _10363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23379_ _07619_ _07345_ _07620_ _07803_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__a31o_1
X_26167_ _09396_ _09390_ VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25118_ _08787_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26098_ net1758 _09343_ _09352_ _09346_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_72_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25049_ csr._mcycle_T_2\[21\] _08710_ _08645_ csr.mcycle\[21\] VGND VGND VPWR VPWR
+ _08746_ sky130_fd_sc_hd__a211oi_1
X_29926_ clknet_leaf_340_clock _02939_ VGND VGND VPWR VPWR decode.regfile.registers_21\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_17940_ decode.regfile.registers_20\[29\] _12525_ _12552_ _12523_ _12536_ VGND VGND
+ VPWR VPWR _03338_ sky130_fd_sc_hd__a41o_1
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17871_ _12630_ decode.regfile.registers_0\[27\] VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__nand2_1
X_29857_ clknet_leaf_306_clock _02870_ VGND VGND VPWR VPWR decode.regfile.registers_19\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19610_ _04886_ _04887_ _04505_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__o211a_1
X_28808_ clknet_leaf_99_clock _01821_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16822_ decode.regfile.registers_6\[2\] _10602_ _12615_ _12783_ _12784_ VGND VGND
+ VPWR VPWR _12785_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_105_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29788_ clknet_leaf_313_clock _02801_ VGND VGND VPWR VPWR decode.regfile.registers_17\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19541_ _04811_ _04465_ _04817_ _04303_ _04824_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_221_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28739_ clknet_leaf_130_clock _01752_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16753_ decode.regfile.registers_20\[1\] _12525_ _12552_ _12523_ _12536_ VGND VGND
+ VPWR VPWR _12717_ sky130_fd_sc_hd__a41o_1
XFILLER_0_219_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13965_ _10136_ _10198_ VGND VGND VPWR VPWR _10237_ sky130_fd_sc_hd__nand2_1
X_15704_ decode.regfile.registers_11\[10\] _11071_ _11204_ _11407_ VGND VGND VPWR
+ VPWR _11691_ sky130_fd_sc_hd__a31o_1
X_19472_ _04118_ _04112_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__nand2_1
X_16684_ _12637_ VGND VGND VPWR VPWR _12649_ sky130_fd_sc_hd__buf_4
XFILLER_0_201_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13896_ _09930_ _10195_ _10149_ _10196_ VGND VGND VPWR VPWR _10197_ sky130_fd_sc_hd__and4b_1
XFILLER_0_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_302 decode.id_ex_rs1_data_reg\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18423_ decode.id_ex_ex_use_rs2_reg execute.io_mem_regwrite VGND VGND VPWR VPWR _03722_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_1191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15635_ decode.regfile.registers_8\[8\] _11045_ _11175_ VGND VGND VPWR VPWR _11624_
+ sky130_fd_sc_hd__a21o_1
XINSDIODE1_313 decode.id_ex_rs1_data_reg\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_324 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_335 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE1_346 net139 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_201_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XINSDIODE1_357 _11037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18354_ _03652_ execute.io_mem_rd\[4\] VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__nand2_1
XINSDIODE1_368 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _11106_ _11555_ _11556_ VGND VGND VPWR VPWR _11557_ sky130_fd_sc_hd__a21o_1
XINSDIODE1_379 _07099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17305_ _13215_ decode.regfile.registers_28\[12\] _13093_ VGND VGND VPWR VPWR _13258_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14517_ _09879_ _10561_ _09882_ VGND VGND VPWR VPWR _10562_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_135_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18285_ _03607_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15497_ _11489_ decode.regfile.registers_28\[4\] decode.regfile.registers_29\[4\]
+ _11255_ _11246_ VGND VGND VPWR VPWR _11490_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_61_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17236_ decode.regfile.registers_9\[11\] _12602_ _12653_ VGND VGND VPWR VPWR _13190_
+ sky130_fd_sc_hd__o21ai_1
X_14448_ _10505_ VGND VGND VPWR VPWR _10517_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17167_ decode.regfile.registers_18\[9\] _12572_ _13121_ _13122_ _12562_ VGND VGND
+ VPWR VPWR _13123_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold905 fetch.bht.bhtTable_tag\[1\]\[15\] VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14379_ _10031_ _10474_ VGND VGND VPWR VPWR _10478_ sky130_fd_sc_hd__nand2_1
Xhold916 fetch.bht.bhtTable_target_pc\[2\]\[3\] VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold927 decode.regfile.registers_10\[20\] VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16118_ _11761_ net822 _12054_ _12094_ _11760_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__o221a_1
Xhold938 decode.regfile.registers_12\[29\] VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 fetch.bht.bhtTable_tag\[10\]\[21\] VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17098_ _10930_ VGND VGND VPWR VPWR _13055_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16049_ decode.regfile.registers_5\[19\] _11290_ _10636_ _11135_ VGND VGND VPWR VPWR
+ _12027_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2306 csr.msie VGND VGND VPWR VPWR net2533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2317 decode.regfile.registers_9\[27\] VGND VGND VPWR VPWR net2544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2328 decode.regfile.registers_9\[3\] VGND VGND VPWR VPWR net2555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2339 decode.regfile.registers_24\[24\] VGND VGND VPWR VPWR net2566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1605 fetch.bht.bhtTable_target_pc\[10\]\[17\] VGND VGND VPWR VPWR net1832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1616 fetch.bht.bhtTable_target_pc\[0\]\[0\] VGND VGND VPWR VPWR net1843 sky130_fd_sc_hd__dlygate4sd3_1
X_19808_ _05079_ net212 _05080_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__and3_1
Xhold1627 decode.regfile.registers_15\[6\] VGND VGND VPWR VPWR net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1638 fetch.bht.bhtTable_target_pc\[13\]\[7\] VGND VGND VPWR VPWR net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1649 decode.regfile.registers_25\[3\] VGND VGND VPWR VPWR net1876 sky130_fd_sc_hd__dlygate4sd3_1
X_19739_ _04974_ _04995_ _04191_ _04192_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__and4_1
XFILLER_0_205_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22750_ _06124_ net1648 _07265_ VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21701_ csr.minstret\[15\] csr.minstret\[25\] csr.minstret\[26\] csr.io_inst_retired
+ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22681_ csr._mcycle_T_2\[16\] _07223_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24420_ _08387_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__buf_6
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21632_ csr._mcycle_T_2\[10\] _06325_ _06340_ _06349_ csr.minstret\[10\] VGND VGND
+ VPWR VPWR _06351_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_133_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24351_ _08113_ net1742 _06187_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__mux2_1
X_21563_ _06134_ net2225 _06295_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23302_ csr._csr_read_data_T_8\[23\] _07416_ csr.io_mret_vector\[23\] _07621_ _07731_
+ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_211_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20514_ csr.mcycle\[10\] _05588_ _05663_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27070_ clknet_leaf_347_clock _00099_ VGND VGND VPWR VPWR decode.regfile.registers_24\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_24282_ _08316_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__clkbuf_1
X_21494_ _06264_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23233_ fetch.bht.bhtTable_target_pc\[0\]\[19\] fetch.bht.bhtTable_target_pc\[1\]\[19\]
+ _07067_ VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26021_ net2247 _09300_ _09308_ _09305_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__o211a_1
X_20445_ _05565_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__buf_2
XFILLER_0_160_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23164_ net73 _07536_ _07537_ _07601_ _07535_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__o311a_1
X_20376_ _03718_ net293 net358 _03741_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__or4_2
XFILLER_0_24_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_189_Right_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22115_ _06623_ _06705_ _06628_ _06709_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_100_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27972_ clknet_leaf_196_clock _00994_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_23095_ _06248_ VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__buf_2
XFILLER_0_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29711_ clknet_leaf_284_clock _02724_ VGND VGND VPWR VPWR decode.regfile.registers_14\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_22046_ _06640_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__buf_4
X_26923_ _09450_ _09840_ VGND VGND VPWR VPWR _09842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_228_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29642_ clknet_leaf_276_clock _02655_ VGND VGND VPWR VPWR decode.regfile.registers_12\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_162_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26854_ _09381_ _09796_ VGND VGND VPWR VPWR _09802_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_162_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25805_ net1280 _09183_ _09184_ _09182_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__o211a_1
X_29573_ clknet_leaf_273_clock _02586_ VGND VGND VPWR VPWR decode.regfile.registers_10\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26785_ _09387_ _09753_ VGND VGND VPWR VPWR _09762_ sky130_fd_sc_hd__nand2_1
X_23997_ net799 execute.io_target_pc\[19\] _08164_ VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_218_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28524_ clknet_leaf_168_clock _01537_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_218_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13750_ net2547 _10083_ _10093_ _10077_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__o211a_1
X_25736_ net2480 _09139_ _09144_ _09142_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_218_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22948_ csr._csr_read_data_T_8\[3\] _06481_ csr.io_mret_vector\[3\] _06463_ _07397_
+ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__a221o_1
XFILLER_0_168_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_1174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28455_ clknet_leaf_148_clock _01468_ VGND VGND VPWR VPWR decode.io_id_pc\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25667_ _08966_ _09092_ VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13681_ net545 _09988_ _10033_ _10034_ VGND VGND VPWR VPWR _10035_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_85_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22879_ _07336_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_1304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15420_ decode.regfile.registers_3\[3\] _11109_ _11141_ _11145_ VGND VGND VPWR VPWR
+ _11414_ sky130_fd_sc_hd__a31o_1
X_27406_ clknet_leaf_29_clock _00435_ VGND VGND VPWR VPWR decode.id_ex_rs1_data_reg\[15\]
+ sky130_fd_sc_hd__dfxtp_4
X_24618_ _08491_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28386_ clknet_leaf_144_clock _01399_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_167_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25598_ _08973_ _09023_ VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27337_ clknet_leaf_46_clock _00366_ VGND VGND VPWR VPWR decode.id_ex_imm_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15351_ _10961_ VGND VGND VPWR VPWR _11346_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24549_ _08109_ net1794 _09902_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14302_ net703 _10419_ _10433_ _10427_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18070_ _10997_ _03458_ _10969_ _03453_ _10999_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__o41a_1
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27268_ clknet_leaf_12_clock _00297_ VGND VGND VPWR VPWR decode.regfile.registers_30\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_15282_ _11277_ VGND VGND VPWR VPWR _11278_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29007_ clknet_leaf_107_clock _02020_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[13\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17021_ _12499_ _12541_ _12490_ decode.regfile.registers_11\[6\] _12878_ VGND VGND
+ VPWR VPWR _12980_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_130_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14233_ net2242 _10390_ _10393_ _10385_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__o211a_1
X_26219_ _09432_ _09413_ VGND VGND VPWR VPWR _09433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire176 net177 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27199_ clknet_leaf_361_clock _00228_ VGND VGND VPWR VPWR decode.regfile.registers_28\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xwire187 _04366_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
XFILLER_0_184_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_169_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14164_ _10064_ _10342_ VGND VGND VPWR VPWR _10353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_1059 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18972_ _04259_ _04267_ _04270_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__mux2_1
X_14095_ net2160 _10302_ _10313_ _10304_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_91_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ decode.regfile.registers_16\[28\] _13011_ _03305_ _03321_ _12578_ VGND VGND
+ VPWR VPWR _03322_ sky130_fd_sc_hd__o221a_1
XFILLER_0_221_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29909_ clknet_leaf_301_clock _02922_ VGND VGND VPWR VPWR decode.regfile.registers_20\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17854_ _13339_ _03252_ _03253_ _03254_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__a31o_1
XFILLER_0_206_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16805_ _12767_ VGND VGND VPWR VPWR _12768_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17785_ decode.regfile.registers_19\[25\] _12679_ _12906_ VGND VGND VPWR VPWR _03187_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14997_ _11009_ VGND VGND VPWR VPWR _11010_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19524_ _04245_ _04607_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__nor2_1
X_16736_ _10928_ VGND VGND VPWR VPWR _12701_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13948_ _10092_ _10223_ VGND VGND VPWR VPWR _10228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_220_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19455_ _04741_ net263 VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16667_ decode.regfile.registers_1\[0\] decode.regfile.registers_0\[0\] _12631_ VGND
+ VGND VPWR VPWR _12632_ sky130_fd_sc_hd__mux2_1
X_13879_ net2319 _10180_ _10186_ _10175_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__o211a_1
XINSDIODE1_110 _10935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_121 _11085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_202_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18406_ _03704_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__clkbuf_4
XINSDIODE1_132 _11347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_143 _12504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15618_ _11403_ _11605_ _11606_ _11607_ VGND VGND VPWR VPWR _11608_ sky130_fd_sc_hd__a31o_1
X_19386_ _04465_ _04670_ _04428_ _04675_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_158_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XINSDIODE1_154 _12690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16598_ _12546_ _12553_ _12554_ _12562_ decode.regfile.registers_19\[0\] VGND VGND
+ VPWR VPWR _12563_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XINSDIODE1_165 decode.id_ex_rs1_data_reg\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_176 decode.id_ex_rs2_data_reg\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18337_ _03633_ _03634_ _03635_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__or3b_4
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XINSDIODE1_187 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XINSDIODE1_198 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15549_ _11129_ _11147_ _11300_ decode.regfile.registers_1\[6\] VGND VGND VPWR VPWR
+ _11540_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18268_ decode.id_ex_rs2_data_reg\[1\] VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17219_ _13087_ decode.regfile.registers_26\[10\] _12814_ _13047_ _13088_ VGND VGND
+ VPWR VPWR _13174_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_170_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18199_ _10943_ decode.control.io_funct3\[0\] decode.control.io_funct3\[2\] VGND
+ VGND VPWR VPWR _03537_ sky130_fd_sc_hd__or3b_1
XFILLER_0_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold702 fetch.bht.bhtTable_target_pc\[12\]\[24\] VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20230_ _10834_ _10747_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__nand2_1
Xhold713 csr._mcycle_T_3\[56\] VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 fetch.bht.bhtTable_target_pc\[12\]\[10\] VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 decode.regfile.registers_24\[5\] VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 fetch.bht.bhtTable_target_pc\[8\]\[27\] VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 fetch.bht.bhtTable_tag\[8\]\[3\] VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold768 fetch.bht.bhtTable_target_pc\[12\]\[14\] VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__dlygate4sd3_1
X_20161_ _05359_ _05360_ _05361_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__a21oi_2
Xhold779 fetch.bht.bhtTable_tag\[4\]\[16\] VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2103 decode.regfile.registers_15\[1\] VGND VGND VPWR VPWR net2330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2114 csr._csr_read_data_T_8\[9\] VGND VGND VPWR VPWR net2341 sky130_fd_sc_hd__dlygate4sd3_1
X_20092_ _05296_ _05305_ _05301_ _05302_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2125 decode.regfile.registers_22\[24\] VGND VGND VPWR VPWR net2352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2136 decode.regfile.registers_18\[27\] VGND VGND VPWR VPWR net2363 sky130_fd_sc_hd__dlygate4sd3_1
X_23920_ _06155_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__clkbuf_8
Xhold2147 fetch.bht.bhtTable_target_pc\[14\]\[31\] VGND VGND VPWR VPWR net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1402 fetch.bht.bhtTable_tag\[0\]\[8\] VGND VGND VPWR VPWR net1629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1413 fetch.bht.bhtTable_target_pc\[9\]\[17\] VGND VGND VPWR VPWR net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2158 decode.regfile.registers_1\[19\] VGND VGND VPWR VPWR net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1424 decode.regfile.registers_10\[30\] VGND VGND VPWR VPWR net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2169 decode.regfile.registers_13\[14\] VGND VGND VPWR VPWR net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1435 fetch.bht.bhtTable_target_pc\[7\]\[5\] VGND VGND VPWR VPWR net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1446 fetch.bht.bhtTable_target_pc\[7\]\[30\] VGND VGND VPWR VPWR net1673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1457 fetch.bht.bhtTable_target_pc\[9\]\[13\] VGND VGND VPWR VPWR net1684 sky130_fd_sc_hd__dlygate4sd3_1
X_23851_ _08088_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_1342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1468 decode.regfile.registers_23\[26\] VGND VGND VPWR VPWR net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1479 fetch.bht.bhtTable_tag\[13\]\[25\] VGND VGND VPWR VPWR net1706 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_200_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22802_ net769 _10807_ _07286_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_200_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26570_ net1678 _09636_ _09638_ _09635_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_196_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23782_ _08043_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__clkbuf_1
X_20994_ _05980_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25521_ net2067 _09008_ _09019_ _09017_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22733_ _06107_ net1604 _09903_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_213_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28240_ clknet_leaf_73_clock _01262_ VGND VGND VPWR VPWR csr._minstret_T_3\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22664_ csr._mcycle_T_2\[9\] _07210_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__or2_1
X_25452_ _08978_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__buf_2
XFILLER_0_177_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24403_ net942 execute.io_target_pc\[24\] _09911_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__mux2_1
X_21615_ net2799 _06325_ _06338_ _05613_ csr.minstret\[5\] VGND VGND VPWR VPWR _06339_
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_30_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28171_ clknet_leaf_56_clock _01193_ VGND VGND VPWR VPWR csr.io_mret_vector\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_22595_ csr._minstret_T_3\[46\] _07172_ _07173_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__o21ba_1
X_25383_ _08931_ _08923_ VGND VGND VPWR VPWR _08932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27122_ clknet_leaf_351_clock _00151_ VGND VGND VPWR VPWR decode.regfile.registers_26\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_24334_ _08343_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__clkbuf_1
X_21546_ _06117_ net2047 _06284_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24265_ _08093_ net1431 _08300_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27053_ clknet_leaf_331_clock _00082_ VGND VGND VPWR VPWR decode.regfile.registers_23\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_21477_ _06255_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23216_ net76 _07536_ _07537_ _07650_ _07535_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__o311a_1
XFILLER_0_161_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26004_ _08925_ _09297_ VGND VGND VPWR VPWR _09299_ sky130_fd_sc_hd__nand2_1
X_20428_ _05585_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24196_ _08272_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23147_ csr._csr_read_data_T_8\[14\] _06461_ csr.io_mret_vector\[14\] _07417_ _07585_
+ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_164_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20359_ _05521_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_164_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27955_ clknet_leaf_191_clock _00977_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_23078_ net68 _07343_ _07344_ _07520_ _06566_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__o311a_1
XFILLER_0_105_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22029_ _06623_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__clkbuf_4
X_14920_ decode.control.io_opcode\[4\] _10580_ _10579_ decode.control.io_opcode\[5\]
+ VGND VGND VPWR VPWR _10949_ sky130_fd_sc_hd__and4b_1
X_26906_ _09434_ _09819_ VGND VGND VPWR VPWR _09831_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27886_ clknet_leaf_66_clock _00915_ VGND VGND VPWR VPWR csr._mcycle_T_2\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29625_ clknet_leaf_289_clock _02638_ VGND VGND VPWR VPWR decode.regfile.registers_11\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ _10888_ _10890_ _10892_ _10893_ VGND VGND VPWR VPWR _10894_ sky130_fd_sc_hd__a211oi_1
X_26837_ _09441_ _09751_ VGND VGND VPWR VPWR _09791_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13802_ net702 _10083_ _10137_ _10132_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__o211a_1
X_17570_ decode.regfile.registers_19\[19\] _11013_ _10589_ _12519_ _12544_ VGND VGND
+ VPWR VPWR _02978_ sky130_fd_sc_hd__o41a_1
Xhold1980 decode.regfile.registers_25\[30\] VGND VGND VPWR VPWR net2207 sky130_fd_sc_hd__dlygate4sd3_1
X_29556_ clknet_leaf_266_clock _02569_ VGND VGND VPWR VPWR decode.regfile.registers_9\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_14782_ _10748_ _09892_ _09894_ VGND VGND VPWR VPWR _10825_ sky130_fd_sc_hd__nor3_1
Xhold1991 decode.regfile.registers_24\[18\] VGND VGND VPWR VPWR net2218 sky130_fd_sc_hd__dlygate4sd3_1
X_26768_ _09751_ VGND VGND VPWR VPWR _09752_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28507_ clknet_leaf_216_clock _01520_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16521_ _11027_ _11015_ _11012_ _11011_ VGND VGND VPWR VPWR _12486_ sky130_fd_sc_hd__and4_2
X_13733_ _10003_ memory.io_wb_aluresult\[19\] _10001_ memory.io_wb_reg_pc\[19\] _09995_
+ VGND VGND VPWR VPWR _10079_ sky130_fd_sc_hd__a221o_1
X_25719_ net1657 _09125_ _09134_ _09129_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29487_ clknet_leaf_264_clock _02500_ VGND VGND VPWR VPWR decode.regfile.registers_7\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_26699_ _09377_ _09710_ VGND VGND VPWR VPWR _09713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19240_ _04278_ _04267_ net244 VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28438_ clknet_leaf_48_clock _01451_ VGND VGND VPWR VPWR decode.control.io_funct7\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16452_ decode.regfile.registers_11\[30\] net322 _11167_ _11277_ VGND VGND VPWR VPWR
+ _12419_ sky130_fd_sc_hd__a31o_1
X_13664_ net831 _09938_ _10017_ _10020_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15403_ _11347_ _11037_ _11066_ VGND VGND VPWR VPWR _11398_ sky130_fd_sc_hd__and3_1
XFILLER_0_186_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19171_ _04443_ _04362_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28369_ clknet_leaf_211_clock _01382_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_16383_ decode.regfile.registers_1\[28\] _11116_ _11137_ _11157_ VGND VGND VPWR VPWR
+ _12352_ sky130_fd_sc_hd__and4_1
XFILLER_0_27_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_225_Right_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13595_ memory.io_wb_memtoreg\[1\] memory.io_wb_readdata\[1\] _09958_ VGND VGND VPWR
+ VPWR _09959_ sky130_fd_sc_hd__o21a_1
X_18122_ _03482_ _03480_ _03487_ decode.io_id_pc\[17\] VGND VGND VPWR VPWR _03489_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_26_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15334_ decode.regfile.registers_23\[1\] _11262_ _11266_ _11329_ VGND VGND VPWR VPWR
+ _11330_ sky130_fd_sc_hd__o22a_1
XFILLER_0_87_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18053_ _03447_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15265_ _11072_ VGND VGND VPWR VPWR _11261_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_4 _01442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17004_ _12765_ _12768_ _12493_ decode.regfile.registers_29\[5\] _12963_ VGND VGND
+ VPWR VPWR _12964_ sky130_fd_sc_hd__o221a_1
XFILLER_0_227_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14216_ net931 _10376_ _10383_ _10369_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15196_ _11191_ _10630_ _11192_ _11051_ VGND VGND VPWR VPWR _11193_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14147_ _10290_ VGND VGND VPWR VPWR _10344_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14078_ net1990 _10302_ _10303_ _10304_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__o211a_1
X_18955_ _04253_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_197_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17906_ decode.regfile.registers_15\[28\] _12555_ _10619_ _12876_ _13031_ VGND VGND
+ VPWR VPWR _03305_ sky130_fd_sc_hd__a41o_1
X_18886_ _04112_ _04115_ net283 _04103_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17837_ _12612_ _03236_ _03237_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer16 net242 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer27 _04094_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_222_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17768_ _03169_ _12566_ _03170_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__a21oi_1
Xrebuffer38 net263 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
Xrebuffer49 _06615_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_1
XFILLER_0_117_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19507_ _04691_ _04791_ _04272_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__mux2_1
X_16719_ decode.regfile.registers_21\[0\] _12538_ _12683_ VGND VGND VPWR VPWR _12684_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17699_ _02986_ decode.regfile.registers_26\[22\] _13254_ _13484_ _02987_ VGND VGND
+ VPWR VPWR _03104_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_92_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19438_ _04155_ _04714_ _04444_ _04725_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_187_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19369_ _04612_ _04621_ _04132_ _04144_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21400_ _06213_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22380_ _06968_ _06636_ _06974_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_143_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer106 net331 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_1
Xrebuffer117 _11150_ VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21331_ net1386 csr.io_mem_pc\[23\] _06168_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24050_ net1411 execute.io_target_pc\[13\] _08187_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__mux2_1
X_21262_ _10787_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__buf_2
Xhold510 io_fetch_data[7] VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold521 decode.regfile.registers_11\[7\] VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__dlygate4sd3_1
X_23001_ net227 _07427_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__nand2_1
Xhold532 csr._mcycle_T_3\[49\] VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold543 csr.mcycle\[23\] VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__buf_1
X_20213_ decode.id_ex_imm_reg\[31\] decode.id_ex_pc_reg\[31\] VGND VGND VPWR VPWR
+ _05409_ sky130_fd_sc_hd__xor2_1
Xhold554 fetch.bht.bhtTable_tag\[12\]\[13\] VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 decode.regfile.registers_1\[0\] VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__dlygate4sd3_1
X_21193_ _06086_ _06082_ net403 VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold576 decode.regfile.registers_4\[1\] VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 fetch.bht.bhtTable_target_pc\[1\]\[20\] VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_206_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20144_ decode.id_ex_imm_reg\[21\] _10798_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold598 execute.csr_write_data_out_reg\[6\] VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27740_ clknet_leaf_34_clock _00769_ VGND VGND VPWR VPWR decode.io_wb_rd\[3\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_202_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20075_ _05279_ _05285_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__nand2_1
X_24952_ _08681_ VGND VGND VPWR VPWR _08682_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_202_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _08236_ VGND VGND VPWR VPWR net1437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 fetch.bht.bhtTable_target_pc\[3\]\[10\] VGND VGND VPWR VPWR net1448 sky130_fd_sc_hd__dlygate4sd3_1
X_23903_ _08121_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__clkbuf_1
Xhold1232 fetch.bht.bhtTable_tag\[4\]\[19\] VGND VGND VPWR VPWR net1459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1243 fetch.bht.bhtTable_target_pc\[3\]\[1\] VGND VGND VPWR VPWR net1470 sky130_fd_sc_hd__dlygate4sd3_1
X_27671_ clknet_leaf_28_clock _00700_ VGND VGND VPWR VPWR execute.csr_read_data_out_reg\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_24883_ csr.io_csr_write_address\[11\] net216 _06314_ _06459_ VGND VGND VPWR VPWR
+ _08633_ sky130_fd_sc_hd__nand4_4
Xhold1254 fetch.bht.bhtTable_target_pc\[3\]\[8\] VGND VGND VPWR VPWR net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 fetch.bht.bhtTable_target_pc\[8\]\[1\] VGND VGND VPWR VPWR net1492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29410_ clknet_leaf_247_clock _02423_ VGND VGND VPWR VPWR decode.regfile.registers_5\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1276 fetch.bht.bhtTable_target_pc\[3\]\[22\] VGND VGND VPWR VPWR net1503 sky130_fd_sc_hd__dlygate4sd3_1
X_26622_ net2043 _09665_ _09668_ _09660_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__o211a_1
X_23834_ _08076_ net1462 _08058_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_194_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1287 decode.regfile.registers_20\[18\] VGND VGND VPWR VPWR net1514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 decode.regfile.registers_1\[1\] VGND VGND VPWR VPWR net1525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_1309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_29341_ clknet_leaf_244_clock _02354_ VGND VGND VPWR VPWR decode.regfile.registers_3\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26553_ net1116 _09622_ _09628_ _09619_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__o211a_1
X_23765_ _08034_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20977_ net2583 _05965_ _05961_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25504_ decode.regfile.registers_2\[21\] _09008_ _09010_ _09004_ VGND VGND VPWR VPWR
+ _02340_ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22716_ csr._csr_read_data_T_8\[31\] _07235_ _07246_ _07247_ VGND VGND VPWR VPWR
+ _01315_ sky130_fd_sc_hd__o211a_1
X_29272_ clknet_leaf_232_clock _02285_ VGND VGND VPWR VPWR decode.regfile.registers_0\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26484_ net2353 _09578_ _09588_ _09582_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__o211a_1
X_23696_ _07998_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28223_ clknet_leaf_86_clock net527 VGND VGND VPWR VPWR csr.mscratch\[25\] sky130_fd_sc_hd__dfxtp_1
X_25435_ net570 _08951_ _08967_ _08950_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22647_ _07207_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_28154_ clknet_leaf_157_clock _01176_ VGND VGND VPWR VPWR fetch.btb.io_branch sky130_fd_sc_hd__dfxtp_1
X_22578_ csr._minstret_T_3\[40\] _06420_ _07161_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__and3_1
X_25366_ net2340 _08906_ _08919_ _07247_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27105_ clknet_leaf_357_clock _00134_ VGND VGND VPWR VPWR decode.regfile.registers_25\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24317_ _08078_ net2011 _08334_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__mux2_1
X_28085_ clknet_leaf_200_clock _01107_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[13\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_21529_ _06283_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25297_ _08869_ net2701 VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27036_ clknet_leaf_342_clock _00065_ VGND VGND VPWR VPWR decode.regfile.registers_23\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_15050_ _11046_ VGND VGND VPWR VPWR _11047_ sky130_fd_sc_hd__buf_4
X_24248_ _08076_ net1934 _08289_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14001_ net1042 _10258_ _10259_ _10249_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_112_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24179_ _08263_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput74 net74 VGND VGND VPWR VPWR io_fetch_address[16] sky130_fd_sc_hd__clkbuf_4
X_28987_ clknet_leaf_172_clock _02000_ VGND VGND VPWR VPWR fetch.bht.bhtTable_target_pc\[12\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_183_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput85 net85 VGND VGND VPWR VPWR io_fetch_address[26] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 net96 VGND VGND VPWR VPWR io_fetch_address[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18740_ _04034_ _04038_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_27938_ clknet_leaf_223_clock _00960_ VGND VGND VPWR VPWR fetch.bht.bhtTable_tag\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_15952_ decode.regfile.registers_19\[16\] _11453_ _11219_ _11932_ VGND VGND VPWR
+ VPWR _11933_ sky130_fd_sc_hd__o211a_1
X_14903_ _10937_ _10577_ _10673_ _10911_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__nor4_1
X_18671_ decode.id_ex_rs1_data_reg\[3\] net247 VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__nor2_2
X_15883_ _11050_ decode.regfile.registers_25\[14\] _11090_ VGND VGND VPWR VPWR _11866_
+ sky130_fd_sc_hd__or3_1
X_27869_ clknet_leaf_327_clock _00898_ VGND VGND VPWR VPWR memory.csr_read_data_out_reg\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17622_ _13215_ decode.regfile.registers_28\[20\] _02992_ VGND VGND VPWR VPWR _03029_
+ sky130_fd_sc_hd__o21a_1
X_14834_ _10808_ _10876_ VGND VGND VPWR VPWR _10877_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29608_ clknet_leaf_276_clock _02621_ VGND VGND VPWR VPWR decode.regfile.registers_11\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ decode.regfile.registers_3\[19\] _12629_ _13496_ _02960_ VGND VGND VPWR VPWR
+ _02961_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_54_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29539_ clknet_leaf_252_clock _02552_ VGND VGND VPWR VPWR decode.regfile.registers_9\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14765_ csr.io_mem_pc\[13\] csr.io_mem_pc\[14\] _10763_ VGND VGND VPWR VPWR _10808_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_129_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16504_ _10650_ _10625_ _11053_ _12455_ _12469_ VGND VGND VPWR VPWR _12470_ sky130_fd_sc_hd__o32a_1
X_13716_ _10064_ _10016_ VGND VGND VPWR VPWR _10065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17484_ _12599_ _13430_ _13431_ _12791_ VGND VGND VPWR VPWR _13432_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14696_ _10675_ execute.io_target_pc\[16\] _10729_ _10735_ _10738_ VGND VGND VPWR
+ VPWR _10739_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19223_ _04027_ _04028_ _04448_ _04517_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16435_ _11124_ decode.regfile.registers_16\[29\] _11128_ _12402_ VGND VGND VPWR
+ VPWR _12403_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_15_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13647_ _09977_ VGND VGND VPWR VPWR _10005_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19154_ _04006_ _03983_ _04320_ _04003_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16366_ decode.regfile.registers_20\[27\] _11102_ _11327_ _12335_ VGND VGND VPWR
+ VPWR _12336_ sky130_fd_sc_hd__a211o_1
XFILLER_0_186_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13578_ _09939_ VGND VGND VPWR VPWR _09943_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18105_ _03469_ _03467_ _03474_ decode.io_id_pc\[10\] VGND VGND VPWR VPWR _03479_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_147_1027 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15317_ _11042_ VGND VGND VPWR VPWR _11313_ sky130_fd_sc_hd__clkbuf_4
X_19085_ _04280_ _04282_ _04382_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16297_ _11260_ _12266_ _12267_ _12268_ VGND VGND VPWR VPWR _12269_ sky130_fd_sc_hd__a31o_1
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18036_ decode.regfile.registers_18\[31\] _12572_ _03430_ _03431_ _12562_ VGND VGND
+ VPWR VPWR _03432_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15248_ _10958_ _11054_ _11062_ _11244_ VGND VGND VPWR VPWR _11245_ sky130_fd_sc_hd__or4_4
XFILLER_0_169_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15179_ decode.regfile.registers_8\[0\] _11046_ _11175_ VGND VGND VPWR VPWR _11176_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19987_ net2386 _05219_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18938_ _04052_ _04039_ _04025_ _04236_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__and4_1
.ends

